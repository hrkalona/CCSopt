// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module c499(N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,
  N73,N77,N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
  N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
  N137;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
  N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755;

  wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
    N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
    N282,N283,N284,N285,N286,N287,N288,N289,N290,N293,N296,N299,N302,N305,N308,N311,
    N314,N315,N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,N342,N343,N344,N345,
    N346,N347,N348,N349,N350,N351,N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
    N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,
    N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,
    N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,
    N602,N607,N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,N694,N695,N696,N697,
    N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
    N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,extra0,extra1,extra2,extra3,extra4,extra5,
    extra6,extra7;

  XOR2_X1 XOR2_1( .Z(N250), .A(N1), .B(N5) );
  XOR2_X1 XOR2_2( .Z(N251), .A(N9), .B(N13) );
  XOR2_X2 XOR2_3( .Z(N252), .A(N17), .B(N21) );
  XOR2_X2 XOR2_4( .Z(N253), .A(N25), .B(N29) );
  XOR2_X2 XOR2_5( .Z(N254), .A(N33), .B(N37) );
  XOR2_X1 XOR2_6( .Z(N255), .A(N41), .B(N45) );
  XOR2_X1 XOR2_7( .Z(N256), .A(N49), .B(N53) );
  XOR2_X1 XOR2_8( .Z(N257), .A(N57), .B(N61) );
  XOR2_X1 XOR2_9( .Z(N258), .A(N65), .B(N69) );
  XOR2_X1 XOR2_10( .Z(N259), .A(N73), .B(N77) );
  XOR2_X1 XOR2_11( .Z(N260), .A(N81), .B(N85) );
  XOR2_X1 XOR2_12( .Z(N261), .A(N89), .B(N93) );
  XOR2_X1 XOR2_13( .Z(N262), .A(N97), .B(N101) );
  XOR2_X1 XOR2_14( .Z(N263), .A(N105), .B(N109) );
  XOR2_X1 XOR2_15( .Z(N264), .A(N113), .B(N117) );
  XOR2_X1 XOR2_16( .Z(N265), .A(N121), .B(N125) );
  AND2_X1 AND2_17( .ZN(N266), .A1(N129), .A2(N137) );
  AND2_X1 AND2_18( .ZN(N267), .A1(N130), .A2(N137) );
  AND2_X1 AND2_19( .ZN(N268), .A1(N131), .A2(N137) );
  AND2_X1 AND2_20( .ZN(N269), .A1(N132), .A2(N137) );
  AND2_X1 AND2_21( .ZN(N270), .A1(N133), .A2(N137) );
  AND2_X1 AND2_22( .ZN(N271), .A1(N134), .A2(N137) );
  AND2_X1 AND2_23( .ZN(N272), .A1(N135), .A2(N137) );
  AND2_X1 AND2_24( .ZN(N273), .A1(N136), .A2(N137) );
  XOR2_X1 XOR2_25( .Z(N274), .A(N1), .B(N17) );
  XOR2_X1 XOR2_26( .Z(N275), .A(N33), .B(N49) );
  XOR2_X1 XOR2_27( .Z(N276), .A(N5), .B(N21) );
  XOR2_X1 XOR2_28( .Z(N277), .A(N37), .B(N53) );
  XOR2_X2 XOR2_29( .Z(N278), .A(N9), .B(N25) );
  XOR2_X2 XOR2_30( .Z(N279), .A(N41), .B(N57) );
  XOR2_X2 XOR2_31( .Z(N280), .A(N13), .B(N29) );
  XOR2_X2 XOR2_32( .Z(N281), .A(N45), .B(N61) );
  XOR2_X1 XOR2_33( .Z(N282), .A(N65), .B(N81) );
  XOR2_X1 XOR2_34( .Z(N283), .A(N97), .B(N113) );
  XOR2_X1 XOR2_35( .Z(N284), .A(N69), .B(N85) );
  XOR2_X1 XOR2_36( .Z(N285), .A(N101), .B(N117) );
  XOR2_X1 XOR2_37( .Z(N286), .A(N73), .B(N89) );
  XOR2_X1 XOR2_38( .Z(N287), .A(N105), .B(N121) );
  XOR2_X1 XOR2_39( .Z(N288), .A(N77), .B(N93) );
  XOR2_X1 XOR2_40( .Z(N289), .A(N109), .B(N125) );
  XOR2_X1 XOR2_41( .Z(N290), .A(N250), .B(N251) );
  XOR2_X1 XOR2_42( .Z(N293), .A(N252), .B(N253) );
  XOR2_X1 XOR2_43( .Z(N296), .A(N254), .B(N255) );
  XOR2_X1 XOR2_44( .Z(N299), .A(N256), .B(N257) );
  XOR2_X1 XOR2_45( .Z(N302), .A(N258), .B(N259) );
  XOR2_X1 XOR2_46( .Z(N305), .A(N260), .B(N261) );
  XOR2_X1 XOR2_47( .Z(N308), .A(N262), .B(N263) );
  XOR2_X1 XOR2_48( .Z(N311), .A(N264), .B(N265) );
  XOR2_X1 XOR2_49( .Z(N314), .A(N274), .B(N275) );
  XOR2_X1 XOR2_50( .Z(N315), .A(N276), .B(N277) );
  XOR2_X1 XOR2_51( .Z(N316), .A(N278), .B(N279) );
  XOR2_X1 XOR2_52( .Z(N317), .A(N280), .B(N281) );
  XOR2_X1 XOR2_53( .Z(N318), .A(N282), .B(N283) );
  XOR2_X1 XOR2_54( .Z(N319), .A(N284), .B(N285) );
  XOR2_X1 XOR2_55( .Z(N320), .A(N286), .B(N287) );
  XOR2_X1 XOR2_56( .Z(N321), .A(N288), .B(N289) );
  XOR2_X1 XOR2_57( .Z(N338), .A(N290), .B(N293) );
  XOR2_X1 XOR2_58( .Z(N339), .A(N296), .B(N299) );
  XOR2_X1 XOR2_59( .Z(N340), .A(N290), .B(N296) );
  XOR2_X1 XOR2_60( .Z(N341), .A(N293), .B(N299) );
  XOR2_X2 XOR2_61( .Z(N342), .A(N302), .B(N305) );
  XOR2_X2 XOR2_62( .Z(N343), .A(N308), .B(N311) );
  XOR2_X2 XOR2_63( .Z(N344), .A(N302), .B(N308) );
  XOR2_X1 XOR2_64( .Z(N345), .A(N305), .B(N311) );
  XOR2_X1 XOR2_65( .Z(N346), .A(N266), .B(N342) );
  XOR2_X1 XOR2_66( .Z(N347), .A(N267), .B(N343) );
  XOR2_X1 XOR2_67( .Z(N348), .A(N268), .B(N344) );
  XOR2_X1 XOR2_68( .Z(N349), .A(N269), .B(N345) );
  XOR2_X1 XOR2_69( .Z(N350), .A(N270), .B(N338) );
  XOR2_X1 XOR2_70( .Z(N351), .A(N271), .B(N339) );
  XOR2_X1 XOR2_71( .Z(N352), .A(N272), .B(N340) );
  XOR2_X1 XOR2_72( .Z(N353), .A(N273), .B(N341) );
  XOR2_X1 XOR2_73( .Z(N354), .A(N314), .B(N346) );
  XOR2_X1 XOR2_74( .Z(N367), .A(N315), .B(N347) );
  XOR2_X1 XOR2_75( .Z(N380), .A(N316), .B(N348) );
  XOR2_X1 XOR2_76( .Z(N393), .A(N317), .B(N349) );
  XOR2_X1 XOR2_77( .Z(N406), .A(N318), .B(N350) );
  XOR2_X1 XOR2_78( .Z(N419), .A(N319), .B(N351) );
  XOR2_X1 XOR2_79( .Z(N432), .A(N320), .B(N352) );
  XOR2_X1 XOR2_80( .Z(N445), .A(N321), .B(N353) );
  INV_X1 NOT1_81( .ZN(N554), .A(N354) );
  INV_X1 NOT1_82( .ZN(N555), .A(N367) );
  INV_X1 NOT1_83( .ZN(N556), .A(N380) );
  INV_X1 NOT1_84( .ZN(N557), .A(N354) );
  INV_X1 NOT1_85( .ZN(N558), .A(N367) );
  INV_X1 NOT1_86( .ZN(N559), .A(N393) );
  INV_X4 NOT1_87( .ZN(N560), .A(N354) );
  INV_X4 NOT1_88( .ZN(N561), .A(N380) );
  INV_X1 NOT1_89( .ZN(N562), .A(N393) );
  INV_X1 NOT1_90( .ZN(N563), .A(N367) );
  INV_X1 NOT1_91( .ZN(N564), .A(N380) );
  INV_X1 NOT1_92( .ZN(N565), .A(N393) );
  INV_X1 NOT1_93( .ZN(N566), .A(N419) );
  INV_X1 NOT1_94( .ZN(N567), .A(N445) );
  INV_X1 NOT1_95( .ZN(N568), .A(N419) );
  INV_X1 NOT1_96( .ZN(N569), .A(N432) );
  INV_X1 NOT1_97( .ZN(N570), .A(N406) );
  INV_X1 NOT1_98( .ZN(N571), .A(N445) );
  INV_X1 NOT1_99( .ZN(N572), .A(N406) );
  INV_X1 NOT1_100( .ZN(N573), .A(N432) );
  INV_X1 NOT1_101( .ZN(N574), .A(N406) );
  INV_X1 NOT1_102( .ZN(N575), .A(N419) );
  INV_X2 NOT1_103( .ZN(N576), .A(N432) );
  INV_X2 NOT1_104( .ZN(N577), .A(N406) );
  INV_X1 NOT1_105( .ZN(N578), .A(N419) );
  INV_X1 NOT1_106( .ZN(N579), .A(N445) );
  INV_X1 NOT1_107( .ZN(N580), .A(N406) );
  INV_X1 NOT1_108( .ZN(N581), .A(N432) );
  INV_X1 NOT1_109( .ZN(N582), .A(N445) );
  INV_X1 NOT1_110( .ZN(N583), .A(N419) );
  INV_X1 NOT1_111( .ZN(N584), .A(N432) );
  INV_X1 NOT1_112( .ZN(N585), .A(N445) );
  INV_X1 NOT1_113( .ZN(N586), .A(N367) );
  INV_X1 NOT1_114( .ZN(N587), .A(N393) );
  INV_X1 NOT1_115( .ZN(N588), .A(N367) );
  INV_X1 NOT1_116( .ZN(N589), .A(N380) );
  INV_X1 NOT1_117( .ZN(N590), .A(N354) );
  INV_X1 NOT1_118( .ZN(N591), .A(N393) );
  INV_X1 NOT1_119( .ZN(N592), .A(N354) );
  INV_X1 NOT1_120( .ZN(N593), .A(N380) );
  AND4_X1 AND4_121( .ZN(N594), .A1(N554), .A2(N555), .A3(N556), .A4(N393) );
  AND4_X1 AND4_122( .ZN(N595), .A1(N557), .A2(N558), .A3(N380), .A4(N559) );
  AND4_X1 AND4_123( .ZN(N596), .A1(N560), .A2(N367), .A3(N561), .A4(N562) );
  AND4_X4 AND4_124( .ZN(N597), .A1(N354), .A2(N563), .A3(N564), .A4(N565) );
  AND4_X4 AND4_125( .ZN(N598), .A1(N574), .A2(N575), .A3(N576), .A4(N445) );
  AND4_X1 AND4_126( .ZN(N599), .A1(N577), .A2(N578), .A3(N432), .A4(N579) );
  AND4_X1 AND4_127( .ZN(N600), .A1(N580), .A2(N419), .A3(N581), .A4(N582) );
  AND4_X1 AND4_128( .ZN(N601), .A1(N406), .A2(N583), .A3(N584), .A4(N585) );
  OR4_X1 OR4_129( .ZN(N602), .A1(N594), .A2(N595), .A3(N596), .A4(N597) );
  OR4_X1 OR4_130( .ZN(N607), .A1(N598), .A2(N599), .A3(N600), .A4(N601) );
  AND4_X1 AND5_131_A( .ZN(extra0), .A1(N406), .A2(N566), .A3(N432), .A4(N567) );
  AND2_X1 AND5_131( .ZN(N620), .A1(extra0), .A2(N602) );
  AND4_X1 AND5_132_A( .ZN(extra1), .A1(N406), .A2(N568), .A3(N569), .A4(N445) );
  AND2_X1 AND5_132( .ZN(N625), .A1(extra1), .A2(N602) );
  AND4_X1 AND5_133_A( .ZN(extra2), .A1(N570), .A2(N419), .A3(N432), .A4(N571) );
  AND2_X1 AND5_133( .ZN(N630), .A1(extra2), .A2(N602) );
  AND4_X1 AND5_134_A( .ZN(extra3), .A1(N572), .A2(N419), .A3(N573), .A4(N445) );
  AND2_X1 AND5_134( .ZN(N635), .A1(extra3), .A2(N602) );
  AND4_X1 AND5_135_A( .ZN(extra4), .A1(N354), .A2(N586), .A3(N380), .A4(N587) );
  AND2_X1 AND5_135( .ZN(N640), .A1(extra4), .A2(N607) );
  AND4_X1 AND5_136_A( .ZN(extra5), .A1(N354), .A2(N588), .A3(N589), .A4(N393) );
  AND2_X1 AND5_136( .ZN(N645), .A1(extra5), .A2(N607) );
  AND4_X2 AND5_137_A( .ZN(extra6), .A1(N590), .A2(N367), .A3(N380), .A4(N591) );
  AND2_X2 AND5_137( .ZN(N650), .A1(extra6), .A2(N607) );
  AND4_X4 AND5_138_A( .ZN(extra7), .A1(N592), .A2(N367), .A3(N593), .A4(N393) );
  AND2_X4 AND5_138( .ZN(N655), .A1(extra7), .A2(N607) );
  AND2_X1 AND2_139( .ZN(N692), .A1(N354), .A2(N620) );
  AND2_X1 AND2_140( .ZN(N693), .A1(N367), .A2(N620) );
  AND2_X1 AND2_141( .ZN(N694), .A1(N380), .A2(N620) );
  AND2_X1 AND2_142( .ZN(N695), .A1(N393), .A2(N620) );
  AND2_X1 AND2_143( .ZN(N696), .A1(N354), .A2(N625) );
  AND2_X1 AND2_144( .ZN(N697), .A1(N367), .A2(N625) );
  AND2_X1 AND2_145( .ZN(N698), .A1(N380), .A2(N625) );
  AND2_X1 AND2_146( .ZN(N699), .A1(N393), .A2(N625) );
  AND2_X1 AND2_147( .ZN(N700), .A1(N354), .A2(N630) );
  AND2_X1 AND2_148( .ZN(N701), .A1(N367), .A2(N630) );
  AND2_X1 AND2_149( .ZN(N702), .A1(N380), .A2(N630) );
  AND2_X1 AND2_150( .ZN(N703), .A1(N393), .A2(N630) );
  AND2_X1 AND2_151( .ZN(N704), .A1(N354), .A2(N635) );
  AND2_X1 AND2_152( .ZN(N705), .A1(N367), .A2(N635) );
  AND2_X1 AND2_153( .ZN(N706), .A1(N380), .A2(N635) );
  AND2_X1 AND2_154( .ZN(N707), .A1(N393), .A2(N635) );
  AND2_X1 AND2_155( .ZN(N708), .A1(N406), .A2(N640) );
  AND2_X1 AND2_156( .ZN(N709), .A1(N419), .A2(N640) );
  AND2_X1 AND2_157( .ZN(N710), .A1(N432), .A2(N640) );
  AND2_X1 AND2_158( .ZN(N711), .A1(N445), .A2(N640) );
  AND2_X1 AND2_159( .ZN(N712), .A1(N406), .A2(N645) );
  AND2_X1 AND2_160( .ZN(N713), .A1(N419), .A2(N645) );
  AND2_X2 AND2_161( .ZN(N714), .A1(N432), .A2(N645) );
  AND2_X2 AND2_162( .ZN(N715), .A1(N445), .A2(N645) );
  AND2_X2 AND2_163( .ZN(N716), .A1(N406), .A2(N650) );
  AND2_X2 AND2_164( .ZN(N717), .A1(N419), .A2(N650) );
  AND2_X2 AND2_165( .ZN(N718), .A1(N432), .A2(N650) );
  AND2_X1 AND2_166( .ZN(N719), .A1(N445), .A2(N650) );
  AND2_X1 AND2_167( .ZN(N720), .A1(N406), .A2(N655) );
  AND2_X1 AND2_168( .ZN(N721), .A1(N419), .A2(N655) );
  AND2_X1 AND2_169( .ZN(N722), .A1(N432), .A2(N655) );
  AND2_X1 AND2_170( .ZN(N723), .A1(N445), .A2(N655) );
  XOR2_X1 XOR2_171( .Z(N724), .A(N1), .B(N692) );
  XOR2_X1 XOR2_172( .Z(N725), .A(N5), .B(N693) );
  XOR2_X1 XOR2_173( .Z(N726), .A(N9), .B(N694) );
  XOR2_X1 XOR2_174( .Z(N727), .A(N13), .B(N695) );
  XOR2_X1 XOR2_175( .Z(N728), .A(N17), .B(N696) );
  XOR2_X1 XOR2_176( .Z(N729), .A(N21), .B(N697) );
  XOR2_X1 XOR2_177( .Z(N730), .A(N25), .B(N698) );
  XOR2_X1 XOR2_178( .Z(N731), .A(N29), .B(N699) );
  XOR2_X1 XOR2_179( .Z(N732), .A(N33), .B(N700) );
  XOR2_X1 XOR2_180( .Z(N733), .A(N37), .B(N701) );
  XOR2_X1 XOR2_181( .Z(N734), .A(N41), .B(N702) );
  XOR2_X1 XOR2_182( .Z(N735), .A(N45), .B(N703) );
  XOR2_X1 XOR2_183( .Z(N736), .A(N49), .B(N704) );
  XOR2_X1 XOR2_184( .Z(N737), .A(N53), .B(N705) );
  XOR2_X1 XOR2_185( .Z(N738), .A(N57), .B(N706) );
  XOR2_X1 XOR2_186( .Z(N739), .A(N61), .B(N707) );
  XOR2_X1 XOR2_187( .Z(N740), .A(N65), .B(N708) );
  XOR2_X1 XOR2_188( .Z(N741), .A(N69), .B(N709) );
  XOR2_X1 XOR2_189( .Z(N742), .A(N73), .B(N710) );
  XOR2_X2 XOR2_190( .Z(N743), .A(N77), .B(N711) );
  XOR2_X2 XOR2_191( .Z(N744), .A(N81), .B(N712) );
  XOR2_X1 XOR2_192( .Z(N745), .A(N85), .B(N713) );
  XOR2_X1 XOR2_193( .Z(N746), .A(N89), .B(N714) );
  XOR2_X1 XOR2_194( .Z(N747), .A(N93), .B(N715) );
  XOR2_X1 XOR2_195( .Z(N748), .A(N97), .B(N716) );
  XOR2_X1 XOR2_196( .Z(N749), .A(N101), .B(N717) );
  XOR2_X1 XOR2_197( .Z(N750), .A(N105), .B(N718) );
  XOR2_X1 XOR2_198( .Z(N751), .A(N109), .B(N719) );
  XOR2_X1 XOR2_199( .Z(N752), .A(N113), .B(N720) );
  XOR2_X1 XOR2_200( .Z(N753), .A(N117), .B(N721) );
  XOR2_X1 XOR2_201( .Z(N754), .A(N121), .B(N722) );
  XOR2_X1 XOR2_202( .Z(N755), .A(N125), .B(N723) );

endmodule
