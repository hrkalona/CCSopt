// Verilog
// c6288
// Ninputs 32
// Noutputs 32
// NtotalGates 2416
// AND2 256
// NOT1 32
// NOR2 2128

module c6288(N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,
  N307,N324,N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528,N545,N1581,N1901,N2223,
  N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,N6190,N6200,
  N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288);
input N1,N18,N35,N52,N69,N86,N103,N120,N137,N154,N171,N188,N205,N222,N239,N256,N273,N290,N307,N324,
  N341,N358,N375,N392,N409,N426,N443,N460,N477,N494,N511,N528;
output N545,N1581,N1901,N2223,N2548,N2877,N3211,N3552,N3895,N4241,N4591,N4946,N5308,N5672,N5971,N6123,N6150,N6160,N6170,N6180,
  N6190,N6200,N6210,N6220,N6230,N6240,N6250,N6260,N6270,N6280,N6287,N6288;

  wire N546,N549,N552,N555,N558,N561,N564,N567,N570,N573,N576,N579,N582,N585,N588,N591,
    N594,N597,N600,N603,N606,N609,N612,N615,N618,N621,N624,N627,N630,N633,N636,N639,
    N642,N645,N648,N651,N654,N657,N660,N663,N666,N669,N672,N675,N678,N681,N684,N687,
    N690,N693,N696,N699,N702,N705,N708,N711,N714,N717,N720,N723,N726,N729,N732,N735,
    N738,N741,N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,
    N786,N789,N792,N795,N798,N801,N804,N807,N810,N813,N816,N819,N822,N825,N828,N831,
    N834,N837,N840,N843,N846,N849,N852,N855,N858,N861,N864,N867,N870,N873,N876,N879,
    N882,N885,N888,N891,N894,N897,N900,N903,N906,N909,N912,N915,N918,N921,N924,N927,
    N930,N933,N936,N939,N942,N945,N948,N951,N954,N957,N960,N963,N966,N969,N972,N975,
    N978,N981,N984,N987,N990,N993,N996,N999,N1002,N1005,N1008,N1011,N1014,N1017,N1020,N1023,
    N1026,N1029,N1032,N1035,N1038,N1041,N1044,N1047,N1050,N1053,N1056,N1059,N1062,N1065,N1068,N1071,
    N1074,N1077,N1080,N1083,N1086,N1089,N1092,N1095,N1098,N1101,N1104,N1107,N1110,N1113,N1116,N1119,
    N1122,N1125,N1128,N1131,N1134,N1137,N1140,N1143,N1146,N1149,N1152,N1155,N1158,N1161,N1164,N1167,
    N1170,N1173,N1176,N1179,N1182,N1185,N1188,N1191,N1194,N1197,N1200,N1203,N1206,N1209,N1212,N1215,
    N1218,N1221,N1224,N1227,N1230,N1233,N1236,N1239,N1242,N1245,N1248,N1251,N1254,N1257,N1260,N1263,
    N1266,N1269,N1272,N1275,N1278,N1281,N1284,N1287,N1290,N1293,N1296,N1299,N1302,N1305,N1308,N1311,
    N1315,N1319,N1323,N1327,N1331,N1335,N1339,N1343,N1347,N1351,N1355,N1359,N1363,N1367,N1371,N1372,
    N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
    N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1404,N1407,N1410,
    N1413,N1416,N1419,N1422,N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1450,N1454,N1458,N1462,
    N1466,N1470,N1474,N1478,N1482,N1486,N1490,N1494,N1498,N1502,N1506,N1507,N1508,N1511,N1512,N1513,
    N1516,N1517,N1518,N1521,N1522,N1523,N1526,N1527,N1528,N1531,N1532,N1533,N1536,N1537,N1538,N1541,
    N1542,N1543,N1546,N1547,N1548,N1551,N1552,N1553,N1556,N1557,N1558,N1561,N1562,N1563,N1566,N1567,
    N1568,N1571,N1572,N1573,N1576,N1577,N1578,N1582,N1585,N1588,N1591,N1594,N1597,N1600,N1603,N1606,
    N1609,N1612,N1615,N1618,N1621,N1624,N1628,N1632,N1636,N1640,N1644,N1648,N1652,N1656,N1660,N1664,
    N1668,N1672,N1676,N1680,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,
    N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,
    N1712,N1713,N1714,N1717,N1720,N1723,N1726,N1729,N1732,N1735,N1738,N1741,N1744,N1747,N1750,N1753,
    N1756,N1759,N1763,N1767,N1771,N1775,N1779,N1783,N1787,N1791,N1795,N1799,N1803,N1807,N1811,N1815,
    N1819,N1820,N1821,N1824,N1825,N1826,N1829,N1830,N1831,N1834,N1835,N1836,N1839,N1840,N1841,N1844,
    N1845,N1846,N1849,N1850,N1851,N1854,N1855,N1856,N1859,N1860,N1861,N1864,N1865,N1866,N1869,N1870,
    N1871,N1874,N1875,N1876,N1879,N1880,N1881,N1884,N1885,N1886,N1889,N1890,N1891,N1894,N1897,N1902,
    N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,N1932,N1935,N1938,N1941,N1945,N1946,N1947,
    N1951,N1955,N1959,N1963,N1967,N1971,N1975,N1979,N1983,N1987,N1991,N1995,N1999,N2000,N2001,N2004,
    N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,
    N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2033,N2037,N2040,N2043,N2046,N2049,
    N2052,N2055,N2058,N2061,N2064,N2067,N2070,N2073,N2076,N2080,N2081,N2082,N2085,N2089,N2093,N2097,
    N2101,N2105,N2109,N2113,N2117,N2121,N2125,N2129,N2133,N2137,N2138,N2139,N2142,N2145,N2149,N2150,
    N2151,N2154,N2155,N2156,N2159,N2160,N2161,N2164,N2165,N2166,N2169,N2170,N2171,N2174,N2175,N2176,
    N2179,N2180,N2181,N2184,N2185,N2186,N2189,N2190,N2191,N2194,N2195,N2196,N2199,N2200,N2201,N2204,
    N2205,N2206,N2209,N2210,N2211,N2214,N2217,N2221,N2222,N2224,N2227,N2230,N2233,N2236,N2239,N2242,
    N2245,N2248,N2251,N2254,N2257,N2260,N2264,N2265,N2266,N2269,N2273,N2277,N2281,N2285,N2289,N2293,
    N2297,N2301,N2305,N2309,N2313,N2317,N2318,N2319,N2322,N2326,N2327,N2328,N2329,N2330,N2331,N2332,
    N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,
    N2349,N2350,N2353,N2357,N2358,N2359,N2362,N2365,N2368,N2371,N2374,N2377,N2380,N2383,N2386,N2389,
    N2392,N2395,N2398,N2402,N2403,N2404,N2407,N2410,N2414,N2418,N2422,N2426,N2430,N2434,N2438,N2442,
    N2446,N2450,N2454,N2458,N2462,N2463,N2464,N2467,N2470,N2474,N2475,N2476,N2477,N2478,N2481,N2482,
    N2483,N2486,N2487,N2488,N2491,N2492,N2493,N2496,N2497,N2498,N2501,N2502,N2503,N2506,N2507,N2508,
    N2511,N2512,N2513,N2516,N2517,N2518,N2521,N2522,N2523,N2526,N2527,N2528,N2531,N2532,N2533,N2536,
    N2539,N2543,N2544,N2545,N2549,N2552,N2555,N2558,N2561,N2564,N2567,N2570,N2573,N2576,N2579,N2582,
    N2586,N2587,N2588,N2591,N2595,N2599,N2603,N2607,N2611,N2615,N2619,N2623,N2627,N2631,N2635,N2639,
    N2640,N2641,N2644,N2648,N2649,N2650,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,
    N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2678,N2682,N2683,
    N2684,N2687,N2690,N2694,N2697,N2700,N2703,N2706,N2709,N2712,N2715,N2718,N2721,N2724,N2727,N2731,
    N2732,N2733,N2736,N2739,N2743,N2744,N2745,N2749,N2753,N2757,N2761,N2765,N2769,N2773,N2777,N2781,
    N2785,N2789,N2790,N2791,N2794,N2797,N2801,N2802,N2803,N2806,N2807,N2808,N2811,N2812,N2813,N2816,
    N2817,N2818,N2821,N2822,N2823,N2826,N2827,N2828,N2831,N2832,N2833,N2836,N2837,N2838,N2841,N2842,
    N2843,N2846,N2847,N2848,N2851,N2852,N2853,N2856,N2857,N2858,N2861,N2864,N2868,N2869,N2870,N2873,
    N2878,N2881,N2884,N2887,N2890,N2893,N2896,N2899,N2902,N2905,N2908,N2912,N2913,N2914,N2917,N2921,
    N2922,N2923,N2926,N2930,N2934,N2938,N2942,N2946,N2950,N2954,N2958,N2962,N2966,N2967,N2968,N2971,
    N2975,N2976,N2977,N2980,N2983,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
    N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3010,N3014,N3015,N3016,N3019,N3022,
    N3026,N3027,N3028,N3031,N3034,N3037,N3040,N3043,N3046,N3049,N3052,N3055,N3058,N3062,N3063,N3064,
    N3067,N3070,N3074,N3075,N3076,N3079,N3083,N3087,N3091,N3095,N3099,N3103,N3107,N3111,N3115,N3119,
    N3120,N3121,N3124,N3127,N3131,N3132,N3133,N3136,N3140,N3141,N3142,N3145,N3146,N3147,N3150,N3151,
    N3152,N3155,N3156,N3157,N3160,N3161,N3162,N3165,N3166,N3167,N3170,N3171,N3172,N3175,N3176,N3177,
    N3180,N3181,N3182,N3185,N3186,N3187,N3190,N3193,N3197,N3198,N3199,N3202,N3206,N3207,N3208,N3212,
    N3215,N3218,N3221,N3224,N3227,N3230,N3233,N3236,N3239,N3243,N3244,N3245,N3248,N3252,N3253,N3254,
    N3257,N3260,N3264,N3268,N3272,N3276,N3280,N3284,N3288,N3292,N3296,N3300,N3301,N3302,N3305,N3309,
    N3310,N3311,N3314,N3317,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,
    N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3344,N3348,N3349,N3350,N3353,N3356,N3360,
    N3361,N3362,N3365,N3368,N3371,N3374,N3377,N3380,N3383,N3386,N3389,N3392,N3396,N3397,N3398,N3401,
    N3404,N3408,N3409,N3410,N3413,N3417,N3421,N3425,N3429,N3433,N3437,N3441,N3445,N3449,N3453,N3454,
    N3455,N3458,N3461,N3465,N3466,N3467,N3470,N3474,N3475,N3476,N3479,N3480,N3481,N3484,N3485,N3486,
    N3489,N3490,N3491,N3494,N3495,N3496,N3499,N3500,N3501,N3504,N3505,N3506,N3509,N3510,N3511,N3514,
    N3515,N3516,N3519,N3520,N3521,N3524,N3527,N3531,N3532,N3533,N3536,N3540,N3541,N3542,N3545,N3548,
    N3553,N3556,N3559,N3562,N3565,N3568,N3571,N3574,N3577,N3581,N3582,N3583,N3586,N3590,N3591,N3592,
    N3595,N3598,N3602,N3603,N3604,N3608,N3612,N3616,N3620,N3624,N3628,N3632,N3636,N3637,N3638,N3641,
    N3645,N3646,N3647,N3650,N3653,N3657,N3658,N3659,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,
    N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3681,N3685,N3686,N3687,N3690,N3693,N3697,
    N3698,N3699,N3702,N3706,N3709,N3712,N3715,N3718,N3721,N3724,N3727,N3730,N3734,N3735,N3736,N3739,
    N3742,N3746,N3747,N3748,N3751,N3755,N3756,N3757,N3760,N3764,N3768,N3772,N3776,N3780,N3784,N3788,
    N3792,N3793,N3794,N3797,N3800,N3804,N3805,N3806,N3809,N3813,N3814,N3815,N3818,N3821,N3825,N3826,
    N3827,N3830,N3831,N3832,N3835,N3836,N3837,N3840,N3841,N3842,N3845,N3846,N3847,N3850,N3851,N3852,
    N3855,N3856,N3857,N3860,N3861,N3862,N3865,N3868,N3872,N3873,N3874,N3877,N3881,N3882,N3883,N3886,
    N3889,N3893,N3894,N3896,N3899,N3902,N3905,N3908,N3911,N3914,N3917,N3921,N3922,N3923,N3926,N3930,
    N3931,N3932,N3935,N3938,N3942,N3943,N3944,N3947,N3951,N3955,N3959,N3963,N3967,N3971,N3975,N3976,
    N3977,N3980,N3984,N3985,N3986,N3989,N3992,N3996,N3997,N3998,N4001,N4005,N4006,N4007,N4008,N4009,
    N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4022,N4026,N4027,N4028,N4031,N4034,
    N4038,N4039,N4040,N4043,N4047,N4048,N4049,N4052,N4055,N4058,N4061,N4064,N4067,N4070,N4073,N4077,
    N4078,N4079,N4082,N4085,N4089,N4090,N4091,N4094,N4098,N4099,N4100,N4103,N4106,N4110,N4114,N4118,
    N4122,N4126,N4130,N4134,N4138,N4139,N4140,N4143,N4146,N4150,N4151,N4152,N4155,N4159,N4160,N4161,
    N4164,N4167,N4171,N4172,N4173,N4174,N4175,N4178,N4179,N4180,N4183,N4184,N4185,N4188,N4189,N4190,
    N4193,N4194,N4195,N4198,N4199,N4200,N4203,N4204,N4205,N4208,N4211,N4215,N4216,N4217,N4220,N4224,
    N4225,N4226,N4229,N4232,N4236,N4237,N4238,N4242,N4245,N4248,N4251,N4254,N4257,N4260,N4264,N4265,
    N4266,N4269,N4273,N4274,N4275,N4278,N4281,N4285,N4286,N4287,N4290,N4294,N4298,N4302,N4306,N4310,
    N4314,N4318,N4319,N4320,N4323,N4327,N4328,N4329,N4332,N4335,N4339,N4340,N4341,N4344,N4348,N4349,
    N4350,N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4368,N4372,
    N4373,N4374,N4377,N4380,N4384,N4385,N4386,N4389,N4393,N4394,N4395,N4398,N4401,N4405,N4408,N4411,
    N4414,N4417,N4420,N4423,N4427,N4428,N4429,N4432,N4435,N4439,N4440,N4441,N4444,N4448,N4449,N4450,
    N4453,N4456,N4460,N4461,N4462,N4466,N4470,N4474,N4478,N4482,N4486,N4487,N4488,N4491,N4494,N4498,
    N4499,N4500,N4503,N4507,N4508,N4509,N4512,N4515,N4519,N4520,N4521,N4524,N4525,N4526,N4529,N4530,
    N4531,N4534,N4535,N4536,N4539,N4540,N4541,N4544,N4545,N4546,N4549,N4550,N4551,N4554,N4557,N4561,
    N4562,N4563,N4566,N4570,N4571,N4572,N4575,N4578,N4582,N4583,N4584,N4587,N4592,N4595,N4598,N4601,
    N4604,N4607,N4611,N4612,N4613,N4616,N4620,N4621,N4622,N4625,N4628,N4632,N4633,N4634,N4637,N4641,
    N4642,N4643,N4646,N4650,N4654,N4658,N4662,N4666,N4667,N4668,N4671,N4675,N4676,N4677,N4680,N4683,
    N4687,N4688,N4689,N4692,N4696,N4697,N4698,N4701,N4704,N4708,N4709,N4710,N4711,N4712,N4713,N4714,
    N4715,N4716,N4717,N4718,N4721,N4725,N4726,N4727,N4730,N4733,N4737,N4738,N4739,N4742,N4746,N4747,
    N4748,N4751,N4754,N4758,N4759,N4760,N4763,N4766,N4769,N4772,N4775,N4779,N4780,N4781,N4784,N4787,
    N4791,N4792,N4793,N4796,N4800,N4801,N4802,N4805,N4808,N4812,N4813,N4814,N4817,N4821,N4825,N4829,
    N4833,N4837,N4838,N4839,N4842,N4845,N4849,N4850,N4851,N4854,N4858,N4859,N4860,N4863,N4866,N4870,
    N4871,N4872,N4875,N4879,N4880,N4881,N4884,N4885,N4886,N4889,N4890,N4891,N4894,N4895,N4896,N4899,
    N4900,N4901,N4904,N4907,N4911,N4912,N4913,N4916,N4920,N4921,N4922,N4925,N4928,N4932,N4933,N4934,
    N4937,N4941,N4942,N4943,N4947,N4950,N4953,N4956,N4959,N4963,N4964,N4965,N4968,N4972,N4973,N4974,
    N4977,N4980,N4984,N4985,N4986,N4989,N4993,N4994,N4995,N4998,N5001,N5005,N5009,N5013,N5017,N5021,
    N5022,N5023,N5026,N5030,N5031,N5032,N5035,N5038,N5042,N5043,N5044,N5047,N5051,N5052,N5053,N5056,
    N5059,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5076,N5080,N5081,N5082,
    N5085,N5088,N5092,N5093,N5094,N5097,N5101,N5102,N5103,N5106,N5109,N5113,N5114,N5115,N5118,N5121,
    N5124,N5127,N5130,N5134,N5135,N5136,N5139,N5142,N5146,N5147,N5148,N5151,N5155,N5156,N5157,N5160,
    N5163,N5167,N5168,N5169,N5172,N5176,N5180,N5184,N5188,N5192,N5193,N5194,N5197,N5200,N5204,N5205,
    N5206,N5209,N5213,N5214,N5215,N5218,N5221,N5225,N5226,N5227,N5230,N5234,N5235,N5236,N5239,N5240,
    N5241,N5244,N5245,N5246,N5249,N5250,N5251,N5254,N5255,N5256,N5259,N5262,N5266,N5267,N5268,N5271,
    N5275,N5276,N5277,N5280,N5283,N5287,N5288,N5289,N5292,N5296,N5297,N5298,N5301,N5304,N5309,N5312,
    N5315,N5318,N5322,N5323,N5324,N5327,N5331,N5332,N5333,N5336,N5339,N5343,N5344,N5345,N5348,N5352,
    N5353,N5354,N5357,N5360,N5364,N5365,N5366,N5370,N5374,N5378,N5379,N5380,N5383,N5387,N5388,N5389,
    N5392,N5395,N5399,N5400,N5401,N5404,N5408,N5409,N5410,N5413,N5416,N5420,N5421,N5422,N5425,N5426,
    N5427,N5428,N5429,N5430,N5431,N5434,N5438,N5439,N5440,N5443,N5446,N5450,N5451,N5452,N5455,N5459,
    N5460,N5461,N5464,N5467,N5471,N5472,N5473,N5476,N5480,N5483,N5486,N5489,N5493,N5494,N5495,N5498,
    N5501,N5505,N5506,N5507,N5510,N5514,N5515,N5516,N5519,N5522,N5526,N5527,N5528,N5531,N5535,N5536,
    N5537,N5540,N5544,N5548,N5552,N5553,N5554,N5557,N5560,N5564,N5565,N5566,N5569,N5573,N5574,N5575,
    N5578,N5581,N5585,N5586,N5587,N5590,N5594,N5595,N5596,N5599,N5602,N5606,N5607,N5608,N5611,N5612,
    N5613,N5616,N5617,N5618,N5621,N5624,N5628,N5629,N5630,N5633,N5637,N5638,N5639,N5642,N5645,N5649,
    N5650,N5651,N5654,N5658,N5659,N5660,N5663,N5666,N5670,N5671,N5673,N5676,N5679,N5683,N5684,N5685,
    N5688,N5692,N5693,N5694,N5697,N5700,N5704,N5705,N5706,N5709,N5713,N5714,N5715,N5718,N5721,N5725,
    N5726,N5727,N5730,N5734,N5738,N5739,N5740,N5743,N5747,N5748,N5749,N5752,N5755,N5759,N5760,N5761,
    N5764,N5768,N5769,N5770,N5773,N5776,N5780,N5781,N5782,N5785,N5786,N5787,N5788,N5789,N5792,N5796,
    N5797,N5798,N5801,N5804,N5808,N5809,N5810,N5813,N5817,N5818,N5819,N5822,N5825,N5829,N5830,N5831,
    N5834,N5837,N5840,N5844,N5845,N5846,N5849,N5852,N5856,N5857,N5858,N5861,N5865,N5866,N5867,N5870,
    N5873,N5877,N5878,N5879,N5882,N5886,N5890,N5891,N5892,N5895,N5898,N5902,N5903,N5904,N5907,N5911,
    N5912,N5913,N5916,N5919,N5923,N5924,N5925,N5928,N5929,N5930,N5933,N5934,N5935,N5938,N5941,N5945,
    N5946,N5947,N5950,N5954,N5955,N5956,N5959,N5962,N5966,N5967,N5968,N5972,N5975,N5979,N5980,N5981,
    N5984,N5988,N5989,N5990,N5993,N5996,N6000,N6001,N6002,N6005,N6009,N6010,N6011,N6014,N6018,N6019,
    N6020,N6023,N6026,N6030,N6031,N6032,N6035,N6036,N6037,N6040,N6044,N6045,N6046,N6049,N6052,N6056,
    N6057,N6058,N6061,N6064,N6068,N6069,N6070,N6073,N6076,N6080,N6081,N6082,N6085,N6089,N6090,N6091,
    N6094,N6097,N6101,N6102,N6103,N6106,N6107,N6108,N6111,N6114,N6118,N6119,N6120,N6124,N6128,N6129,
    N6130,N6133,N6134,N6135,N6138,N6141,N6145,N6146,N6147,N6151,N6155,N6156,N6157,N6161,N6165,N6166,
    N6167,N6171,N6175,N6176,N6177,N6181,N6185,N6186,N6187,N6191,N6195,N6196,N6197,N6201,N6205,N6206,
    N6207,N6211,N6215,N6216,N6217,N6221,N6225,N6226,N6227,N6231,N6235,N6236,N6237,N6241,N6245,N6246,
    N6247,N6251,N6255,N6256,N6257,N6261,N6265,N6266,N6267,N6271,N6275,N6276,N6277,N6281,N6285,N6286;

  AND2_X1 AND2_1( .ZN(N545), .A1(N1), .A2(N273) );
  AND2_X2 AND2_2( .ZN(N546), .A1(N1), .A2(N290) );
  AND2_X2 AND2_3( .ZN(N549), .A1(N1), .A2(N307) );
  AND2_X2 AND2_4( .ZN(N552), .A1(N1), .A2(N324) );
  AND2_X2 AND2_5( .ZN(N555), .A1(N1), .A2(N341) );
  AND2_X2 AND2_6( .ZN(N558), .A1(N1), .A2(N358) );
  AND2_X1 AND2_7( .ZN(N561), .A1(N1), .A2(N375) );
  AND2_X1 AND2_8( .ZN(N564), .A1(N1), .A2(N392) );
  AND2_X1 AND2_9( .ZN(N567), .A1(N1), .A2(N409) );
  AND2_X1 AND2_10( .ZN(N570), .A1(N1), .A2(N426) );
  AND2_X1 AND2_11( .ZN(N573), .A1(N1), .A2(N443) );
  AND2_X1 AND2_12( .ZN(N576), .A1(N1), .A2(N460) );
  AND2_X1 AND2_13( .ZN(N579), .A1(N1), .A2(N477) );
  AND2_X1 AND2_14( .ZN(N582), .A1(N1), .A2(N494) );
  AND2_X1 AND2_15( .ZN(N585), .A1(N1), .A2(N511) );
  AND2_X1 AND2_16( .ZN(N588), .A1(N1), .A2(N528) );
  AND2_X1 AND2_17( .ZN(N591), .A1(N18), .A2(N273) );
  AND2_X1 AND2_18( .ZN(N594), .A1(N18), .A2(N290) );
  AND2_X1 AND2_19( .ZN(N597), .A1(N18), .A2(N307) );
  AND2_X1 AND2_20( .ZN(N600), .A1(N18), .A2(N324) );
  AND2_X1 AND2_21( .ZN(N603), .A1(N18), .A2(N341) );
  AND2_X1 AND2_22( .ZN(N606), .A1(N18), .A2(N358) );
  AND2_X1 AND2_23( .ZN(N609), .A1(N18), .A2(N375) );
  AND2_X1 AND2_24( .ZN(N612), .A1(N18), .A2(N392) );
  AND2_X1 AND2_25( .ZN(N615), .A1(N18), .A2(N409) );
  AND2_X1 AND2_26( .ZN(N618), .A1(N18), .A2(N426) );
  AND2_X1 AND2_27( .ZN(N621), .A1(N18), .A2(N443) );
  AND2_X1 AND2_28( .ZN(N624), .A1(N18), .A2(N460) );
  AND2_X1 AND2_29( .ZN(N627), .A1(N18), .A2(N477) );
  AND2_X1 AND2_30( .ZN(N630), .A1(N18), .A2(N494) );
  AND2_X1 AND2_31( .ZN(N633), .A1(N18), .A2(N511) );
  AND2_X1 AND2_32( .ZN(N636), .A1(N18), .A2(N528) );
  AND2_X1 AND2_33( .ZN(N639), .A1(N35), .A2(N273) );
  AND2_X1 AND2_34( .ZN(N642), .A1(N35), .A2(N290) );
  AND2_X1 AND2_35( .ZN(N645), .A1(N35), .A2(N307) );
  AND2_X1 AND2_36( .ZN(N648), .A1(N35), .A2(N324) );
  AND2_X1 AND2_37( .ZN(N651), .A1(N35), .A2(N341) );
  AND2_X1 AND2_38( .ZN(N654), .A1(N35), .A2(N358) );
  AND2_X1 AND2_39( .ZN(N657), .A1(N35), .A2(N375) );
  AND2_X1 AND2_40( .ZN(N660), .A1(N35), .A2(N392) );
  AND2_X1 AND2_41( .ZN(N663), .A1(N35), .A2(N409) );
  AND2_X1 AND2_42( .ZN(N666), .A1(N35), .A2(N426) );
  AND2_X1 AND2_43( .ZN(N669), .A1(N35), .A2(N443) );
  AND2_X1 AND2_44( .ZN(N672), .A1(N35), .A2(N460) );
  AND2_X1 AND2_45( .ZN(N675), .A1(N35), .A2(N477) );
  AND2_X1 AND2_46( .ZN(N678), .A1(N35), .A2(N494) );
  AND2_X1 AND2_47( .ZN(N681), .A1(N35), .A2(N511) );
  AND2_X1 AND2_48( .ZN(N684), .A1(N35), .A2(N528) );
  AND2_X1 AND2_49( .ZN(N687), .A1(N52), .A2(N273) );
  AND2_X1 AND2_50( .ZN(N690), .A1(N52), .A2(N290) );
  AND2_X1 AND2_51( .ZN(N693), .A1(N52), .A2(N307) );
  AND2_X1 AND2_52( .ZN(N696), .A1(N52), .A2(N324) );
  AND2_X1 AND2_53( .ZN(N699), .A1(N52), .A2(N341) );
  AND2_X1 AND2_54( .ZN(N702), .A1(N52), .A2(N358) );
  AND2_X1 AND2_55( .ZN(N705), .A1(N52), .A2(N375) );
  AND2_X1 AND2_56( .ZN(N708), .A1(N52), .A2(N392) );
  AND2_X1 AND2_57( .ZN(N711), .A1(N52), .A2(N409) );
  AND2_X1 AND2_58( .ZN(N714), .A1(N52), .A2(N426) );
  AND2_X2 AND2_59( .ZN(N717), .A1(N52), .A2(N443) );
  AND2_X2 AND2_60( .ZN(N720), .A1(N52), .A2(N460) );
  AND2_X2 AND2_61( .ZN(N723), .A1(N52), .A2(N477) );
  AND2_X2 AND2_62( .ZN(N726), .A1(N52), .A2(N494) );
  AND2_X2 AND2_63( .ZN(N729), .A1(N52), .A2(N511) );
  AND2_X2 AND2_64( .ZN(N732), .A1(N52), .A2(N528) );
  AND2_X1 AND2_65( .ZN(N735), .A1(N69), .A2(N273) );
  AND2_X1 AND2_66( .ZN(N738), .A1(N69), .A2(N290) );
  AND2_X1 AND2_67( .ZN(N741), .A1(N69), .A2(N307) );
  AND2_X1 AND2_68( .ZN(N744), .A1(N69), .A2(N324) );
  AND2_X1 AND2_69( .ZN(N747), .A1(N69), .A2(N341) );
  AND2_X1 AND2_70( .ZN(N750), .A1(N69), .A2(N358) );
  AND2_X1 AND2_71( .ZN(N753), .A1(N69), .A2(N375) );
  AND2_X1 AND2_72( .ZN(N756), .A1(N69), .A2(N392) );
  AND2_X1 AND2_73( .ZN(N759), .A1(N69), .A2(N409) );
  AND2_X1 AND2_74( .ZN(N762), .A1(N69), .A2(N426) );
  AND2_X1 AND2_75( .ZN(N765), .A1(N69), .A2(N443) );
  AND2_X1 AND2_76( .ZN(N768), .A1(N69), .A2(N460) );
  AND2_X1 AND2_77( .ZN(N771), .A1(N69), .A2(N477) );
  AND2_X1 AND2_78( .ZN(N774), .A1(N69), .A2(N494) );
  AND2_X1 AND2_79( .ZN(N777), .A1(N69), .A2(N511) );
  AND2_X1 AND2_80( .ZN(N780), .A1(N69), .A2(N528) );
  AND2_X1 AND2_81( .ZN(N783), .A1(N86), .A2(N273) );
  AND2_X1 AND2_82( .ZN(N786), .A1(N86), .A2(N290) );
  AND2_X1 AND2_83( .ZN(N789), .A1(N86), .A2(N307) );
  AND2_X1 AND2_84( .ZN(N792), .A1(N86), .A2(N324) );
  AND2_X1 AND2_85( .ZN(N795), .A1(N86), .A2(N341) );
  AND2_X1 AND2_86( .ZN(N798), .A1(N86), .A2(N358) );
  AND2_X1 AND2_87( .ZN(N801), .A1(N86), .A2(N375) );
  AND2_X1 AND2_88( .ZN(N804), .A1(N86), .A2(N392) );
  AND2_X1 AND2_89( .ZN(N807), .A1(N86), .A2(N409) );
  AND2_X1 AND2_90( .ZN(N810), .A1(N86), .A2(N426) );
  AND2_X1 AND2_91( .ZN(N813), .A1(N86), .A2(N443) );
  AND2_X1 AND2_92( .ZN(N816), .A1(N86), .A2(N460) );
  AND2_X1 AND2_93( .ZN(N819), .A1(N86), .A2(N477) );
  AND2_X1 AND2_94( .ZN(N822), .A1(N86), .A2(N494) );
  AND2_X1 AND2_95( .ZN(N825), .A1(N86), .A2(N511) );
  AND2_X1 AND2_96( .ZN(N828), .A1(N86), .A2(N528) );
  AND2_X1 AND2_97( .ZN(N831), .A1(N103), .A2(N273) );
  AND2_X1 AND2_98( .ZN(N834), .A1(N103), .A2(N290) );
  AND2_X1 AND2_99( .ZN(N837), .A1(N103), .A2(N307) );
  AND2_X1 AND2_100( .ZN(N840), .A1(N103), .A2(N324) );
  AND2_X1 AND2_101( .ZN(N843), .A1(N103), .A2(N341) );
  AND2_X1 AND2_102( .ZN(N846), .A1(N103), .A2(N358) );
  AND2_X1 AND2_103( .ZN(N849), .A1(N103), .A2(N375) );
  AND2_X1 AND2_104( .ZN(N852), .A1(N103), .A2(N392) );
  AND2_X1 AND2_105( .ZN(N855), .A1(N103), .A2(N409) );
  AND2_X1 AND2_106( .ZN(N858), .A1(N103), .A2(N426) );
  AND2_X1 AND2_107( .ZN(N861), .A1(N103), .A2(N443) );
  AND2_X1 AND2_108( .ZN(N864), .A1(N103), .A2(N460) );
  AND2_X1 AND2_109( .ZN(N867), .A1(N103), .A2(N477) );
  AND2_X1 AND2_110( .ZN(N870), .A1(N103), .A2(N494) );
  AND2_X1 AND2_111( .ZN(N873), .A1(N103), .A2(N511) );
  AND2_X1 AND2_112( .ZN(N876), .A1(N103), .A2(N528) );
  AND2_X1 AND2_113( .ZN(N879), .A1(N120), .A2(N273) );
  AND2_X1 AND2_114( .ZN(N882), .A1(N120), .A2(N290) );
  AND2_X1 AND2_115( .ZN(N885), .A1(N120), .A2(N307) );
  AND2_X1 AND2_116( .ZN(N888), .A1(N120), .A2(N324) );
  AND2_X1 AND2_117( .ZN(N891), .A1(N120), .A2(N341) );
  AND2_X1 AND2_118( .ZN(N894), .A1(N120), .A2(N358) );
  AND2_X1 AND2_119( .ZN(N897), .A1(N120), .A2(N375) );
  AND2_X1 AND2_120( .ZN(N900), .A1(N120), .A2(N392) );
  AND2_X1 AND2_121( .ZN(N903), .A1(N120), .A2(N409) );
  AND2_X1 AND2_122( .ZN(N906), .A1(N120), .A2(N426) );
  AND2_X1 AND2_123( .ZN(N909), .A1(N120), .A2(N443) );
  AND2_X1 AND2_124( .ZN(N912), .A1(N120), .A2(N460) );
  AND2_X1 AND2_125( .ZN(N915), .A1(N120), .A2(N477) );
  AND2_X1 AND2_126( .ZN(N918), .A1(N120), .A2(N494) );
  AND2_X1 AND2_127( .ZN(N921), .A1(N120), .A2(N511) );
  AND2_X1 AND2_128( .ZN(N924), .A1(N120), .A2(N528) );
  AND2_X1 AND2_129( .ZN(N927), .A1(N137), .A2(N273) );
  AND2_X1 AND2_130( .ZN(N930), .A1(N137), .A2(N290) );
  AND2_X1 AND2_131( .ZN(N933), .A1(N137), .A2(N307) );
  AND2_X1 AND2_132( .ZN(N936), .A1(N137), .A2(N324) );
  AND2_X1 AND2_133( .ZN(N939), .A1(N137), .A2(N341) );
  AND2_X1 AND2_134( .ZN(N942), .A1(N137), .A2(N358) );
  AND2_X1 AND2_135( .ZN(N945), .A1(N137), .A2(N375) );
  AND2_X1 AND2_136( .ZN(N948), .A1(N137), .A2(N392) );
  AND2_X1 AND2_137( .ZN(N951), .A1(N137), .A2(N409) );
  AND2_X1 AND2_138( .ZN(N954), .A1(N137), .A2(N426) );
  AND2_X1 AND2_139( .ZN(N957), .A1(N137), .A2(N443) );
  AND2_X1 AND2_140( .ZN(N960), .A1(N137), .A2(N460) );
  AND2_X1 AND2_141( .ZN(N963), .A1(N137), .A2(N477) );
  AND2_X1 AND2_142( .ZN(N966), .A1(N137), .A2(N494) );
  AND2_X1 AND2_143( .ZN(N969), .A1(N137), .A2(N511) );
  AND2_X1 AND2_144( .ZN(N972), .A1(N137), .A2(N528) );
  AND2_X1 AND2_145( .ZN(N975), .A1(N154), .A2(N273) );
  AND2_X1 AND2_146( .ZN(N978), .A1(N154), .A2(N290) );
  AND2_X1 AND2_147( .ZN(N981), .A1(N154), .A2(N307) );
  AND2_X1 AND2_148( .ZN(N984), .A1(N154), .A2(N324) );
  AND2_X1 AND2_149( .ZN(N987), .A1(N154), .A2(N341) );
  AND2_X1 AND2_150( .ZN(N990), .A1(N154), .A2(N358) );
  AND2_X1 AND2_151( .ZN(N993), .A1(N154), .A2(N375) );
  AND2_X1 AND2_152( .ZN(N996), .A1(N154), .A2(N392) );
  AND2_X1 AND2_153( .ZN(N999), .A1(N154), .A2(N409) );
  AND2_X1 AND2_154( .ZN(N1002), .A1(N154), .A2(N426) );
  AND2_X1 AND2_155( .ZN(N1005), .A1(N154), .A2(N443) );
  AND2_X1 AND2_156( .ZN(N1008), .A1(N154), .A2(N460) );
  AND2_X1 AND2_157( .ZN(N1011), .A1(N154), .A2(N477) );
  AND2_X1 AND2_158( .ZN(N1014), .A1(N154), .A2(N494) );
  AND2_X1 AND2_159( .ZN(N1017), .A1(N154), .A2(N511) );
  AND2_X4 AND2_160( .ZN(N1020), .A1(N154), .A2(N528) );
  AND2_X4 AND2_161( .ZN(N1023), .A1(N171), .A2(N273) );
  AND2_X4 AND2_162( .ZN(N1026), .A1(N171), .A2(N290) );
  AND2_X4 AND2_163( .ZN(N1029), .A1(N171), .A2(N307) );
  AND2_X4 AND2_164( .ZN(N1032), .A1(N171), .A2(N324) );
  AND2_X1 AND2_165( .ZN(N1035), .A1(N171), .A2(N341) );
  AND2_X1 AND2_166( .ZN(N1038), .A1(N171), .A2(N358) );
  AND2_X1 AND2_167( .ZN(N1041), .A1(N171), .A2(N375) );
  AND2_X1 AND2_168( .ZN(N1044), .A1(N171), .A2(N392) );
  AND2_X1 AND2_169( .ZN(N1047), .A1(N171), .A2(N409) );
  AND2_X1 AND2_170( .ZN(N1050), .A1(N171), .A2(N426) );
  AND2_X1 AND2_171( .ZN(N1053), .A1(N171), .A2(N443) );
  AND2_X1 AND2_172( .ZN(N1056), .A1(N171), .A2(N460) );
  AND2_X1 AND2_173( .ZN(N1059), .A1(N171), .A2(N477) );
  AND2_X1 AND2_174( .ZN(N1062), .A1(N171), .A2(N494) );
  AND2_X1 AND2_175( .ZN(N1065), .A1(N171), .A2(N511) );
  AND2_X1 AND2_176( .ZN(N1068), .A1(N171), .A2(N528) );
  AND2_X1 AND2_177( .ZN(N1071), .A1(N188), .A2(N273) );
  AND2_X1 AND2_178( .ZN(N1074), .A1(N188), .A2(N290) );
  AND2_X1 AND2_179( .ZN(N1077), .A1(N188), .A2(N307) );
  AND2_X1 AND2_180( .ZN(N1080), .A1(N188), .A2(N324) );
  AND2_X1 AND2_181( .ZN(N1083), .A1(N188), .A2(N341) );
  AND2_X1 AND2_182( .ZN(N1086), .A1(N188), .A2(N358) );
  AND2_X1 AND2_183( .ZN(N1089), .A1(N188), .A2(N375) );
  AND2_X1 AND2_184( .ZN(N1092), .A1(N188), .A2(N392) );
  AND2_X1 AND2_185( .ZN(N1095), .A1(N188), .A2(N409) );
  AND2_X1 AND2_186( .ZN(N1098), .A1(N188), .A2(N426) );
  AND2_X1 AND2_187( .ZN(N1101), .A1(N188), .A2(N443) );
  AND2_X1 AND2_188( .ZN(N1104), .A1(N188), .A2(N460) );
  AND2_X1 AND2_189( .ZN(N1107), .A1(N188), .A2(N477) );
  AND2_X1 AND2_190( .ZN(N1110), .A1(N188), .A2(N494) );
  AND2_X1 AND2_191( .ZN(N1113), .A1(N188), .A2(N511) );
  AND2_X1 AND2_192( .ZN(N1116), .A1(N188), .A2(N528) );
  AND2_X1 AND2_193( .ZN(N1119), .A1(N205), .A2(N273) );
  AND2_X1 AND2_194( .ZN(N1122), .A1(N205), .A2(N290) );
  AND2_X1 AND2_195( .ZN(N1125), .A1(N205), .A2(N307) );
  AND2_X1 AND2_196( .ZN(N1128), .A1(N205), .A2(N324) );
  AND2_X1 AND2_197( .ZN(N1131), .A1(N205), .A2(N341) );
  AND2_X1 AND2_198( .ZN(N1134), .A1(N205), .A2(N358) );
  AND2_X1 AND2_199( .ZN(N1137), .A1(N205), .A2(N375) );
  AND2_X1 AND2_200( .ZN(N1140), .A1(N205), .A2(N392) );
  AND2_X1 AND2_201( .ZN(N1143), .A1(N205), .A2(N409) );
  AND2_X1 AND2_202( .ZN(N1146), .A1(N205), .A2(N426) );
  AND2_X1 AND2_203( .ZN(N1149), .A1(N205), .A2(N443) );
  AND2_X1 AND2_204( .ZN(N1152), .A1(N205), .A2(N460) );
  AND2_X1 AND2_205( .ZN(N1155), .A1(N205), .A2(N477) );
  AND2_X1 AND2_206( .ZN(N1158), .A1(N205), .A2(N494) );
  AND2_X1 AND2_207( .ZN(N1161), .A1(N205), .A2(N511) );
  AND2_X1 AND2_208( .ZN(N1164), .A1(N205), .A2(N528) );
  AND2_X1 AND2_209( .ZN(N1167), .A1(N222), .A2(N273) );
  AND2_X1 AND2_210( .ZN(N1170), .A1(N222), .A2(N290) );
  AND2_X1 AND2_211( .ZN(N1173), .A1(N222), .A2(N307) );
  AND2_X1 AND2_212( .ZN(N1176), .A1(N222), .A2(N324) );
  AND2_X1 AND2_213( .ZN(N1179), .A1(N222), .A2(N341) );
  AND2_X1 AND2_214( .ZN(N1182), .A1(N222), .A2(N358) );
  AND2_X1 AND2_215( .ZN(N1185), .A1(N222), .A2(N375) );
  AND2_X1 AND2_216( .ZN(N1188), .A1(N222), .A2(N392) );
  AND2_X1 AND2_217( .ZN(N1191), .A1(N222), .A2(N409) );
  AND2_X1 AND2_218( .ZN(N1194), .A1(N222), .A2(N426) );
  AND2_X1 AND2_219( .ZN(N1197), .A1(N222), .A2(N443) );
  AND2_X1 AND2_220( .ZN(N1200), .A1(N222), .A2(N460) );
  AND2_X1 AND2_221( .ZN(N1203), .A1(N222), .A2(N477) );
  AND2_X1 AND2_222( .ZN(N1206), .A1(N222), .A2(N494) );
  AND2_X1 AND2_223( .ZN(N1209), .A1(N222), .A2(N511) );
  AND2_X1 AND2_224( .ZN(N1212), .A1(N222), .A2(N528) );
  AND2_X1 AND2_225( .ZN(N1215), .A1(N239), .A2(N273) );
  AND2_X1 AND2_226( .ZN(N1218), .A1(N239), .A2(N290) );
  AND2_X1 AND2_227( .ZN(N1221), .A1(N239), .A2(N307) );
  AND2_X1 AND2_228( .ZN(N1224), .A1(N239), .A2(N324) );
  AND2_X1 AND2_229( .ZN(N1227), .A1(N239), .A2(N341) );
  AND2_X1 AND2_230( .ZN(N1230), .A1(N239), .A2(N358) );
  AND2_X1 AND2_231( .ZN(N1233), .A1(N239), .A2(N375) );
  AND2_X1 AND2_232( .ZN(N1236), .A1(N239), .A2(N392) );
  AND2_X1 AND2_233( .ZN(N1239), .A1(N239), .A2(N409) );
  AND2_X1 AND2_234( .ZN(N1242), .A1(N239), .A2(N426) );
  AND2_X1 AND2_235( .ZN(N1245), .A1(N239), .A2(N443) );
  AND2_X1 AND2_236( .ZN(N1248), .A1(N239), .A2(N460) );
  AND2_X1 AND2_237( .ZN(N1251), .A1(N239), .A2(N477) );
  AND2_X1 AND2_238( .ZN(N1254), .A1(N239), .A2(N494) );
  AND2_X1 AND2_239( .ZN(N1257), .A1(N239), .A2(N511) );
  AND2_X1 AND2_240( .ZN(N1260), .A1(N239), .A2(N528) );
  AND2_X1 AND2_241( .ZN(N1263), .A1(N256), .A2(N273) );
  AND2_X1 AND2_242( .ZN(N1266), .A1(N256), .A2(N290) );
  AND2_X1 AND2_243( .ZN(N1269), .A1(N256), .A2(N307) );
  AND2_X1 AND2_244( .ZN(N1272), .A1(N256), .A2(N324) );
  AND2_X1 AND2_245( .ZN(N1275), .A1(N256), .A2(N341) );
  AND2_X1 AND2_246( .ZN(N1278), .A1(N256), .A2(N358) );
  AND2_X1 AND2_247( .ZN(N1281), .A1(N256), .A2(N375) );
  AND2_X1 AND2_248( .ZN(N1284), .A1(N256), .A2(N392) );
  AND2_X1 AND2_249( .ZN(N1287), .A1(N256), .A2(N409) );
  AND2_X1 AND2_250( .ZN(N1290), .A1(N256), .A2(N426) );
  AND2_X1 AND2_251( .ZN(N1293), .A1(N256), .A2(N443) );
  AND2_X1 AND2_252( .ZN(N1296), .A1(N256), .A2(N460) );
  AND2_X1 AND2_253( .ZN(N1299), .A1(N256), .A2(N477) );
  AND2_X1 AND2_254( .ZN(N1302), .A1(N256), .A2(N494) );
  AND2_X1 AND2_255( .ZN(N1305), .A1(N256), .A2(N511) );
  AND2_X1 AND2_256( .ZN(N1308), .A1(N256), .A2(N528) );
  INV_X1 NOT1_257( .ZN(N1311), .A(N591) );
  INV_X8 NOT1_258( .ZN(N1315), .A(N639) );
  INV_X8 NOT1_259( .ZN(N1319), .A(N687) );
  INV_X8 NOT1_260( .ZN(N1323), .A(N735) );
  INV_X8 NOT1_261( .ZN(N1327), .A(N783) );
  INV_X8 NOT1_262( .ZN(N1331), .A(N831) );
  INV_X8 NOT1_263( .ZN(N1335), .A(N879) );
  INV_X1 NOT1_264( .ZN(N1339), .A(N927) );
  INV_X1 NOT1_265( .ZN(N1343), .A(N975) );
  INV_X1 NOT1_266( .ZN(N1347), .A(N1023) );
  INV_X1 NOT1_267( .ZN(N1351), .A(N1071) );
  INV_X1 NOT1_268( .ZN(N1355), .A(N1119) );
  INV_X1 NOT1_269( .ZN(N1359), .A(N1167) );
  INV_X1 NOT1_270( .ZN(N1363), .A(N1215) );
  INV_X1 NOT1_271( .ZN(N1367), .A(N1263) );
  NOR2_X1 NOR2_272( .ZN(N1371), .A1(N591), .A2(N1311) );
  INV_X1 NOT1_273( .ZN(N1372), .A(N1311) );
  NOR2_X1 NOR2_274( .ZN(N1373), .A1(N639), .A2(N1315) );
  INV_X1 NOT1_275( .ZN(N1374), .A(N1315) );
  NOR2_X1 NOR2_276( .ZN(N1375), .A1(N687), .A2(N1319) );
  INV_X1 NOT1_277( .ZN(N1376), .A(N1319) );
  NOR2_X1 NOR2_278( .ZN(N1377), .A1(N735), .A2(N1323) );
  INV_X1 NOT1_279( .ZN(N1378), .A(N1323) );
  NOR2_X1 NOR2_280( .ZN(N1379), .A1(N783), .A2(N1327) );
  INV_X1 NOT1_281( .ZN(N1380), .A(N1327) );
  NOR2_X1 NOR2_282( .ZN(N1381), .A1(N831), .A2(N1331) );
  INV_X1 NOT1_283( .ZN(N1382), .A(N1331) );
  NOR2_X1 NOR2_284( .ZN(N1383), .A1(N879), .A2(N1335) );
  INV_X1 NOT1_285( .ZN(N1384), .A(N1335) );
  NOR2_X1 NOR2_286( .ZN(N1385), .A1(N927), .A2(N1339) );
  INV_X1 NOT1_287( .ZN(N1386), .A(N1339) );
  NOR2_X1 NOR2_288( .ZN(N1387), .A1(N975), .A2(N1343) );
  INV_X8 NOT1_289( .ZN(N1388), .A(N1343) );
  NOR2_X1 NOR2_290( .ZN(N1389), .A1(N1023), .A2(N1347) );
  INV_X1 NOT1_291( .ZN(N1390), .A(N1347) );
  NOR2_X1 NOR2_292( .ZN(N1391), .A1(N1071), .A2(N1351) );
  INV_X1 NOT1_293( .ZN(N1392), .A(N1351) );
  NOR2_X1 NOR2_294( .ZN(N1393), .A1(N1119), .A2(N1355) );
  INV_X1 NOT1_295( .ZN(N1394), .A(N1355) );
  NOR2_X1 NOR2_296( .ZN(N1395), .A1(N1167), .A2(N1359) );
  INV_X1 NOT1_297( .ZN(N1396), .A(N1359) );
  NOR2_X1 NOR2_298( .ZN(N1397), .A1(N1215), .A2(N1363) );
  INV_X1 NOT1_299( .ZN(N1398), .A(N1363) );
  NOR2_X1 NOR2_300( .ZN(N1399), .A1(N1263), .A2(N1367) );
  INV_X1 NOT1_301( .ZN(N1400), .A(N1367) );
  NOR2_X1 NOR2_302( .ZN(N1401), .A1(N1371), .A2(N1372) );
  NOR2_X1 NOR2_303( .ZN(N1404), .A1(N1373), .A2(N1374) );
  NOR2_X2 NOR2_304( .ZN(N1407), .A1(N1375), .A2(N1376) );
  NOR2_X2 NOR2_305( .ZN(N1410), .A1(N1377), .A2(N1378) );
  NOR2_X2 NOR2_306( .ZN(N1413), .A1(N1379), .A2(N1380) );
  NOR2_X2 NOR2_307( .ZN(N1416), .A1(N1381), .A2(N1382) );
  NOR2_X2 NOR2_308( .ZN(N1419), .A1(N1383), .A2(N1384) );
  NOR2_X2 NOR2_309( .ZN(N1422), .A1(N1385), .A2(N1386) );
  NOR2_X1 NOR2_310( .ZN(N1425), .A1(N1387), .A2(N1388) );
  NOR2_X1 NOR2_311( .ZN(N1428), .A1(N1389), .A2(N1390) );
  NOR2_X1 NOR2_312( .ZN(N1431), .A1(N1391), .A2(N1392) );
  NOR2_X1 NOR2_313( .ZN(N1434), .A1(N1393), .A2(N1394) );
  NOR2_X1 NOR2_314( .ZN(N1437), .A1(N1395), .A2(N1396) );
  NOR2_X1 NOR2_315( .ZN(N1440), .A1(N1397), .A2(N1398) );
  NOR2_X1 NOR2_316( .ZN(N1443), .A1(N1399), .A2(N1400) );
  NOR2_X1 NOR2_317( .ZN(N1446), .A1(N1401), .A2(N546) );
  NOR2_X1 NOR2_318( .ZN(N1450), .A1(N1404), .A2(N594) );
  NOR2_X1 NOR2_319( .ZN(N1454), .A1(N1407), .A2(N642) );
  NOR2_X1 NOR2_320( .ZN(N1458), .A1(N1410), .A2(N690) );
  NOR2_X1 NOR2_321( .ZN(N1462), .A1(N1413), .A2(N738) );
  NOR2_X1 NOR2_322( .ZN(N1466), .A1(N1416), .A2(N786) );
  NOR2_X1 NOR2_323( .ZN(N1470), .A1(N1419), .A2(N834) );
  NOR2_X1 NOR2_324( .ZN(N1474), .A1(N1422), .A2(N882) );
  NOR2_X1 NOR2_325( .ZN(N1478), .A1(N1425), .A2(N930) );
  NOR2_X1 NOR2_326( .ZN(N1482), .A1(N1428), .A2(N978) );
  NOR2_X1 NOR2_327( .ZN(N1486), .A1(N1431), .A2(N1026) );
  NOR2_X1 NOR2_328( .ZN(N1490), .A1(N1434), .A2(N1074) );
  NOR2_X1 NOR2_329( .ZN(N1494), .A1(N1437), .A2(N1122) );
  NOR2_X1 NOR2_330( .ZN(N1498), .A1(N1440), .A2(N1170) );
  NOR2_X1 NOR2_331( .ZN(N1502), .A1(N1443), .A2(N1218) );
  NOR2_X1 NOR2_332( .ZN(N1506), .A1(N1401), .A2(N1446) );
  NOR2_X1 NOR2_333( .ZN(N1507), .A1(N1446), .A2(N546) );
  NOR2_X1 NOR2_334( .ZN(N1508), .A1(N1311), .A2(N1446) );
  NOR2_X1 NOR2_335( .ZN(N1511), .A1(N1404), .A2(N1450) );
  NOR2_X1 NOR2_336( .ZN(N1512), .A1(N1450), .A2(N594) );
  NOR2_X1 NOR2_337( .ZN(N1513), .A1(N1315), .A2(N1450) );
  NOR2_X1 NOR2_338( .ZN(N1516), .A1(N1407), .A2(N1454) );
  NOR2_X1 NOR2_339( .ZN(N1517), .A1(N1454), .A2(N642) );
  NOR2_X1 NOR2_340( .ZN(N1518), .A1(N1319), .A2(N1454) );
  NOR2_X1 NOR2_341( .ZN(N1521), .A1(N1410), .A2(N1458) );
  NOR2_X1 NOR2_342( .ZN(N1522), .A1(N1458), .A2(N690) );
  NOR2_X1 NOR2_343( .ZN(N1523), .A1(N1323), .A2(N1458) );
  NOR2_X1 NOR2_344( .ZN(N1526), .A1(N1413), .A2(N1462) );
  NOR2_X1 NOR2_345( .ZN(N1527), .A1(N1462), .A2(N738) );
  NOR2_X1 NOR2_346( .ZN(N1528), .A1(N1327), .A2(N1462) );
  NOR2_X1 NOR2_347( .ZN(N1531), .A1(N1416), .A2(N1466) );
  NOR2_X1 NOR2_348( .ZN(N1532), .A1(N1466), .A2(N786) );
  NOR2_X1 NOR2_349( .ZN(N1533), .A1(N1331), .A2(N1466) );
  NOR2_X1 NOR2_350( .ZN(N1536), .A1(N1419), .A2(N1470) );
  NOR2_X1 NOR2_351( .ZN(N1537), .A1(N1470), .A2(N834) );
  NOR2_X1 NOR2_352( .ZN(N1538), .A1(N1335), .A2(N1470) );
  NOR2_X1 NOR2_353( .ZN(N1541), .A1(N1422), .A2(N1474) );
  NOR2_X1 NOR2_354( .ZN(N1542), .A1(N1474), .A2(N882) );
  NOR2_X1 NOR2_355( .ZN(N1543), .A1(N1339), .A2(N1474) );
  NOR2_X1 NOR2_356( .ZN(N1546), .A1(N1425), .A2(N1478) );
  NOR2_X1 NOR2_357( .ZN(N1547), .A1(N1478), .A2(N930) );
  NOR2_X1 NOR2_358( .ZN(N1548), .A1(N1343), .A2(N1478) );
  NOR2_X1 NOR2_359( .ZN(N1551), .A1(N1428), .A2(N1482) );
  NOR2_X1 NOR2_360( .ZN(N1552), .A1(N1482), .A2(N978) );
  NOR2_X1 NOR2_361( .ZN(N1553), .A1(N1347), .A2(N1482) );
  NOR2_X1 NOR2_362( .ZN(N1556), .A1(N1431), .A2(N1486) );
  NOR2_X1 NOR2_363( .ZN(N1557), .A1(N1486), .A2(N1026) );
  NOR2_X1 NOR2_364( .ZN(N1558), .A1(N1351), .A2(N1486) );
  NOR2_X1 NOR2_365( .ZN(N1561), .A1(N1434), .A2(N1490) );
  NOR2_X1 NOR2_366( .ZN(N1562), .A1(N1490), .A2(N1074) );
  NOR2_X1 NOR2_367( .ZN(N1563), .A1(N1355), .A2(N1490) );
  NOR2_X1 NOR2_368( .ZN(N1566), .A1(N1437), .A2(N1494) );
  NOR2_X1 NOR2_369( .ZN(N1567), .A1(N1494), .A2(N1122) );
  NOR2_X1 NOR2_370( .ZN(N1568), .A1(N1359), .A2(N1494) );
  NOR2_X1 NOR2_371( .ZN(N1571), .A1(N1440), .A2(N1498) );
  NOR2_X1 NOR2_372( .ZN(N1572), .A1(N1498), .A2(N1170) );
  NOR2_X1 NOR2_373( .ZN(N1573), .A1(N1363), .A2(N1498) );
  NOR2_X1 NOR2_374( .ZN(N1576), .A1(N1443), .A2(N1502) );
  NOR2_X1 NOR2_375( .ZN(N1577), .A1(N1502), .A2(N1218) );
  NOR2_X1 NOR2_376( .ZN(N1578), .A1(N1367), .A2(N1502) );
  NOR2_X1 NOR2_377( .ZN(N1581), .A1(N1506), .A2(N1507) );
  NOR2_X1 NOR2_378( .ZN(N1582), .A1(N1511), .A2(N1512) );
  NOR2_X1 NOR2_379( .ZN(N1585), .A1(N1516), .A2(N1517) );
  NOR2_X1 NOR2_380( .ZN(N1588), .A1(N1521), .A2(N1522) );
  NOR2_X1 NOR2_381( .ZN(N1591), .A1(N1526), .A2(N1527) );
  NOR2_X1 NOR2_382( .ZN(N1594), .A1(N1531), .A2(N1532) );
  NOR2_X1 NOR2_383( .ZN(N1597), .A1(N1536), .A2(N1537) );
  NOR2_X1 NOR2_384( .ZN(N1600), .A1(N1541), .A2(N1542) );
  NOR2_X1 NOR2_385( .ZN(N1603), .A1(N1546), .A2(N1547) );
  NOR2_X1 NOR2_386( .ZN(N1606), .A1(N1551), .A2(N1552) );
  NOR2_X1 NOR2_387( .ZN(N1609), .A1(N1556), .A2(N1557) );
  NOR2_X1 NOR2_388( .ZN(N1612), .A1(N1561), .A2(N1562) );
  NOR2_X1 NOR2_389( .ZN(N1615), .A1(N1566), .A2(N1567) );
  NOR2_X1 NOR2_390( .ZN(N1618), .A1(N1571), .A2(N1572) );
  NOR2_X1 NOR2_391( .ZN(N1621), .A1(N1576), .A2(N1577) );
  NOR2_X1 NOR2_392( .ZN(N1624), .A1(N1266), .A2(N1578) );
  NOR2_X1 NOR2_393( .ZN(N1628), .A1(N1582), .A2(N1508) );
  NOR2_X1 NOR2_394( .ZN(N1632), .A1(N1585), .A2(N1513) );
  NOR2_X1 NOR2_395( .ZN(N1636), .A1(N1588), .A2(N1518) );
  NOR2_X1 NOR2_396( .ZN(N1640), .A1(N1591), .A2(N1523) );
  NOR2_X1 NOR2_397( .ZN(N1644), .A1(N1594), .A2(N1528) );
  NOR2_X2 NOR2_398( .ZN(N1648), .A1(N1597), .A2(N1533) );
  NOR2_X2 NOR2_399( .ZN(N1652), .A1(N1600), .A2(N1538) );
  NOR2_X2 NOR2_400( .ZN(N1656), .A1(N1603), .A2(N1543) );
  NOR2_X2 NOR2_401( .ZN(N1660), .A1(N1606), .A2(N1548) );
  NOR2_X2 NOR2_402( .ZN(N1664), .A1(N1609), .A2(N1553) );
  NOR2_X2 NOR2_403( .ZN(N1668), .A1(N1612), .A2(N1558) );
  NOR2_X1 NOR2_404( .ZN(N1672), .A1(N1615), .A2(N1563) );
  NOR2_X1 NOR2_405( .ZN(N1676), .A1(N1618), .A2(N1568) );
  NOR2_X1 NOR2_406( .ZN(N1680), .A1(N1621), .A2(N1573) );
  NOR2_X1 NOR2_407( .ZN(N1684), .A1(N1266), .A2(N1624) );
  NOR2_X1 NOR2_408( .ZN(N1685), .A1(N1624), .A2(N1578) );
  NOR2_X1 NOR2_409( .ZN(N1686), .A1(N1582), .A2(N1628) );
  NOR2_X1 NOR2_410( .ZN(N1687), .A1(N1628), .A2(N1508) );
  NOR2_X1 NOR2_411( .ZN(N1688), .A1(N1585), .A2(N1632) );
  NOR2_X1 NOR2_412( .ZN(N1689), .A1(N1632), .A2(N1513) );
  NOR2_X1 NOR2_413( .ZN(N1690), .A1(N1588), .A2(N1636) );
  NOR2_X1 NOR2_414( .ZN(N1691), .A1(N1636), .A2(N1518) );
  NOR2_X1 NOR2_415( .ZN(N1692), .A1(N1591), .A2(N1640) );
  NOR2_X1 NOR2_416( .ZN(N1693), .A1(N1640), .A2(N1523) );
  NOR2_X1 NOR2_417( .ZN(N1694), .A1(N1594), .A2(N1644) );
  NOR2_X1 NOR2_418( .ZN(N1695), .A1(N1644), .A2(N1528) );
  NOR2_X1 NOR2_419( .ZN(N1696), .A1(N1597), .A2(N1648) );
  NOR2_X1 NOR2_420( .ZN(N1697), .A1(N1648), .A2(N1533) );
  NOR2_X1 NOR2_421( .ZN(N1698), .A1(N1600), .A2(N1652) );
  NOR2_X1 NOR2_422( .ZN(N1699), .A1(N1652), .A2(N1538) );
  NOR2_X1 NOR2_423( .ZN(N1700), .A1(N1603), .A2(N1656) );
  NOR2_X1 NOR2_424( .ZN(N1701), .A1(N1656), .A2(N1543) );
  NOR2_X1 NOR2_425( .ZN(N1702), .A1(N1606), .A2(N1660) );
  NOR2_X1 NOR2_426( .ZN(N1703), .A1(N1660), .A2(N1548) );
  NOR2_X1 NOR2_427( .ZN(N1704), .A1(N1609), .A2(N1664) );
  NOR2_X1 NOR2_428( .ZN(N1705), .A1(N1664), .A2(N1553) );
  NOR2_X1 NOR2_429( .ZN(N1706), .A1(N1612), .A2(N1668) );
  NOR2_X1 NOR2_430( .ZN(N1707), .A1(N1668), .A2(N1558) );
  NOR2_X1 NOR2_431( .ZN(N1708), .A1(N1615), .A2(N1672) );
  NOR2_X1 NOR2_432( .ZN(N1709), .A1(N1672), .A2(N1563) );
  NOR2_X1 NOR2_433( .ZN(N1710), .A1(N1618), .A2(N1676) );
  NOR2_X1 NOR2_434( .ZN(N1711), .A1(N1676), .A2(N1568) );
  NOR2_X1 NOR2_435( .ZN(N1712), .A1(N1621), .A2(N1680) );
  NOR2_X1 NOR2_436( .ZN(N1713), .A1(N1680), .A2(N1573) );
  NOR2_X1 NOR2_437( .ZN(N1714), .A1(N1684), .A2(N1685) );
  NOR2_X1 NOR2_438( .ZN(N1717), .A1(N1686), .A2(N1687) );
  NOR2_X1 NOR2_439( .ZN(N1720), .A1(N1688), .A2(N1689) );
  NOR2_X1 NOR2_440( .ZN(N1723), .A1(N1690), .A2(N1691) );
  NOR2_X1 NOR2_441( .ZN(N1726), .A1(N1692), .A2(N1693) );
  NOR2_X1 NOR2_442( .ZN(N1729), .A1(N1694), .A2(N1695) );
  NOR2_X1 NOR2_443( .ZN(N1732), .A1(N1696), .A2(N1697) );
  NOR2_X1 NOR2_444( .ZN(N1735), .A1(N1698), .A2(N1699) );
  NOR2_X1 NOR2_445( .ZN(N1738), .A1(N1700), .A2(N1701) );
  NOR2_X1 NOR2_446( .ZN(N1741), .A1(N1702), .A2(N1703) );
  NOR2_X1 NOR2_447( .ZN(N1744), .A1(N1704), .A2(N1705) );
  NOR2_X1 NOR2_448( .ZN(N1747), .A1(N1706), .A2(N1707) );
  NOR2_X1 NOR2_449( .ZN(N1750), .A1(N1708), .A2(N1709) );
  NOR2_X1 NOR2_450( .ZN(N1753), .A1(N1710), .A2(N1711) );
  NOR2_X1 NOR2_451( .ZN(N1756), .A1(N1712), .A2(N1713) );
  NOR2_X1 NOR2_452( .ZN(N1759), .A1(N1714), .A2(N1221) );
  NOR2_X1 NOR2_453( .ZN(N1763), .A1(N1717), .A2(N549) );
  NOR2_X1 NOR2_454( .ZN(N1767), .A1(N1720), .A2(N597) );
  NOR2_X1 NOR2_455( .ZN(N1771), .A1(N1723), .A2(N645) );
  NOR2_X1 NOR2_456( .ZN(N1775), .A1(N1726), .A2(N693) );
  NOR2_X1 NOR2_457( .ZN(N1779), .A1(N1729), .A2(N741) );
  NOR2_X1 NOR2_458( .ZN(N1783), .A1(N1732), .A2(N789) );
  NOR2_X1 NOR2_459( .ZN(N1787), .A1(N1735), .A2(N837) );
  NOR2_X1 NOR2_460( .ZN(N1791), .A1(N1738), .A2(N885) );
  NOR2_X1 NOR2_461( .ZN(N1795), .A1(N1741), .A2(N933) );
  NOR2_X1 NOR2_462( .ZN(N1799), .A1(N1744), .A2(N981) );
  NOR2_X1 NOR2_463( .ZN(N1803), .A1(N1747), .A2(N1029) );
  NOR2_X1 NOR2_464( .ZN(N1807), .A1(N1750), .A2(N1077) );
  NOR2_X1 NOR2_465( .ZN(N1811), .A1(N1753), .A2(N1125) );
  NOR2_X1 NOR2_466( .ZN(N1815), .A1(N1756), .A2(N1173) );
  NOR2_X1 NOR2_467( .ZN(N1819), .A1(N1714), .A2(N1759) );
  NOR2_X1 NOR2_468( .ZN(N1820), .A1(N1759), .A2(N1221) );
  NOR2_X1 NOR2_469( .ZN(N1821), .A1(N1624), .A2(N1759) );
  NOR2_X1 NOR2_470( .ZN(N1824), .A1(N1717), .A2(N1763) );
  NOR2_X1 NOR2_471( .ZN(N1825), .A1(N1763), .A2(N549) );
  NOR2_X1 NOR2_472( .ZN(N1826), .A1(N1628), .A2(N1763) );
  NOR2_X1 NOR2_473( .ZN(N1829), .A1(N1720), .A2(N1767) );
  NOR2_X1 NOR2_474( .ZN(N1830), .A1(N1767), .A2(N597) );
  NOR2_X1 NOR2_475( .ZN(N1831), .A1(N1632), .A2(N1767) );
  NOR2_X1 NOR2_476( .ZN(N1834), .A1(N1723), .A2(N1771) );
  NOR2_X1 NOR2_477( .ZN(N1835), .A1(N1771), .A2(N645) );
  NOR2_X1 NOR2_478( .ZN(N1836), .A1(N1636), .A2(N1771) );
  NOR2_X1 NOR2_479( .ZN(N1839), .A1(N1726), .A2(N1775) );
  NOR2_X1 NOR2_480( .ZN(N1840), .A1(N1775), .A2(N693) );
  NOR2_X1 NOR2_481( .ZN(N1841), .A1(N1640), .A2(N1775) );
  NOR2_X1 NOR2_482( .ZN(N1844), .A1(N1729), .A2(N1779) );
  NOR2_X1 NOR2_483( .ZN(N1845), .A1(N1779), .A2(N741) );
  NOR2_X1 NOR2_484( .ZN(N1846), .A1(N1644), .A2(N1779) );
  NOR2_X1 NOR2_485( .ZN(N1849), .A1(N1732), .A2(N1783) );
  NOR2_X1 NOR2_486( .ZN(N1850), .A1(N1783), .A2(N789) );
  NOR2_X1 NOR2_487( .ZN(N1851), .A1(N1648), .A2(N1783) );
  NOR2_X1 NOR2_488( .ZN(N1854), .A1(N1735), .A2(N1787) );
  NOR2_X1 NOR2_489( .ZN(N1855), .A1(N1787), .A2(N837) );
  NOR2_X1 NOR2_490( .ZN(N1856), .A1(N1652), .A2(N1787) );
  NOR2_X1 NOR2_491( .ZN(N1859), .A1(N1738), .A2(N1791) );
  NOR2_X1 NOR2_492( .ZN(N1860), .A1(N1791), .A2(N885) );
  NOR2_X1 NOR2_493( .ZN(N1861), .A1(N1656), .A2(N1791) );
  NOR2_X1 NOR2_494( .ZN(N1864), .A1(N1741), .A2(N1795) );
  NOR2_X1 NOR2_495( .ZN(N1865), .A1(N1795), .A2(N933) );
  NOR2_X1 NOR2_496( .ZN(N1866), .A1(N1660), .A2(N1795) );
  NOR2_X1 NOR2_497( .ZN(N1869), .A1(N1744), .A2(N1799) );
  NOR2_X1 NOR2_498( .ZN(N1870), .A1(N1799), .A2(N981) );
  NOR2_X1 NOR2_499( .ZN(N1871), .A1(N1664), .A2(N1799) );
  NOR2_X1 NOR2_500( .ZN(N1874), .A1(N1747), .A2(N1803) );
  NOR2_X1 NOR2_501( .ZN(N1875), .A1(N1803), .A2(N1029) );
  NOR2_X1 NOR2_502( .ZN(N1876), .A1(N1668), .A2(N1803) );
  NOR2_X1 NOR2_503( .ZN(N1879), .A1(N1750), .A2(N1807) );
  NOR2_X1 NOR2_504( .ZN(N1880), .A1(N1807), .A2(N1077) );
  NOR2_X1 NOR2_505( .ZN(N1881), .A1(N1672), .A2(N1807) );
  NOR2_X1 NOR2_506( .ZN(N1884), .A1(N1753), .A2(N1811) );
  NOR2_X1 NOR2_507( .ZN(N1885), .A1(N1811), .A2(N1125) );
  NOR2_X1 NOR2_508( .ZN(N1886), .A1(N1676), .A2(N1811) );
  NOR2_X1 NOR2_509( .ZN(N1889), .A1(N1756), .A2(N1815) );
  NOR2_X1 NOR2_510( .ZN(N1890), .A1(N1815), .A2(N1173) );
  NOR2_X1 NOR2_511( .ZN(N1891), .A1(N1680), .A2(N1815) );
  NOR2_X1 NOR2_512( .ZN(N1894), .A1(N1819), .A2(N1820) );
  NOR2_X1 NOR2_513( .ZN(N1897), .A1(N1269), .A2(N1821) );
  NOR2_X1 NOR2_514( .ZN(N1901), .A1(N1824), .A2(N1825) );
  NOR2_X1 NOR2_515( .ZN(N1902), .A1(N1829), .A2(N1830) );
  NOR2_X1 NOR2_516( .ZN(N1905), .A1(N1834), .A2(N1835) );
  NOR2_X1 NOR2_517( .ZN(N1908), .A1(N1839), .A2(N1840) );
  NOR2_X1 NOR2_518( .ZN(N1911), .A1(N1844), .A2(N1845) );
  NOR2_X1 NOR2_519( .ZN(N1914), .A1(N1849), .A2(N1850) );
  NOR2_X1 NOR2_520( .ZN(N1917), .A1(N1854), .A2(N1855) );
  NOR2_X1 NOR2_521( .ZN(N1920), .A1(N1859), .A2(N1860) );
  NOR2_X1 NOR2_522( .ZN(N1923), .A1(N1864), .A2(N1865) );
  NOR2_X1 NOR2_523( .ZN(N1926), .A1(N1869), .A2(N1870) );
  NOR2_X1 NOR2_524( .ZN(N1929), .A1(N1874), .A2(N1875) );
  NOR2_X1 NOR2_525( .ZN(N1932), .A1(N1879), .A2(N1880) );
  NOR2_X1 NOR2_526( .ZN(N1935), .A1(N1884), .A2(N1885) );
  NOR2_X1 NOR2_527( .ZN(N1938), .A1(N1889), .A2(N1890) );
  NOR2_X1 NOR2_528( .ZN(N1941), .A1(N1894), .A2(N1891) );
  NOR2_X1 NOR2_529( .ZN(N1945), .A1(N1269), .A2(N1897) );
  NOR2_X1 NOR2_530( .ZN(N1946), .A1(N1897), .A2(N1821) );
  NOR2_X2 NOR2_531( .ZN(N1947), .A1(N1902), .A2(N1826) );
  NOR2_X2 NOR2_532( .ZN(N1951), .A1(N1905), .A2(N1831) );
  NOR2_X2 NOR2_533( .ZN(N1955), .A1(N1908), .A2(N1836) );
  NOR2_X2 NOR2_534( .ZN(N1959), .A1(N1911), .A2(N1841) );
  NOR2_X1 NOR2_535( .ZN(N1963), .A1(N1914), .A2(N1846) );
  NOR2_X1 NOR2_536( .ZN(N1967), .A1(N1917), .A2(N1851) );
  NOR2_X1 NOR2_537( .ZN(N1971), .A1(N1920), .A2(N1856) );
  NOR2_X1 NOR2_538( .ZN(N1975), .A1(N1923), .A2(N1861) );
  NOR2_X1 NOR2_539( .ZN(N1979), .A1(N1926), .A2(N1866) );
  NOR2_X1 NOR2_540( .ZN(N1983), .A1(N1929), .A2(N1871) );
  NOR2_X1 NOR2_541( .ZN(N1987), .A1(N1932), .A2(N1876) );
  NOR2_X1 NOR2_542( .ZN(N1991), .A1(N1935), .A2(N1881) );
  NOR2_X1 NOR2_543( .ZN(N1995), .A1(N1938), .A2(N1886) );
  NOR2_X1 NOR2_544( .ZN(N1999), .A1(N1894), .A2(N1941) );
  NOR2_X1 NOR2_545( .ZN(N2000), .A1(N1941), .A2(N1891) );
  NOR2_X1 NOR2_546( .ZN(N2001), .A1(N1945), .A2(N1946) );
  NOR2_X1 NOR2_547( .ZN(N2004), .A1(N1902), .A2(N1947) );
  NOR2_X1 NOR2_548( .ZN(N2005), .A1(N1947), .A2(N1826) );
  NOR2_X1 NOR2_549( .ZN(N2006), .A1(N1905), .A2(N1951) );
  NOR2_X1 NOR2_550( .ZN(N2007), .A1(N1951), .A2(N1831) );
  NOR2_X1 NOR2_551( .ZN(N2008), .A1(N1908), .A2(N1955) );
  NOR2_X1 NOR2_552( .ZN(N2009), .A1(N1955), .A2(N1836) );
  NOR2_X1 NOR2_553( .ZN(N2010), .A1(N1911), .A2(N1959) );
  NOR2_X1 NOR2_554( .ZN(N2011), .A1(N1959), .A2(N1841) );
  NOR2_X1 NOR2_555( .ZN(N2012), .A1(N1914), .A2(N1963) );
  NOR2_X1 NOR2_556( .ZN(N2013), .A1(N1963), .A2(N1846) );
  NOR2_X1 NOR2_557( .ZN(N2014), .A1(N1917), .A2(N1967) );
  NOR2_X1 NOR2_558( .ZN(N2015), .A1(N1967), .A2(N1851) );
  NOR2_X1 NOR2_559( .ZN(N2016), .A1(N1920), .A2(N1971) );
  NOR2_X1 NOR2_560( .ZN(N2017), .A1(N1971), .A2(N1856) );
  NOR2_X1 NOR2_561( .ZN(N2018), .A1(N1923), .A2(N1975) );
  NOR2_X1 NOR2_562( .ZN(N2019), .A1(N1975), .A2(N1861) );
  NOR2_X1 NOR2_563( .ZN(N2020), .A1(N1926), .A2(N1979) );
  NOR2_X1 NOR2_564( .ZN(N2021), .A1(N1979), .A2(N1866) );
  NOR2_X1 NOR2_565( .ZN(N2022), .A1(N1929), .A2(N1983) );
  NOR2_X1 NOR2_566( .ZN(N2023), .A1(N1983), .A2(N1871) );
  NOR2_X1 NOR2_567( .ZN(N2024), .A1(N1932), .A2(N1987) );
  NOR2_X1 NOR2_568( .ZN(N2025), .A1(N1987), .A2(N1876) );
  NOR2_X1 NOR2_569( .ZN(N2026), .A1(N1935), .A2(N1991) );
  NOR2_X1 NOR2_570( .ZN(N2027), .A1(N1991), .A2(N1881) );
  NOR2_X1 NOR2_571( .ZN(N2028), .A1(N1938), .A2(N1995) );
  NOR2_X1 NOR2_572( .ZN(N2029), .A1(N1995), .A2(N1886) );
  NOR2_X1 NOR2_573( .ZN(N2030), .A1(N1999), .A2(N2000) );
  NOR2_X1 NOR2_574( .ZN(N2033), .A1(N2001), .A2(N1224) );
  NOR2_X1 NOR2_575( .ZN(N2037), .A1(N2004), .A2(N2005) );
  NOR2_X1 NOR2_576( .ZN(N2040), .A1(N2006), .A2(N2007) );
  NOR2_X1 NOR2_577( .ZN(N2043), .A1(N2008), .A2(N2009) );
  NOR2_X1 NOR2_578( .ZN(N2046), .A1(N2010), .A2(N2011) );
  NOR2_X1 NOR2_579( .ZN(N2049), .A1(N2012), .A2(N2013) );
  NOR2_X1 NOR2_580( .ZN(N2052), .A1(N2014), .A2(N2015) );
  NOR2_X1 NOR2_581( .ZN(N2055), .A1(N2016), .A2(N2017) );
  NOR2_X1 NOR2_582( .ZN(N2058), .A1(N2018), .A2(N2019) );
  NOR2_X1 NOR2_583( .ZN(N2061), .A1(N2020), .A2(N2021) );
  NOR2_X1 NOR2_584( .ZN(N2064), .A1(N2022), .A2(N2023) );
  NOR2_X1 NOR2_585( .ZN(N2067), .A1(N2024), .A2(N2025) );
  NOR2_X1 NOR2_586( .ZN(N2070), .A1(N2026), .A2(N2027) );
  NOR2_X1 NOR2_587( .ZN(N2073), .A1(N2028), .A2(N2029) );
  NOR2_X1 NOR2_588( .ZN(N2076), .A1(N2030), .A2(N1176) );
  NOR2_X1 NOR2_589( .ZN(N2080), .A1(N2001), .A2(N2033) );
  NOR2_X1 NOR2_590( .ZN(N2081), .A1(N2033), .A2(N1224) );
  NOR2_X1 NOR2_591( .ZN(N2082), .A1(N1897), .A2(N2033) );
  NOR2_X1 NOR2_592( .ZN(N2085), .A1(N2037), .A2(N552) );
  NOR2_X1 NOR2_593( .ZN(N2089), .A1(N2040), .A2(N600) );
  NOR2_X1 NOR2_594( .ZN(N2093), .A1(N2043), .A2(N648) );
  NOR2_X1 NOR2_595( .ZN(N2097), .A1(N2046), .A2(N696) );
  NOR2_X1 NOR2_596( .ZN(N2101), .A1(N2049), .A2(N744) );
  NOR2_X1 NOR2_597( .ZN(N2105), .A1(N2052), .A2(N792) );
  NOR2_X1 NOR2_598( .ZN(N2109), .A1(N2055), .A2(N840) );
  NOR2_X1 NOR2_599( .ZN(N2113), .A1(N2058), .A2(N888) );
  NOR2_X1 NOR2_600( .ZN(N2117), .A1(N2061), .A2(N936) );
  NOR2_X1 NOR2_601( .ZN(N2121), .A1(N2064), .A2(N984) );
  NOR2_X1 NOR2_602( .ZN(N2125), .A1(N2067), .A2(N1032) );
  NOR2_X1 NOR2_603( .ZN(N2129), .A1(N2070), .A2(N1080) );
  NOR2_X1 NOR2_604( .ZN(N2133), .A1(N2073), .A2(N1128) );
  NOR2_X1 NOR2_605( .ZN(N2137), .A1(N2030), .A2(N2076) );
  NOR2_X1 NOR2_606( .ZN(N2138), .A1(N2076), .A2(N1176) );
  NOR2_X1 NOR2_607( .ZN(N2139), .A1(N1941), .A2(N2076) );
  NOR2_X1 NOR2_608( .ZN(N2142), .A1(N2080), .A2(N2081) );
  NOR2_X1 NOR2_609( .ZN(N2145), .A1(N1272), .A2(N2082) );
  NOR2_X1 NOR2_610( .ZN(N2149), .A1(N2037), .A2(N2085) );
  NOR2_X1 NOR2_611( .ZN(N2150), .A1(N2085), .A2(N552) );
  NOR2_X1 NOR2_612( .ZN(N2151), .A1(N1947), .A2(N2085) );
  NOR2_X1 NOR2_613( .ZN(N2154), .A1(N2040), .A2(N2089) );
  NOR2_X1 NOR2_614( .ZN(N2155), .A1(N2089), .A2(N600) );
  NOR2_X1 NOR2_615( .ZN(N2156), .A1(N1951), .A2(N2089) );
  NOR2_X1 NOR2_616( .ZN(N2159), .A1(N2043), .A2(N2093) );
  NOR2_X1 NOR2_617( .ZN(N2160), .A1(N2093), .A2(N648) );
  NOR2_X1 NOR2_618( .ZN(N2161), .A1(N1955), .A2(N2093) );
  NOR2_X1 NOR2_619( .ZN(N2164), .A1(N2046), .A2(N2097) );
  NOR2_X1 NOR2_620( .ZN(N2165), .A1(N2097), .A2(N696) );
  NOR2_X1 NOR2_621( .ZN(N2166), .A1(N1959), .A2(N2097) );
  NOR2_X1 NOR2_622( .ZN(N2169), .A1(N2049), .A2(N2101) );
  NOR2_X1 NOR2_623( .ZN(N2170), .A1(N2101), .A2(N744) );
  NOR2_X1 NOR2_624( .ZN(N2171), .A1(N1963), .A2(N2101) );
  NOR2_X1 NOR2_625( .ZN(N2174), .A1(N2052), .A2(N2105) );
  NOR2_X1 NOR2_626( .ZN(N2175), .A1(N2105), .A2(N792) );
  NOR2_X1 NOR2_627( .ZN(N2176), .A1(N1967), .A2(N2105) );
  NOR2_X1 NOR2_628( .ZN(N2179), .A1(N2055), .A2(N2109) );
  NOR2_X1 NOR2_629( .ZN(N2180), .A1(N2109), .A2(N840) );
  NOR2_X1 NOR2_630( .ZN(N2181), .A1(N1971), .A2(N2109) );
  NOR2_X1 NOR2_631( .ZN(N2184), .A1(N2058), .A2(N2113) );
  NOR2_X1 NOR2_632( .ZN(N2185), .A1(N2113), .A2(N888) );
  NOR2_X1 NOR2_633( .ZN(N2186), .A1(N1975), .A2(N2113) );
  NOR2_X1 NOR2_634( .ZN(N2189), .A1(N2061), .A2(N2117) );
  NOR2_X1 NOR2_635( .ZN(N2190), .A1(N2117), .A2(N936) );
  NOR2_X1 NOR2_636( .ZN(N2191), .A1(N1979), .A2(N2117) );
  NOR2_X1 NOR2_637( .ZN(N2194), .A1(N2064), .A2(N2121) );
  NOR2_X1 NOR2_638( .ZN(N2195), .A1(N2121), .A2(N984) );
  NOR2_X1 NOR2_639( .ZN(N2196), .A1(N1983), .A2(N2121) );
  NOR2_X1 NOR2_640( .ZN(N2199), .A1(N2067), .A2(N2125) );
  NOR2_X1 NOR2_641( .ZN(N2200), .A1(N2125), .A2(N1032) );
  NOR2_X1 NOR2_642( .ZN(N2201), .A1(N1987), .A2(N2125) );
  NOR2_X1 NOR2_643( .ZN(N2204), .A1(N2070), .A2(N2129) );
  NOR2_X1 NOR2_644( .ZN(N2205), .A1(N2129), .A2(N1080) );
  NOR2_X1 NOR2_645( .ZN(N2206), .A1(N1991), .A2(N2129) );
  NOR2_X1 NOR2_646( .ZN(N2209), .A1(N2073), .A2(N2133) );
  NOR2_X1 NOR2_647( .ZN(N2210), .A1(N2133), .A2(N1128) );
  NOR2_X1 NOR2_648( .ZN(N2211), .A1(N1995), .A2(N2133) );
  NOR2_X1 NOR2_649( .ZN(N2214), .A1(N2137), .A2(N2138) );
  NOR2_X1 NOR2_650( .ZN(N2217), .A1(N2142), .A2(N2139) );
  NOR2_X1 NOR2_651( .ZN(N2221), .A1(N1272), .A2(N2145) );
  NOR2_X1 NOR2_652( .ZN(N2222), .A1(N2145), .A2(N2082) );
  NOR2_X1 NOR2_653( .ZN(N2223), .A1(N2149), .A2(N2150) );
  NOR2_X1 NOR2_654( .ZN(N2224), .A1(N2154), .A2(N2155) );
  NOR2_X1 NOR2_655( .ZN(N2227), .A1(N2159), .A2(N2160) );
  NOR2_X1 NOR2_656( .ZN(N2230), .A1(N2164), .A2(N2165) );
  NOR2_X1 NOR2_657( .ZN(N2233), .A1(N2169), .A2(N2170) );
  NOR2_X1 NOR2_658( .ZN(N2236), .A1(N2174), .A2(N2175) );
  NOR2_X1 NOR2_659( .ZN(N2239), .A1(N2179), .A2(N2180) );
  NOR2_X1 NOR2_660( .ZN(N2242), .A1(N2184), .A2(N2185) );
  NOR2_X1 NOR2_661( .ZN(N2245), .A1(N2189), .A2(N2190) );
  NOR2_X1 NOR2_662( .ZN(N2248), .A1(N2194), .A2(N2195) );
  NOR2_X1 NOR2_663( .ZN(N2251), .A1(N2199), .A2(N2200) );
  NOR2_X1 NOR2_664( .ZN(N2254), .A1(N2204), .A2(N2205) );
  NOR2_X1 NOR2_665( .ZN(N2257), .A1(N2209), .A2(N2210) );
  NOR2_X1 NOR2_666( .ZN(N2260), .A1(N2214), .A2(N2211) );
  NOR2_X1 NOR2_667( .ZN(N2264), .A1(N2142), .A2(N2217) );
  NOR2_X1 NOR2_668( .ZN(N2265), .A1(N2217), .A2(N2139) );
  NOR2_X1 NOR2_669( .ZN(N2266), .A1(N2221), .A2(N2222) );
  NOR2_X1 NOR2_670( .ZN(N2269), .A1(N2224), .A2(N2151) );
  NOR2_X1 NOR2_671( .ZN(N2273), .A1(N2227), .A2(N2156) );
  NOR2_X1 NOR2_672( .ZN(N2277), .A1(N2230), .A2(N2161) );
  NOR2_X1 NOR2_673( .ZN(N2281), .A1(N2233), .A2(N2166) );
  NOR2_X1 NOR2_674( .ZN(N2285), .A1(N2236), .A2(N2171) );
  NOR2_X1 NOR2_675( .ZN(N2289), .A1(N2239), .A2(N2176) );
  NOR2_X1 NOR2_676( .ZN(N2293), .A1(N2242), .A2(N2181) );
  NOR2_X1 NOR2_677( .ZN(N2297), .A1(N2245), .A2(N2186) );
  NOR2_X1 NOR2_678( .ZN(N2301), .A1(N2248), .A2(N2191) );
  NOR2_X1 NOR2_679( .ZN(N2305), .A1(N2251), .A2(N2196) );
  NOR2_X2 NOR2_680( .ZN(N2309), .A1(N2254), .A2(N2201) );
  NOR2_X2 NOR2_681( .ZN(N2313), .A1(N2257), .A2(N2206) );
  NOR2_X2 NOR2_682( .ZN(N2317), .A1(N2214), .A2(N2260) );
  NOR2_X2 NOR2_683( .ZN(N2318), .A1(N2260), .A2(N2211) );
  NOR2_X2 NOR2_684( .ZN(N2319), .A1(N2264), .A2(N2265) );
  NOR2_X2 NOR2_685( .ZN(N2322), .A1(N2266), .A2(N1227) );
  NOR2_X1 NOR2_686( .ZN(N2326), .A1(N2224), .A2(N2269) );
  NOR2_X1 NOR2_687( .ZN(N2327), .A1(N2269), .A2(N2151) );
  NOR2_X1 NOR2_688( .ZN(N2328), .A1(N2227), .A2(N2273) );
  NOR2_X1 NOR2_689( .ZN(N2329), .A1(N2273), .A2(N2156) );
  NOR2_X1 NOR2_690( .ZN(N2330), .A1(N2230), .A2(N2277) );
  NOR2_X1 NOR2_691( .ZN(N2331), .A1(N2277), .A2(N2161) );
  NOR2_X1 NOR2_692( .ZN(N2332), .A1(N2233), .A2(N2281) );
  NOR2_X1 NOR2_693( .ZN(N2333), .A1(N2281), .A2(N2166) );
  NOR2_X1 NOR2_694( .ZN(N2334), .A1(N2236), .A2(N2285) );
  NOR2_X1 NOR2_695( .ZN(N2335), .A1(N2285), .A2(N2171) );
  NOR2_X1 NOR2_696( .ZN(N2336), .A1(N2239), .A2(N2289) );
  NOR2_X1 NOR2_697( .ZN(N2337), .A1(N2289), .A2(N2176) );
  NOR2_X1 NOR2_698( .ZN(N2338), .A1(N2242), .A2(N2293) );
  NOR2_X1 NOR2_699( .ZN(N2339), .A1(N2293), .A2(N2181) );
  NOR2_X1 NOR2_700( .ZN(N2340), .A1(N2245), .A2(N2297) );
  NOR2_X1 NOR2_701( .ZN(N2341), .A1(N2297), .A2(N2186) );
  NOR2_X1 NOR2_702( .ZN(N2342), .A1(N2248), .A2(N2301) );
  NOR2_X1 NOR2_703( .ZN(N2343), .A1(N2301), .A2(N2191) );
  NOR2_X1 NOR2_704( .ZN(N2344), .A1(N2251), .A2(N2305) );
  NOR2_X1 NOR2_705( .ZN(N2345), .A1(N2305), .A2(N2196) );
  NOR2_X1 NOR2_706( .ZN(N2346), .A1(N2254), .A2(N2309) );
  NOR2_X1 NOR2_707( .ZN(N2347), .A1(N2309), .A2(N2201) );
  NOR2_X1 NOR2_708( .ZN(N2348), .A1(N2257), .A2(N2313) );
  NOR2_X1 NOR2_709( .ZN(N2349), .A1(N2313), .A2(N2206) );
  NOR2_X1 NOR2_710( .ZN(N2350), .A1(N2317), .A2(N2318) );
  NOR2_X1 NOR2_711( .ZN(N2353), .A1(N2319), .A2(N1179) );
  NOR2_X1 NOR2_712( .ZN(N2357), .A1(N2266), .A2(N2322) );
  NOR2_X1 NOR2_713( .ZN(N2358), .A1(N2322), .A2(N1227) );
  NOR2_X1 NOR2_714( .ZN(N2359), .A1(N2145), .A2(N2322) );
  NOR2_X1 NOR2_715( .ZN(N2362), .A1(N2326), .A2(N2327) );
  NOR2_X1 NOR2_716( .ZN(N2365), .A1(N2328), .A2(N2329) );
  NOR2_X1 NOR2_717( .ZN(N2368), .A1(N2330), .A2(N2331) );
  NOR2_X1 NOR2_718( .ZN(N2371), .A1(N2332), .A2(N2333) );
  NOR2_X1 NOR2_719( .ZN(N2374), .A1(N2334), .A2(N2335) );
  NOR2_X1 NOR2_720( .ZN(N2377), .A1(N2336), .A2(N2337) );
  NOR2_X1 NOR2_721( .ZN(N2380), .A1(N2338), .A2(N2339) );
  NOR2_X1 NOR2_722( .ZN(N2383), .A1(N2340), .A2(N2341) );
  NOR2_X1 NOR2_723( .ZN(N2386), .A1(N2342), .A2(N2343) );
  NOR2_X1 NOR2_724( .ZN(N2389), .A1(N2344), .A2(N2345) );
  NOR2_X1 NOR2_725( .ZN(N2392), .A1(N2346), .A2(N2347) );
  NOR2_X1 NOR2_726( .ZN(N2395), .A1(N2348), .A2(N2349) );
  NOR2_X1 NOR2_727( .ZN(N2398), .A1(N2350), .A2(N1131) );
  NOR2_X1 NOR2_728( .ZN(N2402), .A1(N2319), .A2(N2353) );
  NOR2_X1 NOR2_729( .ZN(N2403), .A1(N2353), .A2(N1179) );
  NOR2_X1 NOR2_730( .ZN(N2404), .A1(N2217), .A2(N2353) );
  NOR2_X1 NOR2_731( .ZN(N2407), .A1(N2357), .A2(N2358) );
  NOR2_X1 NOR2_732( .ZN(N2410), .A1(N1275), .A2(N2359) );
  NOR2_X1 NOR2_733( .ZN(N2414), .A1(N2362), .A2(N555) );
  NOR2_X1 NOR2_734( .ZN(N2418), .A1(N2365), .A2(N603) );
  NOR2_X1 NOR2_735( .ZN(N2422), .A1(N2368), .A2(N651) );
  NOR2_X1 NOR2_736( .ZN(N2426), .A1(N2371), .A2(N699) );
  NOR2_X1 NOR2_737( .ZN(N2430), .A1(N2374), .A2(N747) );
  NOR2_X1 NOR2_738( .ZN(N2434), .A1(N2377), .A2(N795) );
  NOR2_X1 NOR2_739( .ZN(N2438), .A1(N2380), .A2(N843) );
  NOR2_X1 NOR2_740( .ZN(N2442), .A1(N2383), .A2(N891) );
  NOR2_X1 NOR2_741( .ZN(N2446), .A1(N2386), .A2(N939) );
  NOR2_X1 NOR2_742( .ZN(N2450), .A1(N2389), .A2(N987) );
  NOR2_X1 NOR2_743( .ZN(N2454), .A1(N2392), .A2(N1035) );
  NOR2_X1 NOR2_744( .ZN(N2458), .A1(N2395), .A2(N1083) );
  NOR2_X1 NOR2_745( .ZN(N2462), .A1(N2350), .A2(N2398) );
  NOR2_X1 NOR2_746( .ZN(N2463), .A1(N2398), .A2(N1131) );
  NOR2_X1 NOR2_747( .ZN(N2464), .A1(N2260), .A2(N2398) );
  NOR2_X1 NOR2_748( .ZN(N2467), .A1(N2402), .A2(N2403) );
  NOR2_X1 NOR2_749( .ZN(N2470), .A1(N2407), .A2(N2404) );
  NOR2_X1 NOR2_750( .ZN(N2474), .A1(N1275), .A2(N2410) );
  NOR2_X1 NOR2_751( .ZN(N2475), .A1(N2410), .A2(N2359) );
  NOR2_X1 NOR2_752( .ZN(N2476), .A1(N2362), .A2(N2414) );
  NOR2_X1 NOR2_753( .ZN(N2477), .A1(N2414), .A2(N555) );
  NOR2_X1 NOR2_754( .ZN(N2478), .A1(N2269), .A2(N2414) );
  NOR2_X1 NOR2_755( .ZN(N2481), .A1(N2365), .A2(N2418) );
  NOR2_X1 NOR2_756( .ZN(N2482), .A1(N2418), .A2(N603) );
  NOR2_X1 NOR2_757( .ZN(N2483), .A1(N2273), .A2(N2418) );
  NOR2_X1 NOR2_758( .ZN(N2486), .A1(N2368), .A2(N2422) );
  NOR2_X1 NOR2_759( .ZN(N2487), .A1(N2422), .A2(N651) );
  NOR2_X1 NOR2_760( .ZN(N2488), .A1(N2277), .A2(N2422) );
  NOR2_X1 NOR2_761( .ZN(N2491), .A1(N2371), .A2(N2426) );
  NOR2_X1 NOR2_762( .ZN(N2492), .A1(N2426), .A2(N699) );
  NOR2_X1 NOR2_763( .ZN(N2493), .A1(N2281), .A2(N2426) );
  NOR2_X1 NOR2_764( .ZN(N2496), .A1(N2374), .A2(N2430) );
  NOR2_X1 NOR2_765( .ZN(N2497), .A1(N2430), .A2(N747) );
  NOR2_X1 NOR2_766( .ZN(N2498), .A1(N2285), .A2(N2430) );
  NOR2_X1 NOR2_767( .ZN(N2501), .A1(N2377), .A2(N2434) );
  NOR2_X1 NOR2_768( .ZN(N2502), .A1(N2434), .A2(N795) );
  NOR2_X1 NOR2_769( .ZN(N2503), .A1(N2289), .A2(N2434) );
  NOR2_X1 NOR2_770( .ZN(N2506), .A1(N2380), .A2(N2438) );
  NOR2_X1 NOR2_771( .ZN(N2507), .A1(N2438), .A2(N843) );
  NOR2_X1 NOR2_772( .ZN(N2508), .A1(N2293), .A2(N2438) );
  NOR2_X1 NOR2_773( .ZN(N2511), .A1(N2383), .A2(N2442) );
  NOR2_X1 NOR2_774( .ZN(N2512), .A1(N2442), .A2(N891) );
  NOR2_X1 NOR2_775( .ZN(N2513), .A1(N2297), .A2(N2442) );
  NOR2_X1 NOR2_776( .ZN(N2516), .A1(N2386), .A2(N2446) );
  NOR2_X1 NOR2_777( .ZN(N2517), .A1(N2446), .A2(N939) );
  NOR2_X1 NOR2_778( .ZN(N2518), .A1(N2301), .A2(N2446) );
  NOR2_X1 NOR2_779( .ZN(N2521), .A1(N2389), .A2(N2450) );
  NOR2_X1 NOR2_780( .ZN(N2522), .A1(N2450), .A2(N987) );
  NOR2_X1 NOR2_781( .ZN(N2523), .A1(N2305), .A2(N2450) );
  NOR2_X1 NOR2_782( .ZN(N2526), .A1(N2392), .A2(N2454) );
  NOR2_X1 NOR2_783( .ZN(N2527), .A1(N2454), .A2(N1035) );
  NOR2_X1 NOR2_784( .ZN(N2528), .A1(N2309), .A2(N2454) );
  NOR2_X1 NOR2_785( .ZN(N2531), .A1(N2395), .A2(N2458) );
  NOR2_X1 NOR2_786( .ZN(N2532), .A1(N2458), .A2(N1083) );
  NOR2_X1 NOR2_787( .ZN(N2533), .A1(N2313), .A2(N2458) );
  NOR2_X1 NOR2_788( .ZN(N2536), .A1(N2462), .A2(N2463) );
  NOR2_X1 NOR2_789( .ZN(N2539), .A1(N2467), .A2(N2464) );
  NOR2_X1 NOR2_790( .ZN(N2543), .A1(N2407), .A2(N2470) );
  NOR2_X1 NOR2_791( .ZN(N2544), .A1(N2470), .A2(N2404) );
  NOR2_X1 NOR2_792( .ZN(N2545), .A1(N2474), .A2(N2475) );
  NOR2_X1 NOR2_793( .ZN(N2548), .A1(N2476), .A2(N2477) );
  NOR2_X1 NOR2_794( .ZN(N2549), .A1(N2481), .A2(N2482) );
  NOR2_X1 NOR2_795( .ZN(N2552), .A1(N2486), .A2(N2487) );
  NOR2_X1 NOR2_796( .ZN(N2555), .A1(N2491), .A2(N2492) );
  NOR2_X1 NOR2_797( .ZN(N2558), .A1(N2496), .A2(N2497) );
  NOR2_X1 NOR2_798( .ZN(N2561), .A1(N2501), .A2(N2502) );
  NOR2_X1 NOR2_799( .ZN(N2564), .A1(N2506), .A2(N2507) );
  NOR2_X1 NOR2_800( .ZN(N2567), .A1(N2511), .A2(N2512) );
  NOR2_X1 NOR2_801( .ZN(N2570), .A1(N2516), .A2(N2517) );
  NOR2_X1 NOR2_802( .ZN(N2573), .A1(N2521), .A2(N2522) );
  NOR2_X1 NOR2_803( .ZN(N2576), .A1(N2526), .A2(N2527) );
  NOR2_X1 NOR2_804( .ZN(N2579), .A1(N2531), .A2(N2532) );
  NOR2_X1 NOR2_805( .ZN(N2582), .A1(N2536), .A2(N2533) );
  NOR2_X1 NOR2_806( .ZN(N2586), .A1(N2467), .A2(N2539) );
  NOR2_X1 NOR2_807( .ZN(N2587), .A1(N2539), .A2(N2464) );
  NOR2_X1 NOR2_808( .ZN(N2588), .A1(N2543), .A2(N2544) );
  NOR2_X1 NOR2_809( .ZN(N2591), .A1(N2545), .A2(N1230) );
  NOR2_X1 NOR2_810( .ZN(N2595), .A1(N2549), .A2(N2478) );
  NOR2_X1 NOR2_811( .ZN(N2599), .A1(N2552), .A2(N2483) );
  NOR2_X1 NOR2_812( .ZN(N2603), .A1(N2555), .A2(N2488) );
  NOR2_X1 NOR2_813( .ZN(N2607), .A1(N2558), .A2(N2493) );
  NOR2_X1 NOR2_814( .ZN(N2611), .A1(N2561), .A2(N2498) );
  NOR2_X1 NOR2_815( .ZN(N2615), .A1(N2564), .A2(N2503) );
  NOR2_X1 NOR2_816( .ZN(N2619), .A1(N2567), .A2(N2508) );
  NOR2_X1 NOR2_817( .ZN(N2623), .A1(N2570), .A2(N2513) );
  NOR2_X1 NOR2_818( .ZN(N2627), .A1(N2573), .A2(N2518) );
  NOR2_X1 NOR2_819( .ZN(N2631), .A1(N2576), .A2(N2523) );
  NOR2_X1 NOR2_820( .ZN(N2635), .A1(N2579), .A2(N2528) );
  NOR2_X1 NOR2_821( .ZN(N2639), .A1(N2536), .A2(N2582) );
  NOR2_X1 NOR2_822( .ZN(N2640), .A1(N2582), .A2(N2533) );
  NOR2_X1 NOR2_823( .ZN(N2641), .A1(N2586), .A2(N2587) );
  NOR2_X1 NOR2_824( .ZN(N2644), .A1(N2588), .A2(N1182) );
  NOR2_X1 NOR2_825( .ZN(N2648), .A1(N2545), .A2(N2591) );
  NOR2_X1 NOR2_826( .ZN(N2649), .A1(N2591), .A2(N1230) );
  NOR2_X1 NOR2_827( .ZN(N2650), .A1(N2410), .A2(N2591) );
  NOR2_X1 NOR2_828( .ZN(N2653), .A1(N2549), .A2(N2595) );
  NOR2_X1 NOR2_829( .ZN(N2654), .A1(N2595), .A2(N2478) );
  NOR2_X1 NOR2_830( .ZN(N2655), .A1(N2552), .A2(N2599) );
  NOR2_X1 NOR2_831( .ZN(N2656), .A1(N2599), .A2(N2483) );
  NOR2_X1 NOR2_832( .ZN(N2657), .A1(N2555), .A2(N2603) );
  NOR2_X1 NOR2_833( .ZN(N2658), .A1(N2603), .A2(N2488) );
  NOR2_X1 NOR2_834( .ZN(N2659), .A1(N2558), .A2(N2607) );
  NOR2_X1 NOR2_835( .ZN(N2660), .A1(N2607), .A2(N2493) );
  NOR2_X1 NOR2_836( .ZN(N2661), .A1(N2561), .A2(N2611) );
  NOR2_X1 NOR2_837( .ZN(N2662), .A1(N2611), .A2(N2498) );
  NOR2_X1 NOR2_838( .ZN(N2663), .A1(N2564), .A2(N2615) );
  NOR2_X1 NOR2_839( .ZN(N2664), .A1(N2615), .A2(N2503) );
  NOR2_X1 NOR2_840( .ZN(N2665), .A1(N2567), .A2(N2619) );
  NOR2_X1 NOR2_841( .ZN(N2666), .A1(N2619), .A2(N2508) );
  NOR2_X1 NOR2_842( .ZN(N2667), .A1(N2570), .A2(N2623) );
  NOR2_X1 NOR2_843( .ZN(N2668), .A1(N2623), .A2(N2513) );
  NOR2_X1 NOR2_844( .ZN(N2669), .A1(N2573), .A2(N2627) );
  NOR2_X1 NOR2_845( .ZN(N2670), .A1(N2627), .A2(N2518) );
  NOR2_X1 NOR2_846( .ZN(N2671), .A1(N2576), .A2(N2631) );
  NOR2_X1 NOR2_847( .ZN(N2672), .A1(N2631), .A2(N2523) );
  NOR2_X1 NOR2_848( .ZN(N2673), .A1(N2579), .A2(N2635) );
  NOR2_X1 NOR2_849( .ZN(N2674), .A1(N2635), .A2(N2528) );
  NOR2_X1 NOR2_850( .ZN(N2675), .A1(N2639), .A2(N2640) );
  NOR2_X1 NOR2_851( .ZN(N2678), .A1(N2641), .A2(N1134) );
  NOR2_X1 NOR2_852( .ZN(N2682), .A1(N2588), .A2(N2644) );
  NOR2_X1 NOR2_853( .ZN(N2683), .A1(N2644), .A2(N1182) );
  NOR2_X1 NOR2_854( .ZN(N2684), .A1(N2470), .A2(N2644) );
  NOR2_X1 NOR2_855( .ZN(N2687), .A1(N2648), .A2(N2649) );
  NOR2_X1 NOR2_856( .ZN(N2690), .A1(N1278), .A2(N2650) );
  NOR2_X1 NOR2_857( .ZN(N2694), .A1(N2653), .A2(N2654) );
  NOR2_X1 NOR2_858( .ZN(N2697), .A1(N2655), .A2(N2656) );
  NOR2_X1 NOR2_859( .ZN(N2700), .A1(N2657), .A2(N2658) );
  NOR2_X1 NOR2_860( .ZN(N2703), .A1(N2659), .A2(N2660) );
  NOR2_X1 NOR2_861( .ZN(N2706), .A1(N2661), .A2(N2662) );
  NOR2_X1 NOR2_862( .ZN(N2709), .A1(N2663), .A2(N2664) );
  NOR2_X1 NOR2_863( .ZN(N2712), .A1(N2665), .A2(N2666) );
  NOR2_X1 NOR2_864( .ZN(N2715), .A1(N2667), .A2(N2668) );
  NOR2_X1 NOR2_865( .ZN(N2718), .A1(N2669), .A2(N2670) );
  NOR2_X1 NOR2_866( .ZN(N2721), .A1(N2671), .A2(N2672) );
  NOR2_X1 NOR2_867( .ZN(N2724), .A1(N2673), .A2(N2674) );
  NOR2_X1 NOR2_868( .ZN(N2727), .A1(N2675), .A2(N1086) );
  NOR2_X1 NOR2_869( .ZN(N2731), .A1(N2641), .A2(N2678) );
  NOR2_X1 NOR2_870( .ZN(N2732), .A1(N2678), .A2(N1134) );
  NOR2_X1 NOR2_871( .ZN(N2733), .A1(N2539), .A2(N2678) );
  NOR2_X1 NOR2_872( .ZN(N2736), .A1(N2682), .A2(N2683) );
  NOR2_X1 NOR2_873( .ZN(N2739), .A1(N2687), .A2(N2684) );
  NOR2_X1 NOR2_874( .ZN(N2743), .A1(N1278), .A2(N2690) );
  NOR2_X1 NOR2_875( .ZN(N2744), .A1(N2690), .A2(N2650) );
  NOR2_X1 NOR2_876( .ZN(N2745), .A1(N2694), .A2(N558) );
  NOR2_X1 NOR2_877( .ZN(N2749), .A1(N2697), .A2(N606) );
  NOR2_X1 NOR2_878( .ZN(N2753), .A1(N2700), .A2(N654) );
  NOR2_X1 NOR2_879( .ZN(N2757), .A1(N2703), .A2(N702) );
  NOR2_X1 NOR2_880( .ZN(N2761), .A1(N2706), .A2(N750) );
  NOR2_X1 NOR2_881( .ZN(N2765), .A1(N2709), .A2(N798) );
  NOR2_X1 NOR2_882( .ZN(N2769), .A1(N2712), .A2(N846) );
  NOR2_X1 NOR2_883( .ZN(N2773), .A1(N2715), .A2(N894) );
  NOR2_X1 NOR2_884( .ZN(N2777), .A1(N2718), .A2(N942) );
  NOR2_X1 NOR2_885( .ZN(N2781), .A1(N2721), .A2(N990) );
  NOR2_X1 NOR2_886( .ZN(N2785), .A1(N2724), .A2(N1038) );
  NOR2_X1 NOR2_887( .ZN(N2789), .A1(N2675), .A2(N2727) );
  NOR2_X1 NOR2_888( .ZN(N2790), .A1(N2727), .A2(N1086) );
  NOR2_X1 NOR2_889( .ZN(N2791), .A1(N2582), .A2(N2727) );
  NOR2_X1 NOR2_890( .ZN(N2794), .A1(N2731), .A2(N2732) );
  NOR2_X1 NOR2_891( .ZN(N2797), .A1(N2736), .A2(N2733) );
  NOR2_X1 NOR2_892( .ZN(N2801), .A1(N2687), .A2(N2739) );
  NOR2_X1 NOR2_893( .ZN(N2802), .A1(N2739), .A2(N2684) );
  NOR2_X1 NOR2_894( .ZN(N2803), .A1(N2743), .A2(N2744) );
  NOR2_X1 NOR2_895( .ZN(N2806), .A1(N2694), .A2(N2745) );
  NOR2_X1 NOR2_896( .ZN(N2807), .A1(N2745), .A2(N558) );
  NOR2_X1 NOR2_897( .ZN(N2808), .A1(N2595), .A2(N2745) );
  NOR2_X1 NOR2_898( .ZN(N2811), .A1(N2697), .A2(N2749) );
  NOR2_X1 NOR2_899( .ZN(N2812), .A1(N2749), .A2(N606) );
  NOR2_X1 NOR2_900( .ZN(N2813), .A1(N2599), .A2(N2749) );
  NOR2_X1 NOR2_901( .ZN(N2816), .A1(N2700), .A2(N2753) );
  NOR2_X1 NOR2_902( .ZN(N2817), .A1(N2753), .A2(N654) );
  NOR2_X1 NOR2_903( .ZN(N2818), .A1(N2603), .A2(N2753) );
  NOR2_X1 NOR2_904( .ZN(N2821), .A1(N2703), .A2(N2757) );
  NOR2_X1 NOR2_905( .ZN(N2822), .A1(N2757), .A2(N702) );
  NOR2_X1 NOR2_906( .ZN(N2823), .A1(N2607), .A2(N2757) );
  NOR2_X1 NOR2_907( .ZN(N2826), .A1(N2706), .A2(N2761) );
  NOR2_X1 NOR2_908( .ZN(N2827), .A1(N2761), .A2(N750) );
  NOR2_X1 NOR2_909( .ZN(N2828), .A1(N2611), .A2(N2761) );
  NOR2_X1 NOR2_910( .ZN(N2831), .A1(N2709), .A2(N2765) );
  NOR2_X1 NOR2_911( .ZN(N2832), .A1(N2765), .A2(N798) );
  NOR2_X1 NOR2_912( .ZN(N2833), .A1(N2615), .A2(N2765) );
  NOR2_X1 NOR2_913( .ZN(N2836), .A1(N2712), .A2(N2769) );
  NOR2_X1 NOR2_914( .ZN(N2837), .A1(N2769), .A2(N846) );
  NOR2_X1 NOR2_915( .ZN(N2838), .A1(N2619), .A2(N2769) );
  NOR2_X1 NOR2_916( .ZN(N2841), .A1(N2715), .A2(N2773) );
  NOR2_X1 NOR2_917( .ZN(N2842), .A1(N2773), .A2(N894) );
  NOR2_X1 NOR2_918( .ZN(N2843), .A1(N2623), .A2(N2773) );
  NOR2_X1 NOR2_919( .ZN(N2846), .A1(N2718), .A2(N2777) );
  NOR2_X1 NOR2_920( .ZN(N2847), .A1(N2777), .A2(N942) );
  NOR2_X1 NOR2_921( .ZN(N2848), .A1(N2627), .A2(N2777) );
  NOR2_X1 NOR2_922( .ZN(N2851), .A1(N2721), .A2(N2781) );
  NOR2_X1 NOR2_923( .ZN(N2852), .A1(N2781), .A2(N990) );
  NOR2_X1 NOR2_924( .ZN(N2853), .A1(N2631), .A2(N2781) );
  NOR2_X1 NOR2_925( .ZN(N2856), .A1(N2724), .A2(N2785) );
  NOR2_X1 NOR2_926( .ZN(N2857), .A1(N2785), .A2(N1038) );
  NOR2_X1 NOR2_927( .ZN(N2858), .A1(N2635), .A2(N2785) );
  NOR2_X1 NOR2_928( .ZN(N2861), .A1(N2789), .A2(N2790) );
  NOR2_X1 NOR2_929( .ZN(N2864), .A1(N2794), .A2(N2791) );
  NOR2_X1 NOR2_930( .ZN(N2868), .A1(N2736), .A2(N2797) );
  NOR2_X1 NOR2_931( .ZN(N2869), .A1(N2797), .A2(N2733) );
  NOR2_X1 NOR2_932( .ZN(N2870), .A1(N2801), .A2(N2802) );
  NOR2_X1 NOR2_933( .ZN(N2873), .A1(N2803), .A2(N1233) );
  NOR2_X1 NOR2_934( .ZN(N2877), .A1(N2806), .A2(N2807) );
  NOR2_X1 NOR2_935( .ZN(N2878), .A1(N2811), .A2(N2812) );
  NOR2_X1 NOR2_936( .ZN(N2881), .A1(N2816), .A2(N2817) );
  NOR2_X1 NOR2_937( .ZN(N2884), .A1(N2821), .A2(N2822) );
  NOR2_X1 NOR2_938( .ZN(N2887), .A1(N2826), .A2(N2827) );
  NOR2_X1 NOR2_939( .ZN(N2890), .A1(N2831), .A2(N2832) );
  NOR2_X1 NOR2_940( .ZN(N2893), .A1(N2836), .A2(N2837) );
  NOR2_X1 NOR2_941( .ZN(N2896), .A1(N2841), .A2(N2842) );
  NOR2_X1 NOR2_942( .ZN(N2899), .A1(N2846), .A2(N2847) );
  NOR2_X1 NOR2_943( .ZN(N2902), .A1(N2851), .A2(N2852) );
  NOR2_X1 NOR2_944( .ZN(N2905), .A1(N2856), .A2(N2857) );
  NOR2_X1 NOR2_945( .ZN(N2908), .A1(N2861), .A2(N2858) );
  NOR2_X1 NOR2_946( .ZN(N2912), .A1(N2794), .A2(N2864) );
  NOR2_X1 NOR2_947( .ZN(N2913), .A1(N2864), .A2(N2791) );
  NOR2_X1 NOR2_948( .ZN(N2914), .A1(N2868), .A2(N2869) );
  NOR2_X1 NOR2_949( .ZN(N2917), .A1(N2870), .A2(N1185) );
  NOR2_X1 NOR2_950( .ZN(N2921), .A1(N2803), .A2(N2873) );
  NOR2_X1 NOR2_951( .ZN(N2922), .A1(N2873), .A2(N1233) );
  NOR2_X1 NOR2_952( .ZN(N2923), .A1(N2690), .A2(N2873) );
  NOR2_X1 NOR2_953( .ZN(N2926), .A1(N2878), .A2(N2808) );
  NOR2_X1 NOR2_954( .ZN(N2930), .A1(N2881), .A2(N2813) );
  NOR2_X1 NOR2_955( .ZN(N2934), .A1(N2884), .A2(N2818) );
  NOR2_X1 NOR2_956( .ZN(N2938), .A1(N2887), .A2(N2823) );
  NOR2_X1 NOR2_957( .ZN(N2942), .A1(N2890), .A2(N2828) );
  NOR2_X1 NOR2_958( .ZN(N2946), .A1(N2893), .A2(N2833) );
  NOR2_X1 NOR2_959( .ZN(N2950), .A1(N2896), .A2(N2838) );
  NOR2_X1 NOR2_960( .ZN(N2954), .A1(N2899), .A2(N2843) );
  NOR2_X1 NOR2_961( .ZN(N2958), .A1(N2902), .A2(N2848) );
  NOR2_X1 NOR2_962( .ZN(N2962), .A1(N2905), .A2(N2853) );
  NOR2_X1 NOR2_963( .ZN(N2966), .A1(N2861), .A2(N2908) );
  NOR2_X1 NOR2_964( .ZN(N2967), .A1(N2908), .A2(N2858) );
  NOR2_X1 NOR2_965( .ZN(N2968), .A1(N2912), .A2(N2913) );
  NOR2_X1 NOR2_966( .ZN(N2971), .A1(N2914), .A2(N1137) );
  NOR2_X1 NOR2_967( .ZN(N2975), .A1(N2870), .A2(N2917) );
  NOR2_X1 NOR2_968( .ZN(N2976), .A1(N2917), .A2(N1185) );
  NOR2_X1 NOR2_969( .ZN(N2977), .A1(N2739), .A2(N2917) );
  NOR2_X1 NOR2_970( .ZN(N2980), .A1(N2921), .A2(N2922) );
  NOR2_X1 NOR2_971( .ZN(N2983), .A1(N1281), .A2(N2923) );
  NOR2_X1 NOR2_972( .ZN(N2987), .A1(N2878), .A2(N2926) );
  NOR2_X1 NOR2_973( .ZN(N2988), .A1(N2926), .A2(N2808) );
  NOR2_X1 NOR2_974( .ZN(N2989), .A1(N2881), .A2(N2930) );
  NOR2_X1 NOR2_975( .ZN(N2990), .A1(N2930), .A2(N2813) );
  NOR2_X1 NOR2_976( .ZN(N2991), .A1(N2884), .A2(N2934) );
  NOR2_X1 NOR2_977( .ZN(N2992), .A1(N2934), .A2(N2818) );
  NOR2_X1 NOR2_978( .ZN(N2993), .A1(N2887), .A2(N2938) );
  NOR2_X1 NOR2_979( .ZN(N2994), .A1(N2938), .A2(N2823) );
  NOR2_X1 NOR2_980( .ZN(N2995), .A1(N2890), .A2(N2942) );
  NOR2_X1 NOR2_981( .ZN(N2996), .A1(N2942), .A2(N2828) );
  NOR2_X1 NOR2_982( .ZN(N2997), .A1(N2893), .A2(N2946) );
  NOR2_X1 NOR2_983( .ZN(N2998), .A1(N2946), .A2(N2833) );
  NOR2_X1 NOR2_984( .ZN(N2999), .A1(N2896), .A2(N2950) );
  NOR2_X1 NOR2_985( .ZN(N3000), .A1(N2950), .A2(N2838) );
  NOR2_X1 NOR2_986( .ZN(N3001), .A1(N2899), .A2(N2954) );
  NOR2_X1 NOR2_987( .ZN(N3002), .A1(N2954), .A2(N2843) );
  NOR2_X1 NOR2_988( .ZN(N3003), .A1(N2902), .A2(N2958) );
  NOR2_X1 NOR2_989( .ZN(N3004), .A1(N2958), .A2(N2848) );
  NOR2_X1 NOR2_990( .ZN(N3005), .A1(N2905), .A2(N2962) );
  NOR2_X1 NOR2_991( .ZN(N3006), .A1(N2962), .A2(N2853) );
  NOR2_X1 NOR2_992( .ZN(N3007), .A1(N2966), .A2(N2967) );
  NOR2_X1 NOR2_993( .ZN(N3010), .A1(N2968), .A2(N1089) );
  NOR2_X1 NOR2_994( .ZN(N3014), .A1(N2914), .A2(N2971) );
  NOR2_X1 NOR2_995( .ZN(N3015), .A1(N2971), .A2(N1137) );
  NOR2_X1 NOR2_996( .ZN(N3016), .A1(N2797), .A2(N2971) );
  NOR2_X1 NOR2_997( .ZN(N3019), .A1(N2975), .A2(N2976) );
  NOR2_X1 NOR2_998( .ZN(N3022), .A1(N2980), .A2(N2977) );
  NOR2_X1 NOR2_999( .ZN(N3026), .A1(N1281), .A2(N2983) );
  NOR2_X1 NOR2_1000( .ZN(N3027), .A1(N2983), .A2(N2923) );
  NOR2_X1 NOR2_1001( .ZN(N3028), .A1(N2987), .A2(N2988) );
  NOR2_X1 NOR2_1002( .ZN(N3031), .A1(N2989), .A2(N2990) );
  NOR2_X1 NOR2_1003( .ZN(N3034), .A1(N2991), .A2(N2992) );
  NOR2_X1 NOR2_1004( .ZN(N3037), .A1(N2993), .A2(N2994) );
  NOR2_X1 NOR2_1005( .ZN(N3040), .A1(N2995), .A2(N2996) );
  NOR2_X1 NOR2_1006( .ZN(N3043), .A1(N2997), .A2(N2998) );
  NOR2_X1 NOR2_1007( .ZN(N3046), .A1(N2999), .A2(N3000) );
  NOR2_X1 NOR2_1008( .ZN(N3049), .A1(N3001), .A2(N3002) );
  NOR2_X1 NOR2_1009( .ZN(N3052), .A1(N3003), .A2(N3004) );
  NOR2_X1 NOR2_1010( .ZN(N3055), .A1(N3005), .A2(N3006) );
  NOR2_X1 NOR2_1011( .ZN(N3058), .A1(N3007), .A2(N1041) );
  NOR2_X1 NOR2_1012( .ZN(N3062), .A1(N2968), .A2(N3010) );
  NOR2_X1 NOR2_1013( .ZN(N3063), .A1(N3010), .A2(N1089) );
  NOR2_X1 NOR2_1014( .ZN(N3064), .A1(N2864), .A2(N3010) );
  NOR2_X1 NOR2_1015( .ZN(N3067), .A1(N3014), .A2(N3015) );
  NOR2_X1 NOR2_1016( .ZN(N3070), .A1(N3019), .A2(N3016) );
  NOR2_X1 NOR2_1017( .ZN(N3074), .A1(N2980), .A2(N3022) );
  NOR2_X1 NOR2_1018( .ZN(N3075), .A1(N3022), .A2(N2977) );
  NOR2_X1 NOR2_1019( .ZN(N3076), .A1(N3026), .A2(N3027) );
  NOR2_X1 NOR2_1020( .ZN(N3079), .A1(N3028), .A2(N561) );
  NOR2_X1 NOR2_1021( .ZN(N3083), .A1(N3031), .A2(N609) );
  NOR2_X1 NOR2_1022( .ZN(N3087), .A1(N3034), .A2(N657) );
  NOR2_X1 NOR2_1023( .ZN(N3091), .A1(N3037), .A2(N705) );
  NOR2_X1 NOR2_1024( .ZN(N3095), .A1(N3040), .A2(N753) );
  NOR2_X1 NOR2_1025( .ZN(N3099), .A1(N3043), .A2(N801) );
  NOR2_X1 NOR2_1026( .ZN(N3103), .A1(N3046), .A2(N849) );
  NOR2_X1 NOR2_1027( .ZN(N3107), .A1(N3049), .A2(N897) );
  NOR2_X1 NOR2_1028( .ZN(N3111), .A1(N3052), .A2(N945) );
  NOR2_X1 NOR2_1029( .ZN(N3115), .A1(N3055), .A2(N993) );
  NOR2_X1 NOR2_1030( .ZN(N3119), .A1(N3007), .A2(N3058) );
  NOR2_X1 NOR2_1031( .ZN(N3120), .A1(N3058), .A2(N1041) );
  NOR2_X1 NOR2_1032( .ZN(N3121), .A1(N2908), .A2(N3058) );
  NOR2_X1 NOR2_1033( .ZN(N3124), .A1(N3062), .A2(N3063) );
  NOR2_X1 NOR2_1034( .ZN(N3127), .A1(N3067), .A2(N3064) );
  NOR2_X1 NOR2_1035( .ZN(N3131), .A1(N3019), .A2(N3070) );
  NOR2_X1 NOR2_1036( .ZN(N3132), .A1(N3070), .A2(N3016) );
  NOR2_X1 NOR2_1037( .ZN(N3133), .A1(N3074), .A2(N3075) );
  NOR2_X1 NOR2_1038( .ZN(N3136), .A1(N3076), .A2(N1236) );
  NOR2_X1 NOR2_1039( .ZN(N3140), .A1(N3028), .A2(N3079) );
  NOR2_X1 NOR2_1040( .ZN(N3141), .A1(N3079), .A2(N561) );
  NOR2_X1 NOR2_1041( .ZN(N3142), .A1(N2926), .A2(N3079) );
  NOR2_X1 NOR2_1042( .ZN(N3145), .A1(N3031), .A2(N3083) );
  NOR2_X1 NOR2_1043( .ZN(N3146), .A1(N3083), .A2(N609) );
  NOR2_X1 NOR2_1044( .ZN(N3147), .A1(N2930), .A2(N3083) );
  NOR2_X1 NOR2_1045( .ZN(N3150), .A1(N3034), .A2(N3087) );
  NOR2_X1 NOR2_1046( .ZN(N3151), .A1(N3087), .A2(N657) );
  NOR2_X1 NOR2_1047( .ZN(N3152), .A1(N2934), .A2(N3087) );
  NOR2_X1 NOR2_1048( .ZN(N3155), .A1(N3037), .A2(N3091) );
  NOR2_X1 NOR2_1049( .ZN(N3156), .A1(N3091), .A2(N705) );
  NOR2_X1 NOR2_1050( .ZN(N3157), .A1(N2938), .A2(N3091) );
  NOR2_X1 NOR2_1051( .ZN(N3160), .A1(N3040), .A2(N3095) );
  NOR2_X1 NOR2_1052( .ZN(N3161), .A1(N3095), .A2(N753) );
  NOR2_X1 NOR2_1053( .ZN(N3162), .A1(N2942), .A2(N3095) );
  NOR2_X1 NOR2_1054( .ZN(N3165), .A1(N3043), .A2(N3099) );
  NOR2_X1 NOR2_1055( .ZN(N3166), .A1(N3099), .A2(N801) );
  NOR2_X1 NOR2_1056( .ZN(N3167), .A1(N2946), .A2(N3099) );
  NOR2_X1 NOR2_1057( .ZN(N3170), .A1(N3046), .A2(N3103) );
  NOR2_X1 NOR2_1058( .ZN(N3171), .A1(N3103), .A2(N849) );
  NOR2_X1 NOR2_1059( .ZN(N3172), .A1(N2950), .A2(N3103) );
  NOR2_X1 NOR2_1060( .ZN(N3175), .A1(N3049), .A2(N3107) );
  NOR2_X1 NOR2_1061( .ZN(N3176), .A1(N3107), .A2(N897) );
  NOR2_X1 NOR2_1062( .ZN(N3177), .A1(N2954), .A2(N3107) );
  NOR2_X1 NOR2_1063( .ZN(N3180), .A1(N3052), .A2(N3111) );
  NOR2_X1 NOR2_1064( .ZN(N3181), .A1(N3111), .A2(N945) );
  NOR2_X1 NOR2_1065( .ZN(N3182), .A1(N2958), .A2(N3111) );
  NOR2_X1 NOR2_1066( .ZN(N3185), .A1(N3055), .A2(N3115) );
  NOR2_X1 NOR2_1067( .ZN(N3186), .A1(N3115), .A2(N993) );
  NOR2_X1 NOR2_1068( .ZN(N3187), .A1(N2962), .A2(N3115) );
  NOR2_X1 NOR2_1069( .ZN(N3190), .A1(N3119), .A2(N3120) );
  NOR2_X1 NOR2_1070( .ZN(N3193), .A1(N3124), .A2(N3121) );
  NOR2_X1 NOR2_1071( .ZN(N3197), .A1(N3067), .A2(N3127) );
  NOR2_X1 NOR2_1072( .ZN(N3198), .A1(N3127), .A2(N3064) );
  NOR2_X1 NOR2_1073( .ZN(N3199), .A1(N3131), .A2(N3132) );
  NOR2_X1 NOR2_1074( .ZN(N3202), .A1(N3133), .A2(N1188) );
  NOR2_X1 NOR2_1075( .ZN(N3206), .A1(N3076), .A2(N3136) );
  NOR2_X1 NOR2_1076( .ZN(N3207), .A1(N3136), .A2(N1236) );
  NOR2_X1 NOR2_1077( .ZN(N3208), .A1(N2983), .A2(N3136) );
  NOR2_X1 NOR2_1078( .ZN(N3211), .A1(N3140), .A2(N3141) );
  NOR2_X1 NOR2_1079( .ZN(N3212), .A1(N3145), .A2(N3146) );
  NOR2_X1 NOR2_1080( .ZN(N3215), .A1(N3150), .A2(N3151) );
  NOR2_X1 NOR2_1081( .ZN(N3218), .A1(N3155), .A2(N3156) );
  NOR2_X1 NOR2_1082( .ZN(N3221), .A1(N3160), .A2(N3161) );
  NOR2_X1 NOR2_1083( .ZN(N3224), .A1(N3165), .A2(N3166) );
  NOR2_X1 NOR2_1084( .ZN(N3227), .A1(N3170), .A2(N3171) );
  NOR2_X1 NOR2_1085( .ZN(N3230), .A1(N3175), .A2(N3176) );
  NOR2_X1 NOR2_1086( .ZN(N3233), .A1(N3180), .A2(N3181) );
  NOR2_X1 NOR2_1087( .ZN(N3236), .A1(N3185), .A2(N3186) );
  NOR2_X1 NOR2_1088( .ZN(N3239), .A1(N3190), .A2(N3187) );
  NOR2_X1 NOR2_1089( .ZN(N3243), .A1(N3124), .A2(N3193) );
  NOR2_X1 NOR2_1090( .ZN(N3244), .A1(N3193), .A2(N3121) );
  NOR2_X1 NOR2_1091( .ZN(N3245), .A1(N3197), .A2(N3198) );
  NOR2_X1 NOR2_1092( .ZN(N3248), .A1(N3199), .A2(N1140) );
  NOR2_X1 NOR2_1093( .ZN(N3252), .A1(N3133), .A2(N3202) );
  NOR2_X1 NOR2_1094( .ZN(N3253), .A1(N3202), .A2(N1188) );
  NOR2_X1 NOR2_1095( .ZN(N3254), .A1(N3022), .A2(N3202) );
  NOR2_X1 NOR2_1096( .ZN(N3257), .A1(N3206), .A2(N3207) );
  NOR2_X1 NOR2_1097( .ZN(N3260), .A1(N1284), .A2(N3208) );
  NOR2_X1 NOR2_1098( .ZN(N3264), .A1(N3212), .A2(N3142) );
  NOR2_X1 NOR2_1099( .ZN(N3268), .A1(N3215), .A2(N3147) );
  NOR2_X1 NOR2_1100( .ZN(N3272), .A1(N3218), .A2(N3152) );
  NOR2_X1 NOR2_1101( .ZN(N3276), .A1(N3221), .A2(N3157) );
  NOR2_X1 NOR2_1102( .ZN(N3280), .A1(N3224), .A2(N3162) );
  NOR2_X1 NOR2_1103( .ZN(N3284), .A1(N3227), .A2(N3167) );
  NOR2_X1 NOR2_1104( .ZN(N3288), .A1(N3230), .A2(N3172) );
  NOR2_X1 NOR2_1105( .ZN(N3292), .A1(N3233), .A2(N3177) );
  NOR2_X1 NOR2_1106( .ZN(N3296), .A1(N3236), .A2(N3182) );
  NOR2_X1 NOR2_1107( .ZN(N3300), .A1(N3190), .A2(N3239) );
  NOR2_X1 NOR2_1108( .ZN(N3301), .A1(N3239), .A2(N3187) );
  NOR2_X1 NOR2_1109( .ZN(N3302), .A1(N3243), .A2(N3244) );
  NOR2_X1 NOR2_1110( .ZN(N3305), .A1(N3245), .A2(N1092) );
  NOR2_X1 NOR2_1111( .ZN(N3309), .A1(N3199), .A2(N3248) );
  NOR2_X1 NOR2_1112( .ZN(N3310), .A1(N3248), .A2(N1140) );
  NOR2_X1 NOR2_1113( .ZN(N3311), .A1(N3070), .A2(N3248) );
  NOR2_X1 NOR2_1114( .ZN(N3314), .A1(N3252), .A2(N3253) );
  NOR2_X1 NOR2_1115( .ZN(N3317), .A1(N3257), .A2(N3254) );
  NOR2_X1 NOR2_1116( .ZN(N3321), .A1(N1284), .A2(N3260) );
  NOR2_X1 NOR2_1117( .ZN(N3322), .A1(N3260), .A2(N3208) );
  NOR2_X1 NOR2_1118( .ZN(N3323), .A1(N3212), .A2(N3264) );
  NOR2_X1 NOR2_1119( .ZN(N3324), .A1(N3264), .A2(N3142) );
  NOR2_X1 NOR2_1120( .ZN(N3325), .A1(N3215), .A2(N3268) );
  NOR2_X1 NOR2_1121( .ZN(N3326), .A1(N3268), .A2(N3147) );
  NOR2_X1 NOR2_1122( .ZN(N3327), .A1(N3218), .A2(N3272) );
  NOR2_X1 NOR2_1123( .ZN(N3328), .A1(N3272), .A2(N3152) );
  NOR2_X1 NOR2_1124( .ZN(N3329), .A1(N3221), .A2(N3276) );
  NOR2_X1 NOR2_1125( .ZN(N3330), .A1(N3276), .A2(N3157) );
  NOR2_X1 NOR2_1126( .ZN(N3331), .A1(N3224), .A2(N3280) );
  NOR2_X1 NOR2_1127( .ZN(N3332), .A1(N3280), .A2(N3162) );
  NOR2_X1 NOR2_1128( .ZN(N3333), .A1(N3227), .A2(N3284) );
  NOR2_X1 NOR2_1129( .ZN(N3334), .A1(N3284), .A2(N3167) );
  NOR2_X1 NOR2_1130( .ZN(N3335), .A1(N3230), .A2(N3288) );
  NOR2_X1 NOR2_1131( .ZN(N3336), .A1(N3288), .A2(N3172) );
  NOR2_X1 NOR2_1132( .ZN(N3337), .A1(N3233), .A2(N3292) );
  NOR2_X1 NOR2_1133( .ZN(N3338), .A1(N3292), .A2(N3177) );
  NOR2_X1 NOR2_1134( .ZN(N3339), .A1(N3236), .A2(N3296) );
  NOR2_X1 NOR2_1135( .ZN(N3340), .A1(N3296), .A2(N3182) );
  NOR2_X1 NOR2_1136( .ZN(N3341), .A1(N3300), .A2(N3301) );
  NOR2_X1 NOR2_1137( .ZN(N3344), .A1(N3302), .A2(N1044) );
  NOR2_X1 NOR2_1138( .ZN(N3348), .A1(N3245), .A2(N3305) );
  NOR2_X1 NOR2_1139( .ZN(N3349), .A1(N3305), .A2(N1092) );
  NOR2_X1 NOR2_1140( .ZN(N3350), .A1(N3127), .A2(N3305) );
  NOR2_X1 NOR2_1141( .ZN(N3353), .A1(N3309), .A2(N3310) );
  NOR2_X1 NOR2_1142( .ZN(N3356), .A1(N3314), .A2(N3311) );
  NOR2_X1 NOR2_1143( .ZN(N3360), .A1(N3257), .A2(N3317) );
  NOR2_X1 NOR2_1144( .ZN(N3361), .A1(N3317), .A2(N3254) );
  NOR2_X1 NOR2_1145( .ZN(N3362), .A1(N3321), .A2(N3322) );
  NOR2_X1 NOR2_1146( .ZN(N3365), .A1(N3323), .A2(N3324) );
  NOR2_X1 NOR2_1147( .ZN(N3368), .A1(N3325), .A2(N3326) );
  NOR2_X1 NOR2_1148( .ZN(N3371), .A1(N3327), .A2(N3328) );
  NOR2_X1 NOR2_1149( .ZN(N3374), .A1(N3329), .A2(N3330) );
  NOR2_X1 NOR2_1150( .ZN(N3377), .A1(N3331), .A2(N3332) );
  NOR2_X1 NOR2_1151( .ZN(N3380), .A1(N3333), .A2(N3334) );
  NOR2_X1 NOR2_1152( .ZN(N3383), .A1(N3335), .A2(N3336) );
  NOR2_X1 NOR2_1153( .ZN(N3386), .A1(N3337), .A2(N3338) );
  NOR2_X1 NOR2_1154( .ZN(N3389), .A1(N3339), .A2(N3340) );
  NOR2_X1 NOR2_1155( .ZN(N3392), .A1(N3341), .A2(N996) );
  NOR2_X1 NOR2_1156( .ZN(N3396), .A1(N3302), .A2(N3344) );
  NOR2_X2 NOR2_1157( .ZN(N3397), .A1(N3344), .A2(N1044) );
  NOR2_X2 NOR2_1158( .ZN(N3398), .A1(N3193), .A2(N3344) );
  NOR2_X2 NOR2_1159( .ZN(N3401), .A1(N3348), .A2(N3349) );
  NOR2_X2 NOR2_1160( .ZN(N3404), .A1(N3353), .A2(N3350) );
  NOR2_X1 NOR2_1161( .ZN(N3408), .A1(N3314), .A2(N3356) );
  NOR2_X1 NOR2_1162( .ZN(N3409), .A1(N3356), .A2(N3311) );
  NOR2_X1 NOR2_1163( .ZN(N3410), .A1(N3360), .A2(N3361) );
  NOR2_X1 NOR2_1164( .ZN(N3413), .A1(N3362), .A2(N1239) );
  NOR2_X1 NOR2_1165( .ZN(N3417), .A1(N3365), .A2(N564) );
  NOR2_X1 NOR2_1166( .ZN(N3421), .A1(N3368), .A2(N612) );
  NOR2_X1 NOR2_1167( .ZN(N3425), .A1(N3371), .A2(N660) );
  NOR2_X1 NOR2_1168( .ZN(N3429), .A1(N3374), .A2(N708) );
  NOR2_X1 NOR2_1169( .ZN(N3433), .A1(N3377), .A2(N756) );
  NOR2_X1 NOR2_1170( .ZN(N3437), .A1(N3380), .A2(N804) );
  NOR2_X1 NOR2_1171( .ZN(N3441), .A1(N3383), .A2(N852) );
  NOR2_X1 NOR2_1172( .ZN(N3445), .A1(N3386), .A2(N900) );
  NOR2_X1 NOR2_1173( .ZN(N3449), .A1(N3389), .A2(N948) );
  NOR2_X1 NOR2_1174( .ZN(N3453), .A1(N3341), .A2(N3392) );
  NOR2_X1 NOR2_1175( .ZN(N3454), .A1(N3392), .A2(N996) );
  NOR2_X1 NOR2_1176( .ZN(N3455), .A1(N3239), .A2(N3392) );
  NOR2_X1 NOR2_1177( .ZN(N3458), .A1(N3396), .A2(N3397) );
  NOR2_X1 NOR2_1178( .ZN(N3461), .A1(N3401), .A2(N3398) );
  NOR2_X1 NOR2_1179( .ZN(N3465), .A1(N3353), .A2(N3404) );
  NOR2_X1 NOR2_1180( .ZN(N3466), .A1(N3404), .A2(N3350) );
  NOR2_X1 NOR2_1181( .ZN(N3467), .A1(N3408), .A2(N3409) );
  NOR2_X1 NOR2_1182( .ZN(N3470), .A1(N3410), .A2(N1191) );
  NOR2_X1 NOR2_1183( .ZN(N3474), .A1(N3362), .A2(N3413) );
  NOR2_X1 NOR2_1184( .ZN(N3475), .A1(N3413), .A2(N1239) );
  NOR2_X1 NOR2_1185( .ZN(N3476), .A1(N3260), .A2(N3413) );
  NOR2_X1 NOR2_1186( .ZN(N3479), .A1(N3365), .A2(N3417) );
  NOR2_X1 NOR2_1187( .ZN(N3480), .A1(N3417), .A2(N564) );
  NOR2_X1 NOR2_1188( .ZN(N3481), .A1(N3264), .A2(N3417) );
  NOR2_X1 NOR2_1189( .ZN(N3484), .A1(N3368), .A2(N3421) );
  NOR2_X1 NOR2_1190( .ZN(N3485), .A1(N3421), .A2(N612) );
  NOR2_X1 NOR2_1191( .ZN(N3486), .A1(N3268), .A2(N3421) );
  NOR2_X1 NOR2_1192( .ZN(N3489), .A1(N3371), .A2(N3425) );
  NOR2_X1 NOR2_1193( .ZN(N3490), .A1(N3425), .A2(N660) );
  NOR2_X1 NOR2_1194( .ZN(N3491), .A1(N3272), .A2(N3425) );
  NOR2_X1 NOR2_1195( .ZN(N3494), .A1(N3374), .A2(N3429) );
  NOR2_X1 NOR2_1196( .ZN(N3495), .A1(N3429), .A2(N708) );
  NOR2_X1 NOR2_1197( .ZN(N3496), .A1(N3276), .A2(N3429) );
  NOR2_X1 NOR2_1198( .ZN(N3499), .A1(N3377), .A2(N3433) );
  NOR2_X1 NOR2_1199( .ZN(N3500), .A1(N3433), .A2(N756) );
  NOR2_X1 NOR2_1200( .ZN(N3501), .A1(N3280), .A2(N3433) );
  NOR2_X1 NOR2_1201( .ZN(N3504), .A1(N3380), .A2(N3437) );
  NOR2_X1 NOR2_1202( .ZN(N3505), .A1(N3437), .A2(N804) );
  NOR2_X1 NOR2_1203( .ZN(N3506), .A1(N3284), .A2(N3437) );
  NOR2_X1 NOR2_1204( .ZN(N3509), .A1(N3383), .A2(N3441) );
  NOR2_X1 NOR2_1205( .ZN(N3510), .A1(N3441), .A2(N852) );
  NOR2_X1 NOR2_1206( .ZN(N3511), .A1(N3288), .A2(N3441) );
  NOR2_X1 NOR2_1207( .ZN(N3514), .A1(N3386), .A2(N3445) );
  NOR2_X1 NOR2_1208( .ZN(N3515), .A1(N3445), .A2(N900) );
  NOR2_X1 NOR2_1209( .ZN(N3516), .A1(N3292), .A2(N3445) );
  NOR2_X1 NOR2_1210( .ZN(N3519), .A1(N3389), .A2(N3449) );
  NOR2_X1 NOR2_1211( .ZN(N3520), .A1(N3449), .A2(N948) );
  NOR2_X1 NOR2_1212( .ZN(N3521), .A1(N3296), .A2(N3449) );
  NOR2_X1 NOR2_1213( .ZN(N3524), .A1(N3453), .A2(N3454) );
  NOR2_X1 NOR2_1214( .ZN(N3527), .A1(N3458), .A2(N3455) );
  NOR2_X1 NOR2_1215( .ZN(N3531), .A1(N3401), .A2(N3461) );
  NOR2_X1 NOR2_1216( .ZN(N3532), .A1(N3461), .A2(N3398) );
  NOR2_X1 NOR2_1217( .ZN(N3533), .A1(N3465), .A2(N3466) );
  NOR2_X1 NOR2_1218( .ZN(N3536), .A1(N3467), .A2(N1143) );
  NOR2_X1 NOR2_1219( .ZN(N3540), .A1(N3410), .A2(N3470) );
  NOR2_X1 NOR2_1220( .ZN(N3541), .A1(N3470), .A2(N1191) );
  NOR2_X1 NOR2_1221( .ZN(N3542), .A1(N3317), .A2(N3470) );
  NOR2_X1 NOR2_1222( .ZN(N3545), .A1(N3474), .A2(N3475) );
  NOR2_X1 NOR2_1223( .ZN(N3548), .A1(N1287), .A2(N3476) );
  NOR2_X1 NOR2_1224( .ZN(N3552), .A1(N3479), .A2(N3480) );
  NOR2_X1 NOR2_1225( .ZN(N3553), .A1(N3484), .A2(N3485) );
  NOR2_X1 NOR2_1226( .ZN(N3556), .A1(N3489), .A2(N3490) );
  NOR2_X1 NOR2_1227( .ZN(N3559), .A1(N3494), .A2(N3495) );
  NOR2_X1 NOR2_1228( .ZN(N3562), .A1(N3499), .A2(N3500) );
  NOR2_X1 NOR2_1229( .ZN(N3565), .A1(N3504), .A2(N3505) );
  NOR2_X1 NOR2_1230( .ZN(N3568), .A1(N3509), .A2(N3510) );
  NOR2_X1 NOR2_1231( .ZN(N3571), .A1(N3514), .A2(N3515) );
  NOR2_X1 NOR2_1232( .ZN(N3574), .A1(N3519), .A2(N3520) );
  NOR2_X1 NOR2_1233( .ZN(N3577), .A1(N3524), .A2(N3521) );
  NOR2_X1 NOR2_1234( .ZN(N3581), .A1(N3458), .A2(N3527) );
  NOR2_X1 NOR2_1235( .ZN(N3582), .A1(N3527), .A2(N3455) );
  NOR2_X1 NOR2_1236( .ZN(N3583), .A1(N3531), .A2(N3532) );
  NOR2_X1 NOR2_1237( .ZN(N3586), .A1(N3533), .A2(N1095) );
  NOR2_X1 NOR2_1238( .ZN(N3590), .A1(N3467), .A2(N3536) );
  NOR2_X1 NOR2_1239( .ZN(N3591), .A1(N3536), .A2(N1143) );
  NOR2_X1 NOR2_1240( .ZN(N3592), .A1(N3356), .A2(N3536) );
  NOR2_X1 NOR2_1241( .ZN(N3595), .A1(N3540), .A2(N3541) );
  NOR2_X1 NOR2_1242( .ZN(N3598), .A1(N3545), .A2(N3542) );
  NOR2_X1 NOR2_1243( .ZN(N3602), .A1(N1287), .A2(N3548) );
  NOR2_X1 NOR2_1244( .ZN(N3603), .A1(N3548), .A2(N3476) );
  NOR2_X1 NOR2_1245( .ZN(N3604), .A1(N3553), .A2(N3481) );
  NOR2_X1 NOR2_1246( .ZN(N3608), .A1(N3556), .A2(N3486) );
  NOR2_X1 NOR2_1247( .ZN(N3612), .A1(N3559), .A2(N3491) );
  NOR2_X1 NOR2_1248( .ZN(N3616), .A1(N3562), .A2(N3496) );
  NOR2_X1 NOR2_1249( .ZN(N3620), .A1(N3565), .A2(N3501) );
  NOR2_X1 NOR2_1250( .ZN(N3624), .A1(N3568), .A2(N3506) );
  NOR2_X1 NOR2_1251( .ZN(N3628), .A1(N3571), .A2(N3511) );
  NOR2_X1 NOR2_1252( .ZN(N3632), .A1(N3574), .A2(N3516) );
  NOR2_X1 NOR2_1253( .ZN(N3636), .A1(N3524), .A2(N3577) );
  NOR2_X1 NOR2_1254( .ZN(N3637), .A1(N3577), .A2(N3521) );
  NOR2_X1 NOR2_1255( .ZN(N3638), .A1(N3581), .A2(N3582) );
  NOR2_X1 NOR2_1256( .ZN(N3641), .A1(N3583), .A2(N1047) );
  NOR2_X1 NOR2_1257( .ZN(N3645), .A1(N3533), .A2(N3586) );
  NOR2_X1 NOR2_1258( .ZN(N3646), .A1(N3586), .A2(N1095) );
  NOR2_X1 NOR2_1259( .ZN(N3647), .A1(N3404), .A2(N3586) );
  NOR2_X1 NOR2_1260( .ZN(N3650), .A1(N3590), .A2(N3591) );
  NOR2_X1 NOR2_1261( .ZN(N3653), .A1(N3595), .A2(N3592) );
  NOR2_X1 NOR2_1262( .ZN(N3657), .A1(N3545), .A2(N3598) );
  NOR2_X1 NOR2_1263( .ZN(N3658), .A1(N3598), .A2(N3542) );
  NOR2_X1 NOR2_1264( .ZN(N3659), .A1(N3602), .A2(N3603) );
  NOR2_X1 NOR2_1265( .ZN(N3662), .A1(N3553), .A2(N3604) );
  NOR2_X1 NOR2_1266( .ZN(N3663), .A1(N3604), .A2(N3481) );
  NOR2_X1 NOR2_1267( .ZN(N3664), .A1(N3556), .A2(N3608) );
  NOR2_X1 NOR2_1268( .ZN(N3665), .A1(N3608), .A2(N3486) );
  NOR2_X1 NOR2_1269( .ZN(N3666), .A1(N3559), .A2(N3612) );
  NOR2_X1 NOR2_1270( .ZN(N3667), .A1(N3612), .A2(N3491) );
  NOR2_X1 NOR2_1271( .ZN(N3668), .A1(N3562), .A2(N3616) );
  NOR2_X1 NOR2_1272( .ZN(N3669), .A1(N3616), .A2(N3496) );
  NOR2_X1 NOR2_1273( .ZN(N3670), .A1(N3565), .A2(N3620) );
  NOR2_X1 NOR2_1274( .ZN(N3671), .A1(N3620), .A2(N3501) );
  NOR2_X1 NOR2_1275( .ZN(N3672), .A1(N3568), .A2(N3624) );
  NOR2_X1 NOR2_1276( .ZN(N3673), .A1(N3624), .A2(N3506) );
  NOR2_X1 NOR2_1277( .ZN(N3674), .A1(N3571), .A2(N3628) );
  NOR2_X1 NOR2_1278( .ZN(N3675), .A1(N3628), .A2(N3511) );
  NOR2_X1 NOR2_1279( .ZN(N3676), .A1(N3574), .A2(N3632) );
  NOR2_X1 NOR2_1280( .ZN(N3677), .A1(N3632), .A2(N3516) );
  NOR2_X1 NOR2_1281( .ZN(N3678), .A1(N3636), .A2(N3637) );
  NOR2_X1 NOR2_1282( .ZN(N3681), .A1(N3638), .A2(N999) );
  NOR2_X1 NOR2_1283( .ZN(N3685), .A1(N3583), .A2(N3641) );
  NOR2_X1 NOR2_1284( .ZN(N3686), .A1(N3641), .A2(N1047) );
  NOR2_X1 NOR2_1285( .ZN(N3687), .A1(N3461), .A2(N3641) );
  NOR2_X1 NOR2_1286( .ZN(N3690), .A1(N3645), .A2(N3646) );
  NOR2_X1 NOR2_1287( .ZN(N3693), .A1(N3650), .A2(N3647) );
  NOR2_X1 NOR2_1288( .ZN(N3697), .A1(N3595), .A2(N3653) );
  NOR2_X1 NOR2_1289( .ZN(N3698), .A1(N3653), .A2(N3592) );
  NOR2_X1 NOR2_1290( .ZN(N3699), .A1(N3657), .A2(N3658) );
  NOR2_X1 NOR2_1291( .ZN(N3702), .A1(N3659), .A2(N1242) );
  NOR2_X1 NOR2_1292( .ZN(N3706), .A1(N3662), .A2(N3663) );
  NOR2_X1 NOR2_1293( .ZN(N3709), .A1(N3664), .A2(N3665) );
  NOR2_X1 NOR2_1294( .ZN(N3712), .A1(N3666), .A2(N3667) );
  NOR2_X1 NOR2_1295( .ZN(N3715), .A1(N3668), .A2(N3669) );
  NOR2_X1 NOR2_1296( .ZN(N3718), .A1(N3670), .A2(N3671) );
  NOR2_X1 NOR2_1297( .ZN(N3721), .A1(N3672), .A2(N3673) );
  NOR2_X1 NOR2_1298( .ZN(N3724), .A1(N3674), .A2(N3675) );
  NOR2_X1 NOR2_1299( .ZN(N3727), .A1(N3676), .A2(N3677) );
  NOR2_X1 NOR2_1300( .ZN(N3730), .A1(N3678), .A2(N951) );
  NOR2_X1 NOR2_1301( .ZN(N3734), .A1(N3638), .A2(N3681) );
  NOR2_X1 NOR2_1302( .ZN(N3735), .A1(N3681), .A2(N999) );
  NOR2_X1 NOR2_1303( .ZN(N3736), .A1(N3527), .A2(N3681) );
  NOR2_X1 NOR2_1304( .ZN(N3739), .A1(N3685), .A2(N3686) );
  NOR2_X1 NOR2_1305( .ZN(N3742), .A1(N3690), .A2(N3687) );
  NOR2_X1 NOR2_1306( .ZN(N3746), .A1(N3650), .A2(N3693) );
  NOR2_X1 NOR2_1307( .ZN(N3747), .A1(N3693), .A2(N3647) );
  NOR2_X1 NOR2_1308( .ZN(N3748), .A1(N3697), .A2(N3698) );
  NOR2_X1 NOR2_1309( .ZN(N3751), .A1(N3699), .A2(N1194) );
  NOR2_X1 NOR2_1310( .ZN(N3755), .A1(N3659), .A2(N3702) );
  NOR2_X1 NOR2_1311( .ZN(N3756), .A1(N3702), .A2(N1242) );
  NOR2_X1 NOR2_1312( .ZN(N3757), .A1(N3548), .A2(N3702) );
  NOR2_X1 NOR2_1313( .ZN(N3760), .A1(N3706), .A2(N567) );
  NOR2_X1 NOR2_1314( .ZN(N3764), .A1(N3709), .A2(N615) );
  NOR2_X1 NOR2_1315( .ZN(N3768), .A1(N3712), .A2(N663) );
  NOR2_X1 NOR2_1316( .ZN(N3772), .A1(N3715), .A2(N711) );
  NOR2_X1 NOR2_1317( .ZN(N3776), .A1(N3718), .A2(N759) );
  NOR2_X1 NOR2_1318( .ZN(N3780), .A1(N3721), .A2(N807) );
  NOR2_X1 NOR2_1319( .ZN(N3784), .A1(N3724), .A2(N855) );
  NOR2_X1 NOR2_1320( .ZN(N3788), .A1(N3727), .A2(N903) );
  NOR2_X1 NOR2_1321( .ZN(N3792), .A1(N3678), .A2(N3730) );
  NOR2_X1 NOR2_1322( .ZN(N3793), .A1(N3730), .A2(N951) );
  NOR2_X1 NOR2_1323( .ZN(N3794), .A1(N3577), .A2(N3730) );
  NOR2_X1 NOR2_1324( .ZN(N3797), .A1(N3734), .A2(N3735) );
  NOR2_X1 NOR2_1325( .ZN(N3800), .A1(N3739), .A2(N3736) );
  NOR2_X1 NOR2_1326( .ZN(N3804), .A1(N3690), .A2(N3742) );
  NOR2_X1 NOR2_1327( .ZN(N3805), .A1(N3742), .A2(N3687) );
  NOR2_X1 NOR2_1328( .ZN(N3806), .A1(N3746), .A2(N3747) );
  NOR2_X1 NOR2_1329( .ZN(N3809), .A1(N3748), .A2(N1146) );
  NOR2_X1 NOR2_1330( .ZN(N3813), .A1(N3699), .A2(N3751) );
  NOR2_X1 NOR2_1331( .ZN(N3814), .A1(N3751), .A2(N1194) );
  NOR2_X1 NOR2_1332( .ZN(N3815), .A1(N3598), .A2(N3751) );
  NOR2_X1 NOR2_1333( .ZN(N3818), .A1(N3755), .A2(N3756) );
  NOR2_X1 NOR2_1334( .ZN(N3821), .A1(N1290), .A2(N3757) );
  NOR2_X1 NOR2_1335( .ZN(N3825), .A1(N3706), .A2(N3760) );
  NOR2_X1 NOR2_1336( .ZN(N3826), .A1(N3760), .A2(N567) );
  NOR2_X1 NOR2_1337( .ZN(N3827), .A1(N3604), .A2(N3760) );
  NOR2_X1 NOR2_1338( .ZN(N3830), .A1(N3709), .A2(N3764) );
  NOR2_X1 NOR2_1339( .ZN(N3831), .A1(N3764), .A2(N615) );
  NOR2_X1 NOR2_1340( .ZN(N3832), .A1(N3608), .A2(N3764) );
  NOR2_X1 NOR2_1341( .ZN(N3835), .A1(N3712), .A2(N3768) );
  NOR2_X1 NOR2_1342( .ZN(N3836), .A1(N3768), .A2(N663) );
  NOR2_X1 NOR2_1343( .ZN(N3837), .A1(N3612), .A2(N3768) );
  NOR2_X1 NOR2_1344( .ZN(N3840), .A1(N3715), .A2(N3772) );
  NOR2_X1 NOR2_1345( .ZN(N3841), .A1(N3772), .A2(N711) );
  NOR2_X1 NOR2_1346( .ZN(N3842), .A1(N3616), .A2(N3772) );
  NOR2_X1 NOR2_1347( .ZN(N3845), .A1(N3718), .A2(N3776) );
  NOR2_X1 NOR2_1348( .ZN(N3846), .A1(N3776), .A2(N759) );
  NOR2_X1 NOR2_1349( .ZN(N3847), .A1(N3620), .A2(N3776) );
  NOR2_X1 NOR2_1350( .ZN(N3850), .A1(N3721), .A2(N3780) );
  NOR2_X1 NOR2_1351( .ZN(N3851), .A1(N3780), .A2(N807) );
  NOR2_X1 NOR2_1352( .ZN(N3852), .A1(N3624), .A2(N3780) );
  NOR2_X1 NOR2_1353( .ZN(N3855), .A1(N3724), .A2(N3784) );
  NOR2_X1 NOR2_1354( .ZN(N3856), .A1(N3784), .A2(N855) );
  NOR2_X1 NOR2_1355( .ZN(N3857), .A1(N3628), .A2(N3784) );
  NOR2_X1 NOR2_1356( .ZN(N3860), .A1(N3727), .A2(N3788) );
  NOR2_X1 NOR2_1357( .ZN(N3861), .A1(N3788), .A2(N903) );
  NOR2_X1 NOR2_1358( .ZN(N3862), .A1(N3632), .A2(N3788) );
  NOR2_X1 NOR2_1359( .ZN(N3865), .A1(N3792), .A2(N3793) );
  NOR2_X1 NOR2_1360( .ZN(N3868), .A1(N3797), .A2(N3794) );
  NOR2_X1 NOR2_1361( .ZN(N3872), .A1(N3739), .A2(N3800) );
  NOR2_X1 NOR2_1362( .ZN(N3873), .A1(N3800), .A2(N3736) );
  NOR2_X1 NOR2_1363( .ZN(N3874), .A1(N3804), .A2(N3805) );
  NOR2_X1 NOR2_1364( .ZN(N3877), .A1(N3806), .A2(N1098) );
  NOR2_X1 NOR2_1365( .ZN(N3881), .A1(N3748), .A2(N3809) );
  NOR2_X1 NOR2_1366( .ZN(N3882), .A1(N3809), .A2(N1146) );
  NOR2_X1 NOR2_1367( .ZN(N3883), .A1(N3653), .A2(N3809) );
  NOR2_X1 NOR2_1368( .ZN(N3886), .A1(N3813), .A2(N3814) );
  NOR2_X1 NOR2_1369( .ZN(N3889), .A1(N3818), .A2(N3815) );
  NOR2_X1 NOR2_1370( .ZN(N3893), .A1(N1290), .A2(N3821) );
  NOR2_X1 NOR2_1371( .ZN(N3894), .A1(N3821), .A2(N3757) );
  NOR2_X1 NOR2_1372( .ZN(N3895), .A1(N3825), .A2(N3826) );
  NOR2_X1 NOR2_1373( .ZN(N3896), .A1(N3830), .A2(N3831) );
  NOR2_X1 NOR2_1374( .ZN(N3899), .A1(N3835), .A2(N3836) );
  NOR2_X1 NOR2_1375( .ZN(N3902), .A1(N3840), .A2(N3841) );
  NOR2_X1 NOR2_1376( .ZN(N3905), .A1(N3845), .A2(N3846) );
  NOR2_X1 NOR2_1377( .ZN(N3908), .A1(N3850), .A2(N3851) );
  NOR2_X1 NOR2_1378( .ZN(N3911), .A1(N3855), .A2(N3856) );
  NOR2_X1 NOR2_1379( .ZN(N3914), .A1(N3860), .A2(N3861) );
  NOR2_X1 NOR2_1380( .ZN(N3917), .A1(N3865), .A2(N3862) );
  NOR2_X1 NOR2_1381( .ZN(N3921), .A1(N3797), .A2(N3868) );
  NOR2_X1 NOR2_1382( .ZN(N3922), .A1(N3868), .A2(N3794) );
  NOR2_X1 NOR2_1383( .ZN(N3923), .A1(N3872), .A2(N3873) );
  NOR2_X1 NOR2_1384( .ZN(N3926), .A1(N3874), .A2(N1050) );
  NOR2_X1 NOR2_1385( .ZN(N3930), .A1(N3806), .A2(N3877) );
  NOR2_X1 NOR2_1386( .ZN(N3931), .A1(N3877), .A2(N1098) );
  NOR2_X1 NOR2_1387( .ZN(N3932), .A1(N3693), .A2(N3877) );
  NOR2_X1 NOR2_1388( .ZN(N3935), .A1(N3881), .A2(N3882) );
  NOR2_X1 NOR2_1389( .ZN(N3938), .A1(N3886), .A2(N3883) );
  NOR2_X1 NOR2_1390( .ZN(N3942), .A1(N3818), .A2(N3889) );
  NOR2_X1 NOR2_1391( .ZN(N3943), .A1(N3889), .A2(N3815) );
  NOR2_X1 NOR2_1392( .ZN(N3944), .A1(N3893), .A2(N3894) );
  NOR2_X1 NOR2_1393( .ZN(N3947), .A1(N3896), .A2(N3827) );
  NOR2_X1 NOR2_1394( .ZN(N3951), .A1(N3899), .A2(N3832) );
  NOR2_X1 NOR2_1395( .ZN(N3955), .A1(N3902), .A2(N3837) );
  NOR2_X1 NOR2_1396( .ZN(N3959), .A1(N3905), .A2(N3842) );
  NOR2_X1 NOR2_1397( .ZN(N3963), .A1(N3908), .A2(N3847) );
  NOR2_X1 NOR2_1398( .ZN(N3967), .A1(N3911), .A2(N3852) );
  NOR2_X1 NOR2_1399( .ZN(N3971), .A1(N3914), .A2(N3857) );
  NOR2_X1 NOR2_1400( .ZN(N3975), .A1(N3865), .A2(N3917) );
  NOR2_X1 NOR2_1401( .ZN(N3976), .A1(N3917), .A2(N3862) );
  NOR2_X1 NOR2_1402( .ZN(N3977), .A1(N3921), .A2(N3922) );
  NOR2_X1 NOR2_1403( .ZN(N3980), .A1(N3923), .A2(N1002) );
  NOR2_X1 NOR2_1404( .ZN(N3984), .A1(N3874), .A2(N3926) );
  NOR2_X1 NOR2_1405( .ZN(N3985), .A1(N3926), .A2(N1050) );
  NOR2_X1 NOR2_1406( .ZN(N3986), .A1(N3742), .A2(N3926) );
  NOR2_X1 NOR2_1407( .ZN(N3989), .A1(N3930), .A2(N3931) );
  NOR2_X1 NOR2_1408( .ZN(N3992), .A1(N3935), .A2(N3932) );
  NOR2_X1 NOR2_1409( .ZN(N3996), .A1(N3886), .A2(N3938) );
  NOR2_X1 NOR2_1410( .ZN(N3997), .A1(N3938), .A2(N3883) );
  NOR2_X1 NOR2_1411( .ZN(N3998), .A1(N3942), .A2(N3943) );
  NOR2_X1 NOR2_1412( .ZN(N4001), .A1(N3944), .A2(N1245) );
  NOR2_X1 NOR2_1413( .ZN(N4005), .A1(N3896), .A2(N3947) );
  NOR2_X1 NOR2_1414( .ZN(N4006), .A1(N3947), .A2(N3827) );
  NOR2_X1 NOR2_1415( .ZN(N4007), .A1(N3899), .A2(N3951) );
  NOR2_X1 NOR2_1416( .ZN(N4008), .A1(N3951), .A2(N3832) );
  NOR2_X1 NOR2_1417( .ZN(N4009), .A1(N3902), .A2(N3955) );
  NOR2_X1 NOR2_1418( .ZN(N4010), .A1(N3955), .A2(N3837) );
  NOR2_X1 NOR2_1419( .ZN(N4011), .A1(N3905), .A2(N3959) );
  NOR2_X1 NOR2_1420( .ZN(N4012), .A1(N3959), .A2(N3842) );
  NOR2_X1 NOR2_1421( .ZN(N4013), .A1(N3908), .A2(N3963) );
  NOR2_X1 NOR2_1422( .ZN(N4014), .A1(N3963), .A2(N3847) );
  NOR2_X1 NOR2_1423( .ZN(N4015), .A1(N3911), .A2(N3967) );
  NOR2_X1 NOR2_1424( .ZN(N4016), .A1(N3967), .A2(N3852) );
  NOR2_X1 NOR2_1425( .ZN(N4017), .A1(N3914), .A2(N3971) );
  NOR2_X1 NOR2_1426( .ZN(N4018), .A1(N3971), .A2(N3857) );
  NOR2_X1 NOR2_1427( .ZN(N4019), .A1(N3975), .A2(N3976) );
  NOR2_X1 NOR2_1428( .ZN(N4022), .A1(N3977), .A2(N954) );
  NOR2_X1 NOR2_1429( .ZN(N4026), .A1(N3923), .A2(N3980) );
  NOR2_X1 NOR2_1430( .ZN(N4027), .A1(N3980), .A2(N1002) );
  NOR2_X1 NOR2_1431( .ZN(N4028), .A1(N3800), .A2(N3980) );
  NOR2_X1 NOR2_1432( .ZN(N4031), .A1(N3984), .A2(N3985) );
  NOR2_X1 NOR2_1433( .ZN(N4034), .A1(N3989), .A2(N3986) );
  NOR2_X1 NOR2_1434( .ZN(N4038), .A1(N3935), .A2(N3992) );
  NOR2_X1 NOR2_1435( .ZN(N4039), .A1(N3992), .A2(N3932) );
  NOR2_X1 NOR2_1436( .ZN(N4040), .A1(N3996), .A2(N3997) );
  NOR2_X1 NOR2_1437( .ZN(N4043), .A1(N3998), .A2(N1197) );
  NOR2_X1 NOR2_1438( .ZN(N4047), .A1(N3944), .A2(N4001) );
  NOR2_X1 NOR2_1439( .ZN(N4048), .A1(N4001), .A2(N1245) );
  NOR2_X1 NOR2_1440( .ZN(N4049), .A1(N3821), .A2(N4001) );
  NOR2_X1 NOR2_1441( .ZN(N4052), .A1(N4005), .A2(N4006) );
  NOR2_X1 NOR2_1442( .ZN(N4055), .A1(N4007), .A2(N4008) );
  NOR2_X1 NOR2_1443( .ZN(N4058), .A1(N4009), .A2(N4010) );
  NOR2_X1 NOR2_1444( .ZN(N4061), .A1(N4011), .A2(N4012) );
  NOR2_X1 NOR2_1445( .ZN(N4064), .A1(N4013), .A2(N4014) );
  NOR2_X1 NOR2_1446( .ZN(N4067), .A1(N4015), .A2(N4016) );
  NOR2_X1 NOR2_1447( .ZN(N4070), .A1(N4017), .A2(N4018) );
  NOR2_X1 NOR2_1448( .ZN(N4073), .A1(N4019), .A2(N906) );
  NOR2_X1 NOR2_1449( .ZN(N4077), .A1(N3977), .A2(N4022) );
  NOR2_X1 NOR2_1450( .ZN(N4078), .A1(N4022), .A2(N954) );
  NOR2_X1 NOR2_1451( .ZN(N4079), .A1(N3868), .A2(N4022) );
  NOR2_X1 NOR2_1452( .ZN(N4082), .A1(N4026), .A2(N4027) );
  NOR2_X1 NOR2_1453( .ZN(N4085), .A1(N4031), .A2(N4028) );
  NOR2_X1 NOR2_1454( .ZN(N4089), .A1(N3989), .A2(N4034) );
  NOR2_X1 NOR2_1455( .ZN(N4090), .A1(N4034), .A2(N3986) );
  NOR2_X1 NOR2_1456( .ZN(N4091), .A1(N4038), .A2(N4039) );
  NOR2_X1 NOR2_1457( .ZN(N4094), .A1(N4040), .A2(N1149) );
  NOR2_X1 NOR2_1458( .ZN(N4098), .A1(N3998), .A2(N4043) );
  NOR2_X1 NOR2_1459( .ZN(N4099), .A1(N4043), .A2(N1197) );
  NOR2_X1 NOR2_1460( .ZN(N4100), .A1(N3889), .A2(N4043) );
  NOR2_X1 NOR2_1461( .ZN(N4103), .A1(N4047), .A2(N4048) );
  NOR2_X1 NOR2_1462( .ZN(N4106), .A1(N1293), .A2(N4049) );
  NOR2_X1 NOR2_1463( .ZN(N4110), .A1(N4052), .A2(N570) );
  NOR2_X1 NOR2_1464( .ZN(N4114), .A1(N4055), .A2(N618) );
  NOR2_X1 NOR2_1465( .ZN(N4118), .A1(N4058), .A2(N666) );
  NOR2_X1 NOR2_1466( .ZN(N4122), .A1(N4061), .A2(N714) );
  NOR2_X1 NOR2_1467( .ZN(N4126), .A1(N4064), .A2(N762) );
  NOR2_X1 NOR2_1468( .ZN(N4130), .A1(N4067), .A2(N810) );
  NOR2_X1 NOR2_1469( .ZN(N4134), .A1(N4070), .A2(N858) );
  NOR2_X1 NOR2_1470( .ZN(N4138), .A1(N4019), .A2(N4073) );
  NOR2_X1 NOR2_1471( .ZN(N4139), .A1(N4073), .A2(N906) );
  NOR2_X1 NOR2_1472( .ZN(N4140), .A1(N3917), .A2(N4073) );
  NOR2_X2 NOR2_1473( .ZN(N4143), .A1(N4077), .A2(N4078) );
  NOR2_X2 NOR2_1474( .ZN(N4146), .A1(N4082), .A2(N4079) );
  NOR2_X2 NOR2_1475( .ZN(N4150), .A1(N4031), .A2(N4085) );
  NOR2_X2 NOR2_1476( .ZN(N4151), .A1(N4085), .A2(N4028) );
  NOR2_X2 NOR2_1477( .ZN(N4152), .A1(N4089), .A2(N4090) );
  NOR2_X2 NOR2_1478( .ZN(N4155), .A1(N4091), .A2(N1101) );
  NOR2_X2 NOR2_1479( .ZN(N4159), .A1(N4040), .A2(N4094) );
  NOR2_X2 NOR2_1480( .ZN(N4160), .A1(N4094), .A2(N1149) );
  NOR2_X1 NOR2_1481( .ZN(N4161), .A1(N3938), .A2(N4094) );
  NOR2_X1 NOR2_1482( .ZN(N4164), .A1(N4098), .A2(N4099) );
  NOR2_X1 NOR2_1483( .ZN(N4167), .A1(N4103), .A2(N4100) );
  NOR2_X1 NOR2_1484( .ZN(N4171), .A1(N1293), .A2(N4106) );
  NOR2_X1 NOR2_1485( .ZN(N4172), .A1(N4106), .A2(N4049) );
  NOR2_X1 NOR2_1486( .ZN(N4173), .A1(N4052), .A2(N4110) );
  NOR2_X1 NOR2_1487( .ZN(N4174), .A1(N4110), .A2(N570) );
  NOR2_X1 NOR2_1488( .ZN(N4175), .A1(N3947), .A2(N4110) );
  NOR2_X1 NOR2_1489( .ZN(N4178), .A1(N4055), .A2(N4114) );
  NOR2_X1 NOR2_1490( .ZN(N4179), .A1(N4114), .A2(N618) );
  NOR2_X1 NOR2_1491( .ZN(N4180), .A1(N3951), .A2(N4114) );
  NOR2_X1 NOR2_1492( .ZN(N4183), .A1(N4058), .A2(N4118) );
  NOR2_X1 NOR2_1493( .ZN(N4184), .A1(N4118), .A2(N666) );
  NOR2_X1 NOR2_1494( .ZN(N4185), .A1(N3955), .A2(N4118) );
  NOR2_X1 NOR2_1495( .ZN(N4188), .A1(N4061), .A2(N4122) );
  NOR2_X1 NOR2_1496( .ZN(N4189), .A1(N4122), .A2(N714) );
  NOR2_X1 NOR2_1497( .ZN(N4190), .A1(N3959), .A2(N4122) );
  NOR2_X1 NOR2_1498( .ZN(N4193), .A1(N4064), .A2(N4126) );
  NOR2_X1 NOR2_1499( .ZN(N4194), .A1(N4126), .A2(N762) );
  NOR2_X1 NOR2_1500( .ZN(N4195), .A1(N3963), .A2(N4126) );
  NOR2_X1 NOR2_1501( .ZN(N4198), .A1(N4067), .A2(N4130) );
  NOR2_X1 NOR2_1502( .ZN(N4199), .A1(N4130), .A2(N810) );
  NOR2_X1 NOR2_1503( .ZN(N4200), .A1(N3967), .A2(N4130) );
  NOR2_X1 NOR2_1504( .ZN(N4203), .A1(N4070), .A2(N4134) );
  NOR2_X1 NOR2_1505( .ZN(N4204), .A1(N4134), .A2(N858) );
  NOR2_X1 NOR2_1506( .ZN(N4205), .A1(N3971), .A2(N4134) );
  NOR2_X1 NOR2_1507( .ZN(N4208), .A1(N4138), .A2(N4139) );
  NOR2_X1 NOR2_1508( .ZN(N4211), .A1(N4143), .A2(N4140) );
  NOR2_X1 NOR2_1509( .ZN(N4215), .A1(N4082), .A2(N4146) );
  NOR2_X1 NOR2_1510( .ZN(N4216), .A1(N4146), .A2(N4079) );
  NOR2_X1 NOR2_1511( .ZN(N4217), .A1(N4150), .A2(N4151) );
  NOR2_X1 NOR2_1512( .ZN(N4220), .A1(N4152), .A2(N1053) );
  NOR2_X1 NOR2_1513( .ZN(N4224), .A1(N4091), .A2(N4155) );
  NOR2_X1 NOR2_1514( .ZN(N4225), .A1(N4155), .A2(N1101) );
  NOR2_X1 NOR2_1515( .ZN(N4226), .A1(N3992), .A2(N4155) );
  NOR2_X1 NOR2_1516( .ZN(N4229), .A1(N4159), .A2(N4160) );
  NOR2_X1 NOR2_1517( .ZN(N4232), .A1(N4164), .A2(N4161) );
  NOR2_X1 NOR2_1518( .ZN(N4236), .A1(N4103), .A2(N4167) );
  NOR2_X1 NOR2_1519( .ZN(N4237), .A1(N4167), .A2(N4100) );
  NOR2_X1 NOR2_1520( .ZN(N4238), .A1(N4171), .A2(N4172) );
  NOR2_X1 NOR2_1521( .ZN(N4241), .A1(N4173), .A2(N4174) );
  NOR2_X1 NOR2_1522( .ZN(N4242), .A1(N4178), .A2(N4179) );
  NOR2_X1 NOR2_1523( .ZN(N4245), .A1(N4183), .A2(N4184) );
  NOR2_X1 NOR2_1524( .ZN(N4248), .A1(N4188), .A2(N4189) );
  NOR2_X1 NOR2_1525( .ZN(N4251), .A1(N4193), .A2(N4194) );
  NOR2_X1 NOR2_1526( .ZN(N4254), .A1(N4198), .A2(N4199) );
  NOR2_X1 NOR2_1527( .ZN(N4257), .A1(N4203), .A2(N4204) );
  NOR2_X1 NOR2_1528( .ZN(N4260), .A1(N4208), .A2(N4205) );
  NOR2_X1 NOR2_1529( .ZN(N4264), .A1(N4143), .A2(N4211) );
  NOR2_X1 NOR2_1530( .ZN(N4265), .A1(N4211), .A2(N4140) );
  NOR2_X1 NOR2_1531( .ZN(N4266), .A1(N4215), .A2(N4216) );
  NOR2_X1 NOR2_1532( .ZN(N4269), .A1(N4217), .A2(N1005) );
  NOR2_X1 NOR2_1533( .ZN(N4273), .A1(N4152), .A2(N4220) );
  NOR2_X1 NOR2_1534( .ZN(N4274), .A1(N4220), .A2(N1053) );
  NOR2_X1 NOR2_1535( .ZN(N4275), .A1(N4034), .A2(N4220) );
  NOR2_X1 NOR2_1536( .ZN(N4278), .A1(N4224), .A2(N4225) );
  NOR2_X1 NOR2_1537( .ZN(N4281), .A1(N4229), .A2(N4226) );
  NOR2_X1 NOR2_1538( .ZN(N4285), .A1(N4164), .A2(N4232) );
  NOR2_X1 NOR2_1539( .ZN(N4286), .A1(N4232), .A2(N4161) );
  NOR2_X1 NOR2_1540( .ZN(N4287), .A1(N4236), .A2(N4237) );
  NOR2_X1 NOR2_1541( .ZN(N4290), .A1(N4238), .A2(N1248) );
  NOR2_X1 NOR2_1542( .ZN(N4294), .A1(N4242), .A2(N4175) );
  NOR2_X1 NOR2_1543( .ZN(N4298), .A1(N4245), .A2(N4180) );
  NOR2_X1 NOR2_1544( .ZN(N4302), .A1(N4248), .A2(N4185) );
  NOR2_X1 NOR2_1545( .ZN(N4306), .A1(N4251), .A2(N4190) );
  NOR2_X1 NOR2_1546( .ZN(N4310), .A1(N4254), .A2(N4195) );
  NOR2_X1 NOR2_1547( .ZN(N4314), .A1(N4257), .A2(N4200) );
  NOR2_X1 NOR2_1548( .ZN(N4318), .A1(N4208), .A2(N4260) );
  NOR2_X1 NOR2_1549( .ZN(N4319), .A1(N4260), .A2(N4205) );
  NOR2_X1 NOR2_1550( .ZN(N4320), .A1(N4264), .A2(N4265) );
  NOR2_X1 NOR2_1551( .ZN(N4323), .A1(N4266), .A2(N957) );
  NOR2_X1 NOR2_1552( .ZN(N4327), .A1(N4217), .A2(N4269) );
  NOR2_X1 NOR2_1553( .ZN(N4328), .A1(N4269), .A2(N1005) );
  NOR2_X1 NOR2_1554( .ZN(N4329), .A1(N4085), .A2(N4269) );
  NOR2_X1 NOR2_1555( .ZN(N4332), .A1(N4273), .A2(N4274) );
  NOR2_X1 NOR2_1556( .ZN(N4335), .A1(N4278), .A2(N4275) );
  NOR2_X1 NOR2_1557( .ZN(N4339), .A1(N4229), .A2(N4281) );
  NOR2_X1 NOR2_1558( .ZN(N4340), .A1(N4281), .A2(N4226) );
  NOR2_X1 NOR2_1559( .ZN(N4341), .A1(N4285), .A2(N4286) );
  NOR2_X1 NOR2_1560( .ZN(N4344), .A1(N4287), .A2(N1200) );
  NOR2_X1 NOR2_1561( .ZN(N4348), .A1(N4238), .A2(N4290) );
  NOR2_X1 NOR2_1562( .ZN(N4349), .A1(N4290), .A2(N1248) );
  NOR2_X1 NOR2_1563( .ZN(N4350), .A1(N4106), .A2(N4290) );
  NOR2_X1 NOR2_1564( .ZN(N4353), .A1(N4242), .A2(N4294) );
  NOR2_X1 NOR2_1565( .ZN(N4354), .A1(N4294), .A2(N4175) );
  NOR2_X1 NOR2_1566( .ZN(N4355), .A1(N4245), .A2(N4298) );
  NOR2_X1 NOR2_1567( .ZN(N4356), .A1(N4298), .A2(N4180) );
  NOR2_X1 NOR2_1568( .ZN(N4357), .A1(N4248), .A2(N4302) );
  NOR2_X1 NOR2_1569( .ZN(N4358), .A1(N4302), .A2(N4185) );
  NOR2_X1 NOR2_1570( .ZN(N4359), .A1(N4251), .A2(N4306) );
  NOR2_X1 NOR2_1571( .ZN(N4360), .A1(N4306), .A2(N4190) );
  NOR2_X1 NOR2_1572( .ZN(N4361), .A1(N4254), .A2(N4310) );
  NOR2_X1 NOR2_1573( .ZN(N4362), .A1(N4310), .A2(N4195) );
  NOR2_X1 NOR2_1574( .ZN(N4363), .A1(N4257), .A2(N4314) );
  NOR2_X1 NOR2_1575( .ZN(N4364), .A1(N4314), .A2(N4200) );
  NOR2_X1 NOR2_1576( .ZN(N4365), .A1(N4318), .A2(N4319) );
  NOR2_X1 NOR2_1577( .ZN(N4368), .A1(N4320), .A2(N909) );
  NOR2_X1 NOR2_1578( .ZN(N4372), .A1(N4266), .A2(N4323) );
  NOR2_X1 NOR2_1579( .ZN(N4373), .A1(N4323), .A2(N957) );
  NOR2_X1 NOR2_1580( .ZN(N4374), .A1(N4146), .A2(N4323) );
  NOR2_X1 NOR2_1581( .ZN(N4377), .A1(N4327), .A2(N4328) );
  NOR2_X1 NOR2_1582( .ZN(N4380), .A1(N4332), .A2(N4329) );
  NOR2_X1 NOR2_1583( .ZN(N4384), .A1(N4278), .A2(N4335) );
  NOR2_X1 NOR2_1584( .ZN(N4385), .A1(N4335), .A2(N4275) );
  NOR2_X1 NOR2_1585( .ZN(N4386), .A1(N4339), .A2(N4340) );
  NOR2_X1 NOR2_1586( .ZN(N4389), .A1(N4341), .A2(N1152) );
  NOR2_X1 NOR2_1587( .ZN(N4393), .A1(N4287), .A2(N4344) );
  NOR2_X1 NOR2_1588( .ZN(N4394), .A1(N4344), .A2(N1200) );
  NOR2_X1 NOR2_1589( .ZN(N4395), .A1(N4167), .A2(N4344) );
  NOR2_X1 NOR2_1590( .ZN(N4398), .A1(N4348), .A2(N4349) );
  NOR2_X1 NOR2_1591( .ZN(N4401), .A1(N1296), .A2(N4350) );
  NOR2_X1 NOR2_1592( .ZN(N4405), .A1(N4353), .A2(N4354) );
  NOR2_X1 NOR2_1593( .ZN(N4408), .A1(N4355), .A2(N4356) );
  NOR2_X1 NOR2_1594( .ZN(N4411), .A1(N4357), .A2(N4358) );
  NOR2_X1 NOR2_1595( .ZN(N4414), .A1(N4359), .A2(N4360) );
  NOR2_X1 NOR2_1596( .ZN(N4417), .A1(N4361), .A2(N4362) );
  NOR2_X1 NOR2_1597( .ZN(N4420), .A1(N4363), .A2(N4364) );
  NOR2_X1 NOR2_1598( .ZN(N4423), .A1(N4365), .A2(N861) );
  NOR2_X1 NOR2_1599( .ZN(N4427), .A1(N4320), .A2(N4368) );
  NOR2_X1 NOR2_1600( .ZN(N4428), .A1(N4368), .A2(N909) );
  NOR2_X1 NOR2_1601( .ZN(N4429), .A1(N4211), .A2(N4368) );
  NOR2_X1 NOR2_1602( .ZN(N4432), .A1(N4372), .A2(N4373) );
  NOR2_X1 NOR2_1603( .ZN(N4435), .A1(N4377), .A2(N4374) );
  NOR2_X1 NOR2_1604( .ZN(N4439), .A1(N4332), .A2(N4380) );
  NOR2_X1 NOR2_1605( .ZN(N4440), .A1(N4380), .A2(N4329) );
  NOR2_X1 NOR2_1606( .ZN(N4441), .A1(N4384), .A2(N4385) );
  NOR2_X1 NOR2_1607( .ZN(N4444), .A1(N4386), .A2(N1104) );
  NOR2_X1 NOR2_1608( .ZN(N4448), .A1(N4341), .A2(N4389) );
  NOR2_X1 NOR2_1609( .ZN(N4449), .A1(N4389), .A2(N1152) );
  NOR2_X1 NOR2_1610( .ZN(N4450), .A1(N4232), .A2(N4389) );
  NOR2_X1 NOR2_1611( .ZN(N4453), .A1(N4393), .A2(N4394) );
  NOR2_X1 NOR2_1612( .ZN(N4456), .A1(N4398), .A2(N4395) );
  NOR2_X1 NOR2_1613( .ZN(N4460), .A1(N1296), .A2(N4401) );
  NOR2_X1 NOR2_1614( .ZN(N4461), .A1(N4401), .A2(N4350) );
  NOR2_X1 NOR2_1615( .ZN(N4462), .A1(N4405), .A2(N573) );
  NOR2_X1 NOR2_1616( .ZN(N4466), .A1(N4408), .A2(N621) );
  NOR2_X1 NOR2_1617( .ZN(N4470), .A1(N4411), .A2(N669) );
  NOR2_X1 NOR2_1618( .ZN(N4474), .A1(N4414), .A2(N717) );
  NOR2_X1 NOR2_1619( .ZN(N4478), .A1(N4417), .A2(N765) );
  NOR2_X1 NOR2_1620( .ZN(N4482), .A1(N4420), .A2(N813) );
  NOR2_X1 NOR2_1621( .ZN(N4486), .A1(N4365), .A2(N4423) );
  NOR2_X1 NOR2_1622( .ZN(N4487), .A1(N4423), .A2(N861) );
  NOR2_X1 NOR2_1623( .ZN(N4488), .A1(N4260), .A2(N4423) );
  NOR2_X1 NOR2_1624( .ZN(N4491), .A1(N4427), .A2(N4428) );
  NOR2_X1 NOR2_1625( .ZN(N4494), .A1(N4432), .A2(N4429) );
  NOR2_X1 NOR2_1626( .ZN(N4498), .A1(N4377), .A2(N4435) );
  NOR2_X1 NOR2_1627( .ZN(N4499), .A1(N4435), .A2(N4374) );
  NOR2_X1 NOR2_1628( .ZN(N4500), .A1(N4439), .A2(N4440) );
  NOR2_X1 NOR2_1629( .ZN(N4503), .A1(N4441), .A2(N1056) );
  NOR2_X1 NOR2_1630( .ZN(N4507), .A1(N4386), .A2(N4444) );
  NOR2_X1 NOR2_1631( .ZN(N4508), .A1(N4444), .A2(N1104) );
  NOR2_X1 NOR2_1632( .ZN(N4509), .A1(N4281), .A2(N4444) );
  NOR2_X1 NOR2_1633( .ZN(N4512), .A1(N4448), .A2(N4449) );
  NOR2_X1 NOR2_1634( .ZN(N4515), .A1(N4453), .A2(N4450) );
  NOR2_X1 NOR2_1635( .ZN(N4519), .A1(N4398), .A2(N4456) );
  NOR2_X1 NOR2_1636( .ZN(N4520), .A1(N4456), .A2(N4395) );
  NOR2_X1 NOR2_1637( .ZN(N4521), .A1(N4460), .A2(N4461) );
  NOR2_X1 NOR2_1638( .ZN(N4524), .A1(N4405), .A2(N4462) );
  NOR2_X1 NOR2_1639( .ZN(N4525), .A1(N4462), .A2(N573) );
  NOR2_X1 NOR2_1640( .ZN(N4526), .A1(N4294), .A2(N4462) );
  NOR2_X1 NOR2_1641( .ZN(N4529), .A1(N4408), .A2(N4466) );
  NOR2_X1 NOR2_1642( .ZN(N4530), .A1(N4466), .A2(N621) );
  NOR2_X1 NOR2_1643( .ZN(N4531), .A1(N4298), .A2(N4466) );
  NOR2_X1 NOR2_1644( .ZN(N4534), .A1(N4411), .A2(N4470) );
  NOR2_X1 NOR2_1645( .ZN(N4535), .A1(N4470), .A2(N669) );
  NOR2_X1 NOR2_1646( .ZN(N4536), .A1(N4302), .A2(N4470) );
  NOR2_X1 NOR2_1647( .ZN(N4539), .A1(N4414), .A2(N4474) );
  NOR2_X1 NOR2_1648( .ZN(N4540), .A1(N4474), .A2(N717) );
  NOR2_X1 NOR2_1649( .ZN(N4541), .A1(N4306), .A2(N4474) );
  NOR2_X1 NOR2_1650( .ZN(N4544), .A1(N4417), .A2(N4478) );
  NOR2_X1 NOR2_1651( .ZN(N4545), .A1(N4478), .A2(N765) );
  NOR2_X1 NOR2_1652( .ZN(N4546), .A1(N4310), .A2(N4478) );
  NOR2_X1 NOR2_1653( .ZN(N4549), .A1(N4420), .A2(N4482) );
  NOR2_X1 NOR2_1654( .ZN(N4550), .A1(N4482), .A2(N813) );
  NOR2_X1 NOR2_1655( .ZN(N4551), .A1(N4314), .A2(N4482) );
  NOR2_X1 NOR2_1656( .ZN(N4554), .A1(N4486), .A2(N4487) );
  NOR2_X1 NOR2_1657( .ZN(N4557), .A1(N4491), .A2(N4488) );
  NOR2_X1 NOR2_1658( .ZN(N4561), .A1(N4432), .A2(N4494) );
  NOR2_X1 NOR2_1659( .ZN(N4562), .A1(N4494), .A2(N4429) );
  NOR2_X1 NOR2_1660( .ZN(N4563), .A1(N4498), .A2(N4499) );
  NOR2_X1 NOR2_1661( .ZN(N4566), .A1(N4500), .A2(N1008) );
  NOR2_X1 NOR2_1662( .ZN(N4570), .A1(N4441), .A2(N4503) );
  NOR2_X1 NOR2_1663( .ZN(N4571), .A1(N4503), .A2(N1056) );
  NOR2_X1 NOR2_1664( .ZN(N4572), .A1(N4335), .A2(N4503) );
  NOR2_X1 NOR2_1665( .ZN(N4575), .A1(N4507), .A2(N4508) );
  NOR2_X1 NOR2_1666( .ZN(N4578), .A1(N4512), .A2(N4509) );
  NOR2_X1 NOR2_1667( .ZN(N4582), .A1(N4453), .A2(N4515) );
  NOR2_X1 NOR2_1668( .ZN(N4583), .A1(N4515), .A2(N4450) );
  NOR2_X1 NOR2_1669( .ZN(N4584), .A1(N4519), .A2(N4520) );
  NOR2_X1 NOR2_1670( .ZN(N4587), .A1(N4521), .A2(N1251) );
  NOR2_X1 NOR2_1671( .ZN(N4591), .A1(N4524), .A2(N4525) );
  NOR2_X1 NOR2_1672( .ZN(N4592), .A1(N4529), .A2(N4530) );
  NOR2_X1 NOR2_1673( .ZN(N4595), .A1(N4534), .A2(N4535) );
  NOR2_X1 NOR2_1674( .ZN(N4598), .A1(N4539), .A2(N4540) );
  NOR2_X1 NOR2_1675( .ZN(N4601), .A1(N4544), .A2(N4545) );
  NOR2_X1 NOR2_1676( .ZN(N4604), .A1(N4549), .A2(N4550) );
  NOR2_X1 NOR2_1677( .ZN(N4607), .A1(N4554), .A2(N4551) );
  NOR2_X1 NOR2_1678( .ZN(N4611), .A1(N4491), .A2(N4557) );
  NOR2_X1 NOR2_1679( .ZN(N4612), .A1(N4557), .A2(N4488) );
  NOR2_X1 NOR2_1680( .ZN(N4613), .A1(N4561), .A2(N4562) );
  NOR2_X1 NOR2_1681( .ZN(N4616), .A1(N4563), .A2(N960) );
  NOR2_X1 NOR2_1682( .ZN(N4620), .A1(N4500), .A2(N4566) );
  NOR2_X1 NOR2_1683( .ZN(N4621), .A1(N4566), .A2(N1008) );
  NOR2_X1 NOR2_1684( .ZN(N4622), .A1(N4380), .A2(N4566) );
  NOR2_X1 NOR2_1685( .ZN(N4625), .A1(N4570), .A2(N4571) );
  NOR2_X1 NOR2_1686( .ZN(N4628), .A1(N4575), .A2(N4572) );
  NOR2_X1 NOR2_1687( .ZN(N4632), .A1(N4512), .A2(N4578) );
  NOR2_X1 NOR2_1688( .ZN(N4633), .A1(N4578), .A2(N4509) );
  NOR2_X1 NOR2_1689( .ZN(N4634), .A1(N4582), .A2(N4583) );
  NOR2_X1 NOR2_1690( .ZN(N4637), .A1(N4584), .A2(N1203) );
  NOR2_X1 NOR2_1691( .ZN(N4641), .A1(N4521), .A2(N4587) );
  NOR2_X1 NOR2_1692( .ZN(N4642), .A1(N4587), .A2(N1251) );
  NOR2_X1 NOR2_1693( .ZN(N4643), .A1(N4401), .A2(N4587) );
  NOR2_X1 NOR2_1694( .ZN(N4646), .A1(N4592), .A2(N4526) );
  NOR2_X1 NOR2_1695( .ZN(N4650), .A1(N4595), .A2(N4531) );
  NOR2_X1 NOR2_1696( .ZN(N4654), .A1(N4598), .A2(N4536) );
  NOR2_X1 NOR2_1697( .ZN(N4658), .A1(N4601), .A2(N4541) );
  NOR2_X1 NOR2_1698( .ZN(N4662), .A1(N4604), .A2(N4546) );
  NOR2_X1 NOR2_1699( .ZN(N4666), .A1(N4554), .A2(N4607) );
  NOR2_X1 NOR2_1700( .ZN(N4667), .A1(N4607), .A2(N4551) );
  NOR2_X1 NOR2_1701( .ZN(N4668), .A1(N4611), .A2(N4612) );
  NOR2_X1 NOR2_1702( .ZN(N4671), .A1(N4613), .A2(N912) );
  NOR2_X1 NOR2_1703( .ZN(N4675), .A1(N4563), .A2(N4616) );
  NOR2_X1 NOR2_1704( .ZN(N4676), .A1(N4616), .A2(N960) );
  NOR2_X1 NOR2_1705( .ZN(N4677), .A1(N4435), .A2(N4616) );
  NOR2_X1 NOR2_1706( .ZN(N4680), .A1(N4620), .A2(N4621) );
  NOR2_X1 NOR2_1707( .ZN(N4683), .A1(N4625), .A2(N4622) );
  NOR2_X1 NOR2_1708( .ZN(N4687), .A1(N4575), .A2(N4628) );
  NOR2_X1 NOR2_1709( .ZN(N4688), .A1(N4628), .A2(N4572) );
  NOR2_X1 NOR2_1710( .ZN(N4689), .A1(N4632), .A2(N4633) );
  NOR2_X1 NOR2_1711( .ZN(N4692), .A1(N4634), .A2(N1155) );
  NOR2_X1 NOR2_1712( .ZN(N4696), .A1(N4584), .A2(N4637) );
  NOR2_X1 NOR2_1713( .ZN(N4697), .A1(N4637), .A2(N1203) );
  NOR2_X1 NOR2_1714( .ZN(N4698), .A1(N4456), .A2(N4637) );
  NOR2_X1 NOR2_1715( .ZN(N4701), .A1(N4641), .A2(N4642) );
  NOR2_X1 NOR2_1716( .ZN(N4704), .A1(N1299), .A2(N4643) );
  NOR2_X1 NOR2_1717( .ZN(N4708), .A1(N4592), .A2(N4646) );
  NOR2_X1 NOR2_1718( .ZN(N4709), .A1(N4646), .A2(N4526) );
  NOR2_X1 NOR2_1719( .ZN(N4710), .A1(N4595), .A2(N4650) );
  NOR2_X1 NOR2_1720( .ZN(N4711), .A1(N4650), .A2(N4531) );
  NOR2_X1 NOR2_1721( .ZN(N4712), .A1(N4598), .A2(N4654) );
  NOR2_X1 NOR2_1722( .ZN(N4713), .A1(N4654), .A2(N4536) );
  NOR2_X1 NOR2_1723( .ZN(N4714), .A1(N4601), .A2(N4658) );
  NOR2_X1 NOR2_1724( .ZN(N4715), .A1(N4658), .A2(N4541) );
  NOR2_X1 NOR2_1725( .ZN(N4716), .A1(N4604), .A2(N4662) );
  NOR2_X1 NOR2_1726( .ZN(N4717), .A1(N4662), .A2(N4546) );
  NOR2_X1 NOR2_1727( .ZN(N4718), .A1(N4666), .A2(N4667) );
  NOR2_X1 NOR2_1728( .ZN(N4721), .A1(N4668), .A2(N864) );
  NOR2_X1 NOR2_1729( .ZN(N4725), .A1(N4613), .A2(N4671) );
  NOR2_X1 NOR2_1730( .ZN(N4726), .A1(N4671), .A2(N912) );
  NOR2_X1 NOR2_1731( .ZN(N4727), .A1(N4494), .A2(N4671) );
  NOR2_X1 NOR2_1732( .ZN(N4730), .A1(N4675), .A2(N4676) );
  NOR2_X1 NOR2_1733( .ZN(N4733), .A1(N4680), .A2(N4677) );
  NOR2_X1 NOR2_1734( .ZN(N4737), .A1(N4625), .A2(N4683) );
  NOR2_X1 NOR2_1735( .ZN(N4738), .A1(N4683), .A2(N4622) );
  NOR2_X1 NOR2_1736( .ZN(N4739), .A1(N4687), .A2(N4688) );
  NOR2_X1 NOR2_1737( .ZN(N4742), .A1(N4689), .A2(N1107) );
  NOR2_X1 NOR2_1738( .ZN(N4746), .A1(N4634), .A2(N4692) );
  NOR2_X1 NOR2_1739( .ZN(N4747), .A1(N4692), .A2(N1155) );
  NOR2_X1 NOR2_1740( .ZN(N4748), .A1(N4515), .A2(N4692) );
  NOR2_X1 NOR2_1741( .ZN(N4751), .A1(N4696), .A2(N4697) );
  NOR2_X2 NOR2_1742( .ZN(N4754), .A1(N4701), .A2(N4698) );
  NOR2_X2 NOR2_1743( .ZN(N4758), .A1(N1299), .A2(N4704) );
  NOR2_X2 NOR2_1744( .ZN(N4759), .A1(N4704), .A2(N4643) );
  NOR2_X2 NOR2_1745( .ZN(N4760), .A1(N4708), .A2(N4709) );
  NOR2_X2 NOR2_1746( .ZN(N4763), .A1(N4710), .A2(N4711) );
  NOR2_X2 NOR2_1747( .ZN(N4766), .A1(N4712), .A2(N4713) );
  NOR2_X2 NOR2_1748( .ZN(N4769), .A1(N4714), .A2(N4715) );
  NOR2_X2 NOR2_1749( .ZN(N4772), .A1(N4716), .A2(N4717) );
  NOR2_X2 NOR2_1750( .ZN(N4775), .A1(N4718), .A2(N816) );
  NOR2_X1 NOR2_1751( .ZN(N4779), .A1(N4668), .A2(N4721) );
  NOR2_X1 NOR2_1752( .ZN(N4780), .A1(N4721), .A2(N864) );
  NOR2_X1 NOR2_1753( .ZN(N4781), .A1(N4557), .A2(N4721) );
  NOR2_X1 NOR2_1754( .ZN(N4784), .A1(N4725), .A2(N4726) );
  NOR2_X1 NOR2_1755( .ZN(N4787), .A1(N4730), .A2(N4727) );
  NOR2_X1 NOR2_1756( .ZN(N4791), .A1(N4680), .A2(N4733) );
  NOR2_X1 NOR2_1757( .ZN(N4792), .A1(N4733), .A2(N4677) );
  NOR2_X1 NOR2_1758( .ZN(N4793), .A1(N4737), .A2(N4738) );
  NOR2_X1 NOR2_1759( .ZN(N4796), .A1(N4739), .A2(N1059) );
  NOR2_X1 NOR2_1760( .ZN(N4800), .A1(N4689), .A2(N4742) );
  NOR2_X1 NOR2_1761( .ZN(N4801), .A1(N4742), .A2(N1107) );
  NOR2_X1 NOR2_1762( .ZN(N4802), .A1(N4578), .A2(N4742) );
  NOR2_X1 NOR2_1763( .ZN(N4805), .A1(N4746), .A2(N4747) );
  NOR2_X1 NOR2_1764( .ZN(N4808), .A1(N4751), .A2(N4748) );
  NOR2_X1 NOR2_1765( .ZN(N4812), .A1(N4701), .A2(N4754) );
  NOR2_X1 NOR2_1766( .ZN(N4813), .A1(N4754), .A2(N4698) );
  NOR2_X1 NOR2_1767( .ZN(N4814), .A1(N4758), .A2(N4759) );
  NOR2_X1 NOR2_1768( .ZN(N4817), .A1(N4760), .A2(N576) );
  NOR2_X1 NOR2_1769( .ZN(N4821), .A1(N4763), .A2(N624) );
  NOR2_X1 NOR2_1770( .ZN(N4825), .A1(N4766), .A2(N672) );
  NOR2_X1 NOR2_1771( .ZN(N4829), .A1(N4769), .A2(N720) );
  NOR2_X1 NOR2_1772( .ZN(N4833), .A1(N4772), .A2(N768) );
  NOR2_X1 NOR2_1773( .ZN(N4837), .A1(N4718), .A2(N4775) );
  NOR2_X1 NOR2_1774( .ZN(N4838), .A1(N4775), .A2(N816) );
  NOR2_X1 NOR2_1775( .ZN(N4839), .A1(N4607), .A2(N4775) );
  NOR2_X1 NOR2_1776( .ZN(N4842), .A1(N4779), .A2(N4780) );
  NOR2_X1 NOR2_1777( .ZN(N4845), .A1(N4784), .A2(N4781) );
  NOR2_X1 NOR2_1778( .ZN(N4849), .A1(N4730), .A2(N4787) );
  NOR2_X1 NOR2_1779( .ZN(N4850), .A1(N4787), .A2(N4727) );
  NOR2_X1 NOR2_1780( .ZN(N4851), .A1(N4791), .A2(N4792) );
  NOR2_X1 NOR2_1781( .ZN(N4854), .A1(N4793), .A2(N1011) );
  NOR2_X1 NOR2_1782( .ZN(N4858), .A1(N4739), .A2(N4796) );
  NOR2_X1 NOR2_1783( .ZN(N4859), .A1(N4796), .A2(N1059) );
  NOR2_X1 NOR2_1784( .ZN(N4860), .A1(N4628), .A2(N4796) );
  NOR2_X1 NOR2_1785( .ZN(N4863), .A1(N4800), .A2(N4801) );
  NOR2_X1 NOR2_1786( .ZN(N4866), .A1(N4805), .A2(N4802) );
  NOR2_X1 NOR2_1787( .ZN(N4870), .A1(N4751), .A2(N4808) );
  NOR2_X1 NOR2_1788( .ZN(N4871), .A1(N4808), .A2(N4748) );
  NOR2_X1 NOR2_1789( .ZN(N4872), .A1(N4812), .A2(N4813) );
  NOR2_X1 NOR2_1790( .ZN(N4875), .A1(N4814), .A2(N1254) );
  NOR2_X1 NOR2_1791( .ZN(N4879), .A1(N4760), .A2(N4817) );
  NOR2_X1 NOR2_1792( .ZN(N4880), .A1(N4817), .A2(N576) );
  NOR2_X1 NOR2_1793( .ZN(N4881), .A1(N4646), .A2(N4817) );
  NOR2_X1 NOR2_1794( .ZN(N4884), .A1(N4763), .A2(N4821) );
  NOR2_X1 NOR2_1795( .ZN(N4885), .A1(N4821), .A2(N624) );
  NOR2_X1 NOR2_1796( .ZN(N4886), .A1(N4650), .A2(N4821) );
  NOR2_X1 NOR2_1797( .ZN(N4889), .A1(N4766), .A2(N4825) );
  NOR2_X1 NOR2_1798( .ZN(N4890), .A1(N4825), .A2(N672) );
  NOR2_X1 NOR2_1799( .ZN(N4891), .A1(N4654), .A2(N4825) );
  NOR2_X1 NOR2_1800( .ZN(N4894), .A1(N4769), .A2(N4829) );
  NOR2_X1 NOR2_1801( .ZN(N4895), .A1(N4829), .A2(N720) );
  NOR2_X1 NOR2_1802( .ZN(N4896), .A1(N4658), .A2(N4829) );
  NOR2_X1 NOR2_1803( .ZN(N4899), .A1(N4772), .A2(N4833) );
  NOR2_X1 NOR2_1804( .ZN(N4900), .A1(N4833), .A2(N768) );
  NOR2_X1 NOR2_1805( .ZN(N4901), .A1(N4662), .A2(N4833) );
  NOR2_X1 NOR2_1806( .ZN(N4904), .A1(N4837), .A2(N4838) );
  NOR2_X1 NOR2_1807( .ZN(N4907), .A1(N4842), .A2(N4839) );
  NOR2_X1 NOR2_1808( .ZN(N4911), .A1(N4784), .A2(N4845) );
  NOR2_X1 NOR2_1809( .ZN(N4912), .A1(N4845), .A2(N4781) );
  NOR2_X1 NOR2_1810( .ZN(N4913), .A1(N4849), .A2(N4850) );
  NOR2_X1 NOR2_1811( .ZN(N4916), .A1(N4851), .A2(N963) );
  NOR2_X1 NOR2_1812( .ZN(N4920), .A1(N4793), .A2(N4854) );
  NOR2_X1 NOR2_1813( .ZN(N4921), .A1(N4854), .A2(N1011) );
  NOR2_X1 NOR2_1814( .ZN(N4922), .A1(N4683), .A2(N4854) );
  NOR2_X1 NOR2_1815( .ZN(N4925), .A1(N4858), .A2(N4859) );
  NOR2_X1 NOR2_1816( .ZN(N4928), .A1(N4863), .A2(N4860) );
  NOR2_X1 NOR2_1817( .ZN(N4932), .A1(N4805), .A2(N4866) );
  NOR2_X1 NOR2_1818( .ZN(N4933), .A1(N4866), .A2(N4802) );
  NOR2_X1 NOR2_1819( .ZN(N4934), .A1(N4870), .A2(N4871) );
  NOR2_X1 NOR2_1820( .ZN(N4937), .A1(N4872), .A2(N1206) );
  NOR2_X1 NOR2_1821( .ZN(N4941), .A1(N4814), .A2(N4875) );
  NOR2_X1 NOR2_1822( .ZN(N4942), .A1(N4875), .A2(N1254) );
  NOR2_X1 NOR2_1823( .ZN(N4943), .A1(N4704), .A2(N4875) );
  NOR2_X1 NOR2_1824( .ZN(N4946), .A1(N4879), .A2(N4880) );
  NOR2_X1 NOR2_1825( .ZN(N4947), .A1(N4884), .A2(N4885) );
  NOR2_X1 NOR2_1826( .ZN(N4950), .A1(N4889), .A2(N4890) );
  NOR2_X1 NOR2_1827( .ZN(N4953), .A1(N4894), .A2(N4895) );
  NOR2_X1 NOR2_1828( .ZN(N4956), .A1(N4899), .A2(N4900) );
  NOR2_X1 NOR2_1829( .ZN(N4959), .A1(N4904), .A2(N4901) );
  NOR2_X1 NOR2_1830( .ZN(N4963), .A1(N4842), .A2(N4907) );
  NOR2_X1 NOR2_1831( .ZN(N4964), .A1(N4907), .A2(N4839) );
  NOR2_X1 NOR2_1832( .ZN(N4965), .A1(N4911), .A2(N4912) );
  NOR2_X1 NOR2_1833( .ZN(N4968), .A1(N4913), .A2(N915) );
  NOR2_X1 NOR2_1834( .ZN(N4972), .A1(N4851), .A2(N4916) );
  NOR2_X1 NOR2_1835( .ZN(N4973), .A1(N4916), .A2(N963) );
  NOR2_X1 NOR2_1836( .ZN(N4974), .A1(N4733), .A2(N4916) );
  NOR2_X1 NOR2_1837( .ZN(N4977), .A1(N4920), .A2(N4921) );
  NOR2_X1 NOR2_1838( .ZN(N4980), .A1(N4925), .A2(N4922) );
  NOR2_X1 NOR2_1839( .ZN(N4984), .A1(N4863), .A2(N4928) );
  NOR2_X1 NOR2_1840( .ZN(N4985), .A1(N4928), .A2(N4860) );
  NOR2_X1 NOR2_1841( .ZN(N4986), .A1(N4932), .A2(N4933) );
  NOR2_X1 NOR2_1842( .ZN(N4989), .A1(N4934), .A2(N1158) );
  NOR2_X1 NOR2_1843( .ZN(N4993), .A1(N4872), .A2(N4937) );
  NOR2_X1 NOR2_1844( .ZN(N4994), .A1(N4937), .A2(N1206) );
  NOR2_X1 NOR2_1845( .ZN(N4995), .A1(N4754), .A2(N4937) );
  NOR2_X1 NOR2_1846( .ZN(N4998), .A1(N4941), .A2(N4942) );
  NOR2_X1 NOR2_1847( .ZN(N5001), .A1(N1302), .A2(N4943) );
  NOR2_X1 NOR2_1848( .ZN(N5005), .A1(N4947), .A2(N4881) );
  NOR2_X1 NOR2_1849( .ZN(N5009), .A1(N4950), .A2(N4886) );
  NOR2_X1 NOR2_1850( .ZN(N5013), .A1(N4953), .A2(N4891) );
  NOR2_X1 NOR2_1851( .ZN(N5017), .A1(N4956), .A2(N4896) );
  NOR2_X1 NOR2_1852( .ZN(N5021), .A1(N4904), .A2(N4959) );
  NOR2_X1 NOR2_1853( .ZN(N5022), .A1(N4959), .A2(N4901) );
  NOR2_X1 NOR2_1854( .ZN(N5023), .A1(N4963), .A2(N4964) );
  NOR2_X1 NOR2_1855( .ZN(N5026), .A1(N4965), .A2(N867) );
  NOR2_X1 NOR2_1856( .ZN(N5030), .A1(N4913), .A2(N4968) );
  NOR2_X1 NOR2_1857( .ZN(N5031), .A1(N4968), .A2(N915) );
  NOR2_X1 NOR2_1858( .ZN(N5032), .A1(N4787), .A2(N4968) );
  NOR2_X1 NOR2_1859( .ZN(N5035), .A1(N4972), .A2(N4973) );
  NOR2_X1 NOR2_1860( .ZN(N5038), .A1(N4977), .A2(N4974) );
  NOR2_X1 NOR2_1861( .ZN(N5042), .A1(N4925), .A2(N4980) );
  NOR2_X1 NOR2_1862( .ZN(N5043), .A1(N4980), .A2(N4922) );
  NOR2_X1 NOR2_1863( .ZN(N5044), .A1(N4984), .A2(N4985) );
  NOR2_X1 NOR2_1864( .ZN(N5047), .A1(N4986), .A2(N1110) );
  NOR2_X1 NOR2_1865( .ZN(N5051), .A1(N4934), .A2(N4989) );
  NOR2_X1 NOR2_1866( .ZN(N5052), .A1(N4989), .A2(N1158) );
  NOR2_X1 NOR2_1867( .ZN(N5053), .A1(N4808), .A2(N4989) );
  NOR2_X1 NOR2_1868( .ZN(N5056), .A1(N4993), .A2(N4994) );
  NOR2_X1 NOR2_1869( .ZN(N5059), .A1(N4998), .A2(N4995) );
  NOR2_X1 NOR2_1870( .ZN(N5063), .A1(N1302), .A2(N5001) );
  NOR2_X1 NOR2_1871( .ZN(N5064), .A1(N5001), .A2(N4943) );
  NOR2_X1 NOR2_1872( .ZN(N5065), .A1(N4947), .A2(N5005) );
  NOR2_X1 NOR2_1873( .ZN(N5066), .A1(N5005), .A2(N4881) );
  NOR2_X1 NOR2_1874( .ZN(N5067), .A1(N4950), .A2(N5009) );
  NOR2_X1 NOR2_1875( .ZN(N5068), .A1(N5009), .A2(N4886) );
  NOR2_X1 NOR2_1876( .ZN(N5069), .A1(N4953), .A2(N5013) );
  NOR2_X1 NOR2_1877( .ZN(N5070), .A1(N5013), .A2(N4891) );
  NOR2_X1 NOR2_1878( .ZN(N5071), .A1(N4956), .A2(N5017) );
  NOR2_X1 NOR2_1879( .ZN(N5072), .A1(N5017), .A2(N4896) );
  NOR2_X1 NOR2_1880( .ZN(N5073), .A1(N5021), .A2(N5022) );
  NOR2_X1 NOR2_1881( .ZN(N5076), .A1(N5023), .A2(N819) );
  NOR2_X1 NOR2_1882( .ZN(N5080), .A1(N4965), .A2(N5026) );
  NOR2_X1 NOR2_1883( .ZN(N5081), .A1(N5026), .A2(N867) );
  NOR2_X1 NOR2_1884( .ZN(N5082), .A1(N4845), .A2(N5026) );
  NOR2_X1 NOR2_1885( .ZN(N5085), .A1(N5030), .A2(N5031) );
  NOR2_X1 NOR2_1886( .ZN(N5088), .A1(N5035), .A2(N5032) );
  NOR2_X1 NOR2_1887( .ZN(N5092), .A1(N4977), .A2(N5038) );
  NOR2_X1 NOR2_1888( .ZN(N5093), .A1(N5038), .A2(N4974) );
  NOR2_X1 NOR2_1889( .ZN(N5094), .A1(N5042), .A2(N5043) );
  NOR2_X1 NOR2_1890( .ZN(N5097), .A1(N5044), .A2(N1062) );
  NOR2_X1 NOR2_1891( .ZN(N5101), .A1(N4986), .A2(N5047) );
  NOR2_X1 NOR2_1892( .ZN(N5102), .A1(N5047), .A2(N1110) );
  NOR2_X1 NOR2_1893( .ZN(N5103), .A1(N4866), .A2(N5047) );
  NOR2_X1 NOR2_1894( .ZN(N5106), .A1(N5051), .A2(N5052) );
  NOR2_X1 NOR2_1895( .ZN(N5109), .A1(N5056), .A2(N5053) );
  NOR2_X1 NOR2_1896( .ZN(N5113), .A1(N4998), .A2(N5059) );
  NOR2_X1 NOR2_1897( .ZN(N5114), .A1(N5059), .A2(N4995) );
  NOR2_X1 NOR2_1898( .ZN(N5115), .A1(N5063), .A2(N5064) );
  NOR2_X1 NOR2_1899( .ZN(N5118), .A1(N5065), .A2(N5066) );
  NOR2_X1 NOR2_1900( .ZN(N5121), .A1(N5067), .A2(N5068) );
  NOR2_X1 NOR2_1901( .ZN(N5124), .A1(N5069), .A2(N5070) );
  NOR2_X1 NOR2_1902( .ZN(N5127), .A1(N5071), .A2(N5072) );
  NOR2_X1 NOR2_1903( .ZN(N5130), .A1(N5073), .A2(N771) );
  NOR2_X1 NOR2_1904( .ZN(N5134), .A1(N5023), .A2(N5076) );
  NOR2_X1 NOR2_1905( .ZN(N5135), .A1(N5076), .A2(N819) );
  NOR2_X1 NOR2_1906( .ZN(N5136), .A1(N4907), .A2(N5076) );
  NOR2_X1 NOR2_1907( .ZN(N5139), .A1(N5080), .A2(N5081) );
  NOR2_X1 NOR2_1908( .ZN(N5142), .A1(N5085), .A2(N5082) );
  NOR2_X1 NOR2_1909( .ZN(N5146), .A1(N5035), .A2(N5088) );
  NOR2_X1 NOR2_1910( .ZN(N5147), .A1(N5088), .A2(N5032) );
  NOR2_X1 NOR2_1911( .ZN(N5148), .A1(N5092), .A2(N5093) );
  NOR2_X1 NOR2_1912( .ZN(N5151), .A1(N5094), .A2(N1014) );
  NOR2_X1 NOR2_1913( .ZN(N5155), .A1(N5044), .A2(N5097) );
  NOR2_X1 NOR2_1914( .ZN(N5156), .A1(N5097), .A2(N1062) );
  NOR2_X1 NOR2_1915( .ZN(N5157), .A1(N4928), .A2(N5097) );
  NOR2_X1 NOR2_1916( .ZN(N5160), .A1(N5101), .A2(N5102) );
  NOR2_X1 NOR2_1917( .ZN(N5163), .A1(N5106), .A2(N5103) );
  NOR2_X1 NOR2_1918( .ZN(N5167), .A1(N5056), .A2(N5109) );
  NOR2_X1 NOR2_1919( .ZN(N5168), .A1(N5109), .A2(N5053) );
  NOR2_X1 NOR2_1920( .ZN(N5169), .A1(N5113), .A2(N5114) );
  NOR2_X1 NOR2_1921( .ZN(N5172), .A1(N5115), .A2(N1257) );
  NOR2_X1 NOR2_1922( .ZN(N5176), .A1(N5118), .A2(N579) );
  NOR2_X1 NOR2_1923( .ZN(N5180), .A1(N5121), .A2(N627) );
  NOR2_X1 NOR2_1924( .ZN(N5184), .A1(N5124), .A2(N675) );
  NOR2_X1 NOR2_1925( .ZN(N5188), .A1(N5127), .A2(N723) );
  NOR2_X1 NOR2_1926( .ZN(N5192), .A1(N5073), .A2(N5130) );
  NOR2_X1 NOR2_1927( .ZN(N5193), .A1(N5130), .A2(N771) );
  NOR2_X1 NOR2_1928( .ZN(N5194), .A1(N4959), .A2(N5130) );
  NOR2_X1 NOR2_1929( .ZN(N5197), .A1(N5134), .A2(N5135) );
  NOR2_X1 NOR2_1930( .ZN(N5200), .A1(N5139), .A2(N5136) );
  NOR2_X1 NOR2_1931( .ZN(N5204), .A1(N5085), .A2(N5142) );
  NOR2_X1 NOR2_1932( .ZN(N5205), .A1(N5142), .A2(N5082) );
  NOR2_X1 NOR2_1933( .ZN(N5206), .A1(N5146), .A2(N5147) );
  NOR2_X1 NOR2_1934( .ZN(N5209), .A1(N5148), .A2(N966) );
  NOR2_X1 NOR2_1935( .ZN(N5213), .A1(N5094), .A2(N5151) );
  NOR2_X1 NOR2_1936( .ZN(N5214), .A1(N5151), .A2(N1014) );
  NOR2_X1 NOR2_1937( .ZN(N5215), .A1(N4980), .A2(N5151) );
  NOR2_X1 NOR2_1938( .ZN(N5218), .A1(N5155), .A2(N5156) );
  NOR2_X1 NOR2_1939( .ZN(N5221), .A1(N5160), .A2(N5157) );
  NOR2_X1 NOR2_1940( .ZN(N5225), .A1(N5106), .A2(N5163) );
  NOR2_X1 NOR2_1941( .ZN(N5226), .A1(N5163), .A2(N5103) );
  NOR2_X1 NOR2_1942( .ZN(N5227), .A1(N5167), .A2(N5168) );
  NOR2_X1 NOR2_1943( .ZN(N5230), .A1(N5169), .A2(N1209) );
  NOR2_X1 NOR2_1944( .ZN(N5234), .A1(N5115), .A2(N5172) );
  NOR2_X1 NOR2_1945( .ZN(N5235), .A1(N5172), .A2(N1257) );
  NOR2_X1 NOR2_1946( .ZN(N5236), .A1(N5001), .A2(N5172) );
  NOR2_X1 NOR2_1947( .ZN(N5239), .A1(N5118), .A2(N5176) );
  NOR2_X1 NOR2_1948( .ZN(N5240), .A1(N5176), .A2(N579) );
  NOR2_X1 NOR2_1949( .ZN(N5241), .A1(N5005), .A2(N5176) );
  NOR2_X1 NOR2_1950( .ZN(N5244), .A1(N5121), .A2(N5180) );
  NOR2_X1 NOR2_1951( .ZN(N5245), .A1(N5180), .A2(N627) );
  NOR2_X1 NOR2_1952( .ZN(N5246), .A1(N5009), .A2(N5180) );
  NOR2_X1 NOR2_1953( .ZN(N5249), .A1(N5124), .A2(N5184) );
  NOR2_X1 NOR2_1954( .ZN(N5250), .A1(N5184), .A2(N675) );
  NOR2_X1 NOR2_1955( .ZN(N5251), .A1(N5013), .A2(N5184) );
  NOR2_X1 NOR2_1956( .ZN(N5254), .A1(N5127), .A2(N5188) );
  NOR2_X1 NOR2_1957( .ZN(N5255), .A1(N5188), .A2(N723) );
  NOR2_X1 NOR2_1958( .ZN(N5256), .A1(N5017), .A2(N5188) );
  NOR2_X1 NOR2_1959( .ZN(N5259), .A1(N5192), .A2(N5193) );
  NOR2_X1 NOR2_1960( .ZN(N5262), .A1(N5197), .A2(N5194) );
  NOR2_X1 NOR2_1961( .ZN(N5266), .A1(N5139), .A2(N5200) );
  NOR2_X1 NOR2_1962( .ZN(N5267), .A1(N5200), .A2(N5136) );
  NOR2_X1 NOR2_1963( .ZN(N5268), .A1(N5204), .A2(N5205) );
  NOR2_X1 NOR2_1964( .ZN(N5271), .A1(N5206), .A2(N918) );
  NOR2_X1 NOR2_1965( .ZN(N5275), .A1(N5148), .A2(N5209) );
  NOR2_X1 NOR2_1966( .ZN(N5276), .A1(N5209), .A2(N966) );
  NOR2_X2 NOR2_1967( .ZN(N5277), .A1(N5038), .A2(N5209) );
  NOR2_X2 NOR2_1968( .ZN(N5280), .A1(N5213), .A2(N5214) );
  NOR2_X2 NOR2_1969( .ZN(N5283), .A1(N5218), .A2(N5215) );
  NOR2_X2 NOR2_1970( .ZN(N5287), .A1(N5160), .A2(N5221) );
  NOR2_X2 NOR2_1971( .ZN(N5288), .A1(N5221), .A2(N5157) );
  NOR2_X2 NOR2_1972( .ZN(N5289), .A1(N5225), .A2(N5226) );
  NOR2_X2 NOR2_1973( .ZN(N5292), .A1(N5227), .A2(N1161) );
  NOR2_X2 NOR2_1974( .ZN(N5296), .A1(N5169), .A2(N5230) );
  NOR2_X2 NOR2_1975( .ZN(N5297), .A1(N5230), .A2(N1209) );
  NOR2_X1 NOR2_1976( .ZN(N5298), .A1(N5059), .A2(N5230) );
  NOR2_X1 NOR2_1977( .ZN(N5301), .A1(N5234), .A2(N5235) );
  NOR2_X1 NOR2_1978( .ZN(N5304), .A1(N1305), .A2(N5236) );
  NOR2_X1 NOR2_1979( .ZN(N5308), .A1(N5239), .A2(N5240) );
  NOR2_X1 NOR2_1980( .ZN(N5309), .A1(N5244), .A2(N5245) );
  NOR2_X1 NOR2_1981( .ZN(N5312), .A1(N5249), .A2(N5250) );
  NOR2_X1 NOR2_1982( .ZN(N5315), .A1(N5254), .A2(N5255) );
  NOR2_X1 NOR2_1983( .ZN(N5318), .A1(N5259), .A2(N5256) );
  NOR2_X1 NOR2_1984( .ZN(N5322), .A1(N5197), .A2(N5262) );
  NOR2_X1 NOR2_1985( .ZN(N5323), .A1(N5262), .A2(N5194) );
  NOR2_X1 NOR2_1986( .ZN(N5324), .A1(N5266), .A2(N5267) );
  NOR2_X1 NOR2_1987( .ZN(N5327), .A1(N5268), .A2(N870) );
  NOR2_X1 NOR2_1988( .ZN(N5331), .A1(N5206), .A2(N5271) );
  NOR2_X1 NOR2_1989( .ZN(N5332), .A1(N5271), .A2(N918) );
  NOR2_X1 NOR2_1990( .ZN(N5333), .A1(N5088), .A2(N5271) );
  NOR2_X1 NOR2_1991( .ZN(N5336), .A1(N5275), .A2(N5276) );
  NOR2_X1 NOR2_1992( .ZN(N5339), .A1(N5280), .A2(N5277) );
  NOR2_X1 NOR2_1993( .ZN(N5343), .A1(N5218), .A2(N5283) );
  NOR2_X1 NOR2_1994( .ZN(N5344), .A1(N5283), .A2(N5215) );
  NOR2_X1 NOR2_1995( .ZN(N5345), .A1(N5287), .A2(N5288) );
  NOR2_X1 NOR2_1996( .ZN(N5348), .A1(N5289), .A2(N1113) );
  NOR2_X1 NOR2_1997( .ZN(N5352), .A1(N5227), .A2(N5292) );
  NOR2_X1 NOR2_1998( .ZN(N5353), .A1(N5292), .A2(N1161) );
  NOR2_X1 NOR2_1999( .ZN(N5354), .A1(N5109), .A2(N5292) );
  NOR2_X1 NOR2_2000( .ZN(N5357), .A1(N5296), .A2(N5297) );
  NOR2_X1 NOR2_2001( .ZN(N5360), .A1(N5301), .A2(N5298) );
  NOR2_X1 NOR2_2002( .ZN(N5364), .A1(N1305), .A2(N5304) );
  NOR2_X1 NOR2_2003( .ZN(N5365), .A1(N5304), .A2(N5236) );
  NOR2_X1 NOR2_2004( .ZN(N5366), .A1(N5309), .A2(N5241) );
  NOR2_X1 NOR2_2005( .ZN(N5370), .A1(N5312), .A2(N5246) );
  NOR2_X1 NOR2_2006( .ZN(N5374), .A1(N5315), .A2(N5251) );
  NOR2_X1 NOR2_2007( .ZN(N5378), .A1(N5259), .A2(N5318) );
  NOR2_X1 NOR2_2008( .ZN(N5379), .A1(N5318), .A2(N5256) );
  NOR2_X1 NOR2_2009( .ZN(N5380), .A1(N5322), .A2(N5323) );
  NOR2_X1 NOR2_2010( .ZN(N5383), .A1(N5324), .A2(N822) );
  NOR2_X1 NOR2_2011( .ZN(N5387), .A1(N5268), .A2(N5327) );
  NOR2_X1 NOR2_2012( .ZN(N5388), .A1(N5327), .A2(N870) );
  NOR2_X1 NOR2_2013( .ZN(N5389), .A1(N5142), .A2(N5327) );
  NOR2_X1 NOR2_2014( .ZN(N5392), .A1(N5331), .A2(N5332) );
  NOR2_X1 NOR2_2015( .ZN(N5395), .A1(N5336), .A2(N5333) );
  NOR2_X1 NOR2_2016( .ZN(N5399), .A1(N5280), .A2(N5339) );
  NOR2_X1 NOR2_2017( .ZN(N5400), .A1(N5339), .A2(N5277) );
  NOR2_X1 NOR2_2018( .ZN(N5401), .A1(N5343), .A2(N5344) );
  NOR2_X1 NOR2_2019( .ZN(N5404), .A1(N5345), .A2(N1065) );
  NOR2_X1 NOR2_2020( .ZN(N5408), .A1(N5289), .A2(N5348) );
  NOR2_X1 NOR2_2021( .ZN(N5409), .A1(N5348), .A2(N1113) );
  NOR2_X1 NOR2_2022( .ZN(N5410), .A1(N5163), .A2(N5348) );
  NOR2_X1 NOR2_2023( .ZN(N5413), .A1(N5352), .A2(N5353) );
  NOR2_X1 NOR2_2024( .ZN(N5416), .A1(N5357), .A2(N5354) );
  NOR2_X1 NOR2_2025( .ZN(N5420), .A1(N5301), .A2(N5360) );
  NOR2_X1 NOR2_2026( .ZN(N5421), .A1(N5360), .A2(N5298) );
  NOR2_X1 NOR2_2027( .ZN(N5422), .A1(N5364), .A2(N5365) );
  NOR2_X1 NOR2_2028( .ZN(N5425), .A1(N5309), .A2(N5366) );
  NOR2_X1 NOR2_2029( .ZN(N5426), .A1(N5366), .A2(N5241) );
  NOR2_X1 NOR2_2030( .ZN(N5427), .A1(N5312), .A2(N5370) );
  NOR2_X1 NOR2_2031( .ZN(N5428), .A1(N5370), .A2(N5246) );
  NOR2_X1 NOR2_2032( .ZN(N5429), .A1(N5315), .A2(N5374) );
  NOR2_X1 NOR2_2033( .ZN(N5430), .A1(N5374), .A2(N5251) );
  NOR2_X1 NOR2_2034( .ZN(N5431), .A1(N5378), .A2(N5379) );
  NOR2_X1 NOR2_2035( .ZN(N5434), .A1(N5380), .A2(N774) );
  NOR2_X1 NOR2_2036( .ZN(N5438), .A1(N5324), .A2(N5383) );
  NOR2_X1 NOR2_2037( .ZN(N5439), .A1(N5383), .A2(N822) );
  NOR2_X1 NOR2_2038( .ZN(N5440), .A1(N5200), .A2(N5383) );
  NOR2_X1 NOR2_2039( .ZN(N5443), .A1(N5387), .A2(N5388) );
  NOR2_X1 NOR2_2040( .ZN(N5446), .A1(N5392), .A2(N5389) );
  NOR2_X1 NOR2_2041( .ZN(N5450), .A1(N5336), .A2(N5395) );
  NOR2_X1 NOR2_2042( .ZN(N5451), .A1(N5395), .A2(N5333) );
  NOR2_X1 NOR2_2043( .ZN(N5452), .A1(N5399), .A2(N5400) );
  NOR2_X1 NOR2_2044( .ZN(N5455), .A1(N5401), .A2(N1017) );
  NOR2_X1 NOR2_2045( .ZN(N5459), .A1(N5345), .A2(N5404) );
  NOR2_X1 NOR2_2046( .ZN(N5460), .A1(N5404), .A2(N1065) );
  NOR2_X1 NOR2_2047( .ZN(N5461), .A1(N5221), .A2(N5404) );
  NOR2_X1 NOR2_2048( .ZN(N5464), .A1(N5408), .A2(N5409) );
  NOR2_X1 NOR2_2049( .ZN(N5467), .A1(N5413), .A2(N5410) );
  NOR2_X1 NOR2_2050( .ZN(N5471), .A1(N5357), .A2(N5416) );
  NOR2_X1 NOR2_2051( .ZN(N5472), .A1(N5416), .A2(N5354) );
  NOR2_X1 NOR2_2052( .ZN(N5473), .A1(N5420), .A2(N5421) );
  NOR2_X1 NOR2_2053( .ZN(N5476), .A1(N5422), .A2(N1260) );
  NOR2_X1 NOR2_2054( .ZN(N5480), .A1(N5425), .A2(N5426) );
  NOR2_X1 NOR2_2055( .ZN(N5483), .A1(N5427), .A2(N5428) );
  NOR2_X1 NOR2_2056( .ZN(N5486), .A1(N5429), .A2(N5430) );
  NOR2_X1 NOR2_2057( .ZN(N5489), .A1(N5431), .A2(N726) );
  NOR2_X1 NOR2_2058( .ZN(N5493), .A1(N5380), .A2(N5434) );
  NOR2_X1 NOR2_2059( .ZN(N5494), .A1(N5434), .A2(N774) );
  NOR2_X1 NOR2_2060( .ZN(N5495), .A1(N5262), .A2(N5434) );
  NOR2_X1 NOR2_2061( .ZN(N5498), .A1(N5438), .A2(N5439) );
  NOR2_X1 NOR2_2062( .ZN(N5501), .A1(N5443), .A2(N5440) );
  NOR2_X1 NOR2_2063( .ZN(N5505), .A1(N5392), .A2(N5446) );
  NOR2_X1 NOR2_2064( .ZN(N5506), .A1(N5446), .A2(N5389) );
  NOR2_X1 NOR2_2065( .ZN(N5507), .A1(N5450), .A2(N5451) );
  NOR2_X1 NOR2_2066( .ZN(N5510), .A1(N5452), .A2(N969) );
  NOR2_X1 NOR2_2067( .ZN(N5514), .A1(N5401), .A2(N5455) );
  NOR2_X1 NOR2_2068( .ZN(N5515), .A1(N5455), .A2(N1017) );
  NOR2_X1 NOR2_2069( .ZN(N5516), .A1(N5283), .A2(N5455) );
  NOR2_X1 NOR2_2070( .ZN(N5519), .A1(N5459), .A2(N5460) );
  NOR2_X1 NOR2_2071( .ZN(N5522), .A1(N5464), .A2(N5461) );
  NOR2_X1 NOR2_2072( .ZN(N5526), .A1(N5413), .A2(N5467) );
  NOR2_X1 NOR2_2073( .ZN(N5527), .A1(N5467), .A2(N5410) );
  NOR2_X1 NOR2_2074( .ZN(N5528), .A1(N5471), .A2(N5472) );
  NOR2_X1 NOR2_2075( .ZN(N5531), .A1(N5473), .A2(N1212) );
  NOR2_X1 NOR2_2076( .ZN(N5535), .A1(N5422), .A2(N5476) );
  NOR2_X1 NOR2_2077( .ZN(N5536), .A1(N5476), .A2(N1260) );
  NOR2_X1 NOR2_2078( .ZN(N5537), .A1(N5304), .A2(N5476) );
  NOR2_X1 NOR2_2079( .ZN(N5540), .A1(N5480), .A2(N582) );
  NOR2_X1 NOR2_2080( .ZN(N5544), .A1(N5483), .A2(N630) );
  NOR2_X1 NOR2_2081( .ZN(N5548), .A1(N5486), .A2(N678) );
  NOR2_X1 NOR2_2082( .ZN(N5552), .A1(N5431), .A2(N5489) );
  NOR2_X1 NOR2_2083( .ZN(N5553), .A1(N5489), .A2(N726) );
  NOR2_X1 NOR2_2084( .ZN(N5554), .A1(N5318), .A2(N5489) );
  NOR2_X1 NOR2_2085( .ZN(N5557), .A1(N5493), .A2(N5494) );
  NOR2_X1 NOR2_2086( .ZN(N5560), .A1(N5498), .A2(N5495) );
  NOR2_X1 NOR2_2087( .ZN(N5564), .A1(N5443), .A2(N5501) );
  NOR2_X1 NOR2_2088( .ZN(N5565), .A1(N5501), .A2(N5440) );
  NOR2_X1 NOR2_2089( .ZN(N5566), .A1(N5505), .A2(N5506) );
  NOR2_X1 NOR2_2090( .ZN(N5569), .A1(N5507), .A2(N921) );
  NOR2_X1 NOR2_2091( .ZN(N5573), .A1(N5452), .A2(N5510) );
  NOR2_X1 NOR2_2092( .ZN(N5574), .A1(N5510), .A2(N969) );
  NOR2_X1 NOR2_2093( .ZN(N5575), .A1(N5339), .A2(N5510) );
  NOR2_X1 NOR2_2094( .ZN(N5578), .A1(N5514), .A2(N5515) );
  NOR2_X1 NOR2_2095( .ZN(N5581), .A1(N5519), .A2(N5516) );
  NOR2_X1 NOR2_2096( .ZN(N5585), .A1(N5464), .A2(N5522) );
  NOR2_X1 NOR2_2097( .ZN(N5586), .A1(N5522), .A2(N5461) );
  NOR2_X1 NOR2_2098( .ZN(N5587), .A1(N5526), .A2(N5527) );
  NOR2_X1 NOR2_2099( .ZN(N5590), .A1(N5528), .A2(N1164) );
  NOR2_X1 NOR2_2100( .ZN(N5594), .A1(N5473), .A2(N5531) );
  NOR2_X1 NOR2_2101( .ZN(N5595), .A1(N5531), .A2(N1212) );
  NOR2_X1 NOR2_2102( .ZN(N5596), .A1(N5360), .A2(N5531) );
  NOR2_X1 NOR2_2103( .ZN(N5599), .A1(N5535), .A2(N5536) );
  NOR2_X1 NOR2_2104( .ZN(N5602), .A1(N1308), .A2(N5537) );
  NOR2_X1 NOR2_2105( .ZN(N5606), .A1(N5480), .A2(N5540) );
  NOR2_X1 NOR2_2106( .ZN(N5607), .A1(N5540), .A2(N582) );
  NOR2_X1 NOR2_2107( .ZN(N5608), .A1(N5366), .A2(N5540) );
  NOR2_X1 NOR2_2108( .ZN(N5611), .A1(N5483), .A2(N5544) );
  NOR2_X1 NOR2_2109( .ZN(N5612), .A1(N5544), .A2(N630) );
  NOR2_X1 NOR2_2110( .ZN(N5613), .A1(N5370), .A2(N5544) );
  NOR2_X1 NOR2_2111( .ZN(N5616), .A1(N5486), .A2(N5548) );
  NOR2_X1 NOR2_2112( .ZN(N5617), .A1(N5548), .A2(N678) );
  NOR2_X1 NOR2_2113( .ZN(N5618), .A1(N5374), .A2(N5548) );
  NOR2_X1 NOR2_2114( .ZN(N5621), .A1(N5552), .A2(N5553) );
  NOR2_X1 NOR2_2115( .ZN(N5624), .A1(N5557), .A2(N5554) );
  NOR2_X1 NOR2_2116( .ZN(N5628), .A1(N5498), .A2(N5560) );
  NOR2_X1 NOR2_2117( .ZN(N5629), .A1(N5560), .A2(N5495) );
  NOR2_X1 NOR2_2118( .ZN(N5630), .A1(N5564), .A2(N5565) );
  NOR2_X1 NOR2_2119( .ZN(N5633), .A1(N5566), .A2(N873) );
  NOR2_X1 NOR2_2120( .ZN(N5637), .A1(N5507), .A2(N5569) );
  NOR2_X1 NOR2_2121( .ZN(N5638), .A1(N5569), .A2(N921) );
  NOR2_X1 NOR2_2122( .ZN(N5639), .A1(N5395), .A2(N5569) );
  NOR2_X1 NOR2_2123( .ZN(N5642), .A1(N5573), .A2(N5574) );
  NOR2_X1 NOR2_2124( .ZN(N5645), .A1(N5578), .A2(N5575) );
  NOR2_X1 NOR2_2125( .ZN(N5649), .A1(N5519), .A2(N5581) );
  NOR2_X1 NOR2_2126( .ZN(N5650), .A1(N5581), .A2(N5516) );
  NOR2_X1 NOR2_2127( .ZN(N5651), .A1(N5585), .A2(N5586) );
  NOR2_X1 NOR2_2128( .ZN(N5654), .A1(N5587), .A2(N1116) );
  NOR2_X1 NOR2_2129( .ZN(N5658), .A1(N5528), .A2(N5590) );
  NOR2_X1 NOR2_2130( .ZN(N5659), .A1(N5590), .A2(N1164) );
  NOR2_X1 NOR2_2131( .ZN(N5660), .A1(N5416), .A2(N5590) );
  NOR2_X1 NOR2_2132( .ZN(N5663), .A1(N5594), .A2(N5595) );
  NOR2_X1 NOR2_2133( .ZN(N5666), .A1(N5599), .A2(N5596) );
  NOR2_X1 NOR2_2134( .ZN(N5670), .A1(N1308), .A2(N5602) );
  NOR2_X1 NOR2_2135( .ZN(N5671), .A1(N5602), .A2(N5537) );
  NOR2_X1 NOR2_2136( .ZN(N5672), .A1(N5606), .A2(N5607) );
  NOR2_X1 NOR2_2137( .ZN(N5673), .A1(N5611), .A2(N5612) );
  NOR2_X1 NOR2_2138( .ZN(N5676), .A1(N5616), .A2(N5617) );
  NOR2_X1 NOR2_2139( .ZN(N5679), .A1(N5621), .A2(N5618) );
  NOR2_X1 NOR2_2140( .ZN(N5683), .A1(N5557), .A2(N5624) );
  NOR2_X1 NOR2_2141( .ZN(N5684), .A1(N5624), .A2(N5554) );
  NOR2_X1 NOR2_2142( .ZN(N5685), .A1(N5628), .A2(N5629) );
  NOR2_X1 NOR2_2143( .ZN(N5688), .A1(N5630), .A2(N825) );
  NOR2_X1 NOR2_2144( .ZN(N5692), .A1(N5566), .A2(N5633) );
  NOR2_X1 NOR2_2145( .ZN(N5693), .A1(N5633), .A2(N873) );
  NOR2_X1 NOR2_2146( .ZN(N5694), .A1(N5446), .A2(N5633) );
  NOR2_X1 NOR2_2147( .ZN(N5697), .A1(N5637), .A2(N5638) );
  NOR2_X1 NOR2_2148( .ZN(N5700), .A1(N5642), .A2(N5639) );
  NOR2_X1 NOR2_2149( .ZN(N5704), .A1(N5578), .A2(N5645) );
  NOR2_X1 NOR2_2150( .ZN(N5705), .A1(N5645), .A2(N5575) );
  NOR2_X1 NOR2_2151( .ZN(N5706), .A1(N5649), .A2(N5650) );
  NOR2_X1 NOR2_2152( .ZN(N5709), .A1(N5651), .A2(N1068) );
  NOR2_X1 NOR2_2153( .ZN(N5713), .A1(N5587), .A2(N5654) );
  NOR2_X1 NOR2_2154( .ZN(N5714), .A1(N5654), .A2(N1116) );
  NOR2_X1 NOR2_2155( .ZN(N5715), .A1(N5467), .A2(N5654) );
  NOR2_X1 NOR2_2156( .ZN(N5718), .A1(N5658), .A2(N5659) );
  NOR2_X1 NOR2_2157( .ZN(N5721), .A1(N5663), .A2(N5660) );
  NOR2_X1 NOR2_2158( .ZN(N5725), .A1(N5599), .A2(N5666) );
  NOR2_X1 NOR2_2159( .ZN(N5726), .A1(N5666), .A2(N5596) );
  NOR2_X1 NOR2_2160( .ZN(N5727), .A1(N5670), .A2(N5671) );
  NOR2_X1 NOR2_2161( .ZN(N5730), .A1(N5673), .A2(N5608) );
  NOR2_X1 NOR2_2162( .ZN(N5734), .A1(N5676), .A2(N5613) );
  NOR2_X1 NOR2_2163( .ZN(N5738), .A1(N5621), .A2(N5679) );
  NOR2_X1 NOR2_2164( .ZN(N5739), .A1(N5679), .A2(N5618) );
  NOR2_X1 NOR2_2165( .ZN(N5740), .A1(N5683), .A2(N5684) );
  NOR2_X1 NOR2_2166( .ZN(N5743), .A1(N5685), .A2(N777) );
  NOR2_X1 NOR2_2167( .ZN(N5747), .A1(N5630), .A2(N5688) );
  NOR2_X1 NOR2_2168( .ZN(N5748), .A1(N5688), .A2(N825) );
  NOR2_X1 NOR2_2169( .ZN(N5749), .A1(N5501), .A2(N5688) );
  NOR2_X1 NOR2_2170( .ZN(N5752), .A1(N5692), .A2(N5693) );
  NOR2_X1 NOR2_2171( .ZN(N5755), .A1(N5697), .A2(N5694) );
  NOR2_X1 NOR2_2172( .ZN(N5759), .A1(N5642), .A2(N5700) );
  NOR2_X1 NOR2_2173( .ZN(N5760), .A1(N5700), .A2(N5639) );
  NOR2_X1 NOR2_2174( .ZN(N5761), .A1(N5704), .A2(N5705) );
  NOR2_X1 NOR2_2175( .ZN(N5764), .A1(N5706), .A2(N1020) );
  NOR2_X1 NOR2_2176( .ZN(N5768), .A1(N5651), .A2(N5709) );
  NOR2_X1 NOR2_2177( .ZN(N5769), .A1(N5709), .A2(N1068) );
  NOR2_X1 NOR2_2178( .ZN(N5770), .A1(N5522), .A2(N5709) );
  NOR2_X1 NOR2_2179( .ZN(N5773), .A1(N5713), .A2(N5714) );
  NOR2_X1 NOR2_2180( .ZN(N5776), .A1(N5718), .A2(N5715) );
  NOR2_X1 NOR2_2181( .ZN(N5780), .A1(N5663), .A2(N5721) );
  NOR2_X1 NOR2_2182( .ZN(N5781), .A1(N5721), .A2(N5660) );
  NOR2_X1 NOR2_2183( .ZN(N5782), .A1(N5725), .A2(N5726) );
  NOR2_X1 NOR2_2184( .ZN(N5785), .A1(N5673), .A2(N5730) );
  NOR2_X1 NOR2_2185( .ZN(N5786), .A1(N5730), .A2(N5608) );
  NOR2_X1 NOR2_2186( .ZN(N5787), .A1(N5676), .A2(N5734) );
  NOR2_X1 NOR2_2187( .ZN(N5788), .A1(N5734), .A2(N5613) );
  NOR2_X1 NOR2_2188( .ZN(N5789), .A1(N5738), .A2(N5739) );
  NOR2_X1 NOR2_2189( .ZN(N5792), .A1(N5740), .A2(N729) );
  NOR2_X1 NOR2_2190( .ZN(N5796), .A1(N5685), .A2(N5743) );
  NOR2_X1 NOR2_2191( .ZN(N5797), .A1(N5743), .A2(N777) );
  NOR2_X1 NOR2_2192( .ZN(N5798), .A1(N5560), .A2(N5743) );
  NOR2_X1 NOR2_2193( .ZN(N5801), .A1(N5747), .A2(N5748) );
  NOR2_X1 NOR2_2194( .ZN(N5804), .A1(N5752), .A2(N5749) );
  NOR2_X1 NOR2_2195( .ZN(N5808), .A1(N5697), .A2(N5755) );
  NOR2_X1 NOR2_2196( .ZN(N5809), .A1(N5755), .A2(N5694) );
  NOR2_X1 NOR2_2197( .ZN(N5810), .A1(N5759), .A2(N5760) );
  NOR2_X1 NOR2_2198( .ZN(N5813), .A1(N5761), .A2(N972) );
  NOR2_X1 NOR2_2199( .ZN(N5817), .A1(N5706), .A2(N5764) );
  NOR2_X1 NOR2_2200( .ZN(N5818), .A1(N5764), .A2(N1020) );
  NOR2_X1 NOR2_2201( .ZN(N5819), .A1(N5581), .A2(N5764) );
  NOR2_X1 NOR2_2202( .ZN(N5822), .A1(N5768), .A2(N5769) );
  NOR2_X1 NOR2_2203( .ZN(N5825), .A1(N5773), .A2(N5770) );
  NOR2_X1 NOR2_2204( .ZN(N5829), .A1(N5718), .A2(N5776) );
  NOR2_X1 NOR2_2205( .ZN(N5830), .A1(N5776), .A2(N5715) );
  NOR2_X1 NOR2_2206( .ZN(N5831), .A1(N5780), .A2(N5781) );
  NOR2_X1 NOR2_2207( .ZN(N5834), .A1(N5785), .A2(N5786) );
  NOR2_X1 NOR2_2208( .ZN(N5837), .A1(N5787), .A2(N5788) );
  NOR2_X1 NOR2_2209( .ZN(N5840), .A1(N5789), .A2(N681) );
  NOR2_X1 NOR2_2210( .ZN(N5844), .A1(N5740), .A2(N5792) );
  NOR2_X1 NOR2_2211( .ZN(N5845), .A1(N5792), .A2(N729) );
  NOR2_X1 NOR2_2212( .ZN(N5846), .A1(N5624), .A2(N5792) );
  NOR2_X1 NOR2_2213( .ZN(N5849), .A1(N5796), .A2(N5797) );
  NOR2_X1 NOR2_2214( .ZN(N5852), .A1(N5801), .A2(N5798) );
  NOR2_X1 NOR2_2215( .ZN(N5856), .A1(N5752), .A2(N5804) );
  NOR2_X1 NOR2_2216( .ZN(N5857), .A1(N5804), .A2(N5749) );
  NOR2_X1 NOR2_2217( .ZN(N5858), .A1(N5808), .A2(N5809) );
  NOR2_X1 NOR2_2218( .ZN(N5861), .A1(N5810), .A2(N924) );
  NOR2_X1 NOR2_2219( .ZN(N5865), .A1(N5761), .A2(N5813) );
  NOR2_X1 NOR2_2220( .ZN(N5866), .A1(N5813), .A2(N972) );
  NOR2_X1 NOR2_2221( .ZN(N5867), .A1(N5645), .A2(N5813) );
  NOR2_X1 NOR2_2222( .ZN(N5870), .A1(N5817), .A2(N5818) );
  NOR2_X1 NOR2_2223( .ZN(N5873), .A1(N5822), .A2(N5819) );
  NOR2_X1 NOR2_2224( .ZN(N5877), .A1(N5773), .A2(N5825) );
  NOR2_X1 NOR2_2225( .ZN(N5878), .A1(N5825), .A2(N5770) );
  NOR2_X1 NOR2_2226( .ZN(N5879), .A1(N5829), .A2(N5830) );
  NOR2_X1 NOR2_2227( .ZN(N5882), .A1(N5834), .A2(N585) );
  NOR2_X1 NOR2_2228( .ZN(N5886), .A1(N5837), .A2(N633) );
  NOR2_X1 NOR2_2229( .ZN(N5890), .A1(N5789), .A2(N5840) );
  NOR2_X1 NOR2_2230( .ZN(N5891), .A1(N5840), .A2(N681) );
  NOR2_X1 NOR2_2231( .ZN(N5892), .A1(N5679), .A2(N5840) );
  NOR2_X1 NOR2_2232( .ZN(N5895), .A1(N5844), .A2(N5845) );
  NOR2_X1 NOR2_2233( .ZN(N5898), .A1(N5849), .A2(N5846) );
  NOR2_X1 NOR2_2234( .ZN(N5902), .A1(N5801), .A2(N5852) );
  NOR2_X1 NOR2_2235( .ZN(N5903), .A1(N5852), .A2(N5798) );
  NOR2_X1 NOR2_2236( .ZN(N5904), .A1(N5856), .A2(N5857) );
  NOR2_X1 NOR2_2237( .ZN(N5907), .A1(N5858), .A2(N876) );
  NOR2_X1 NOR2_2238( .ZN(N5911), .A1(N5810), .A2(N5861) );
  NOR2_X1 NOR2_2239( .ZN(N5912), .A1(N5861), .A2(N924) );
  NOR2_X1 NOR2_2240( .ZN(N5913), .A1(N5700), .A2(N5861) );
  NOR2_X2 NOR2_2241( .ZN(N5916), .A1(N5865), .A2(N5866) );
  NOR2_X2 NOR2_2242( .ZN(N5919), .A1(N5870), .A2(N5867) );
  NOR2_X2 NOR2_2243( .ZN(N5923), .A1(N5822), .A2(N5873) );
  NOR2_X2 NOR2_2244( .ZN(N5924), .A1(N5873), .A2(N5819) );
  NOR2_X2 NOR2_2245( .ZN(N5925), .A1(N5877), .A2(N5878) );
  NOR2_X2 NOR2_2246( .ZN(N5928), .A1(N5834), .A2(N5882) );
  NOR2_X2 NOR2_2247( .ZN(N5929), .A1(N5882), .A2(N585) );
  NOR2_X2 NOR2_2248( .ZN(N5930), .A1(N5730), .A2(N5882) );
  NOR2_X2 NOR2_2249( .ZN(N5933), .A1(N5837), .A2(N5886) );
  NOR2_X1 NOR2_2250( .ZN(N5934), .A1(N5886), .A2(N633) );
  NOR2_X1 NOR2_2251( .ZN(N5935), .A1(N5734), .A2(N5886) );
  NOR2_X1 NOR2_2252( .ZN(N5938), .A1(N5890), .A2(N5891) );
  NOR2_X1 NOR2_2253( .ZN(N5941), .A1(N5895), .A2(N5892) );
  NOR2_X1 NOR2_2254( .ZN(N5945), .A1(N5849), .A2(N5898) );
  NOR2_X1 NOR2_2255( .ZN(N5946), .A1(N5898), .A2(N5846) );
  NOR2_X1 NOR2_2256( .ZN(N5947), .A1(N5902), .A2(N5903) );
  NOR2_X1 NOR2_2257( .ZN(N5950), .A1(N5904), .A2(N828) );
  NOR2_X1 NOR2_2258( .ZN(N5954), .A1(N5858), .A2(N5907) );
  NOR2_X1 NOR2_2259( .ZN(N5955), .A1(N5907), .A2(N876) );
  NOR2_X1 NOR2_2260( .ZN(N5956), .A1(N5755), .A2(N5907) );
  NOR2_X1 NOR2_2261( .ZN(N5959), .A1(N5911), .A2(N5912) );
  NOR2_X1 NOR2_2262( .ZN(N5962), .A1(N5916), .A2(N5913) );
  NOR2_X1 NOR2_2263( .ZN(N5966), .A1(N5870), .A2(N5919) );
  NOR2_X1 NOR2_2264( .ZN(N5967), .A1(N5919), .A2(N5867) );
  NOR2_X1 NOR2_2265( .ZN(N5968), .A1(N5923), .A2(N5924) );
  NOR2_X1 NOR2_2266( .ZN(N5971), .A1(N5928), .A2(N5929) );
  NOR2_X1 NOR2_2267( .ZN(N5972), .A1(N5933), .A2(N5934) );
  NOR2_X1 NOR2_2268( .ZN(N5975), .A1(N5938), .A2(N5935) );
  NOR2_X1 NOR2_2269( .ZN(N5979), .A1(N5895), .A2(N5941) );
  NOR2_X1 NOR2_2270( .ZN(N5980), .A1(N5941), .A2(N5892) );
  NOR2_X1 NOR2_2271( .ZN(N5981), .A1(N5945), .A2(N5946) );
  NOR2_X1 NOR2_2272( .ZN(N5984), .A1(N5947), .A2(N780) );
  NOR2_X1 NOR2_2273( .ZN(N5988), .A1(N5904), .A2(N5950) );
  NOR2_X1 NOR2_2274( .ZN(N5989), .A1(N5950), .A2(N828) );
  NOR2_X1 NOR2_2275( .ZN(N5990), .A1(N5804), .A2(N5950) );
  NOR2_X1 NOR2_2276( .ZN(N5993), .A1(N5954), .A2(N5955) );
  NOR2_X1 NOR2_2277( .ZN(N5996), .A1(N5959), .A2(N5956) );
  NOR2_X1 NOR2_2278( .ZN(N6000), .A1(N5916), .A2(N5962) );
  NOR2_X1 NOR2_2279( .ZN(N6001), .A1(N5962), .A2(N5913) );
  NOR2_X1 NOR2_2280( .ZN(N6002), .A1(N5966), .A2(N5967) );
  NOR2_X1 NOR2_2281( .ZN(N6005), .A1(N5972), .A2(N5930) );
  NOR2_X1 NOR2_2282( .ZN(N6009), .A1(N5938), .A2(N5975) );
  NOR2_X1 NOR2_2283( .ZN(N6010), .A1(N5975), .A2(N5935) );
  NOR2_X1 NOR2_2284( .ZN(N6011), .A1(N5979), .A2(N5980) );
  NOR2_X1 NOR2_2285( .ZN(N6014), .A1(N5981), .A2(N732) );
  NOR2_X1 NOR2_2286( .ZN(N6018), .A1(N5947), .A2(N5984) );
  NOR2_X1 NOR2_2287( .ZN(N6019), .A1(N5984), .A2(N780) );
  NOR2_X1 NOR2_2288( .ZN(N6020), .A1(N5852), .A2(N5984) );
  NOR2_X1 NOR2_2289( .ZN(N6023), .A1(N5988), .A2(N5989) );
  NOR2_X1 NOR2_2290( .ZN(N6026), .A1(N5993), .A2(N5990) );
  NOR2_X1 NOR2_2291( .ZN(N6030), .A1(N5959), .A2(N5996) );
  NOR2_X1 NOR2_2292( .ZN(N6031), .A1(N5996), .A2(N5956) );
  NOR2_X1 NOR2_2293( .ZN(N6032), .A1(N6000), .A2(N6001) );
  NOR2_X1 NOR2_2294( .ZN(N6035), .A1(N5972), .A2(N6005) );
  NOR2_X1 NOR2_2295( .ZN(N6036), .A1(N6005), .A2(N5930) );
  NOR2_X1 NOR2_2296( .ZN(N6037), .A1(N6009), .A2(N6010) );
  NOR2_X1 NOR2_2297( .ZN(N6040), .A1(N6011), .A2(N684) );
  NOR2_X1 NOR2_2298( .ZN(N6044), .A1(N5981), .A2(N6014) );
  NOR2_X1 NOR2_2299( .ZN(N6045), .A1(N6014), .A2(N732) );
  NOR2_X1 NOR2_2300( .ZN(N6046), .A1(N5898), .A2(N6014) );
  NOR2_X1 NOR2_2301( .ZN(N6049), .A1(N6018), .A2(N6019) );
  NOR2_X1 NOR2_2302( .ZN(N6052), .A1(N6023), .A2(N6020) );
  NOR2_X1 NOR2_2303( .ZN(N6056), .A1(N5993), .A2(N6026) );
  NOR2_X1 NOR2_2304( .ZN(N6057), .A1(N6026), .A2(N5990) );
  NOR2_X1 NOR2_2305( .ZN(N6058), .A1(N6030), .A2(N6031) );
  NOR2_X1 NOR2_2306( .ZN(N6061), .A1(N6035), .A2(N6036) );
  NOR2_X1 NOR2_2307( .ZN(N6064), .A1(N6037), .A2(N636) );
  NOR2_X1 NOR2_2308( .ZN(N6068), .A1(N6011), .A2(N6040) );
  NOR2_X1 NOR2_2309( .ZN(N6069), .A1(N6040), .A2(N684) );
  NOR2_X1 NOR2_2310( .ZN(N6070), .A1(N5941), .A2(N6040) );
  NOR2_X1 NOR2_2311( .ZN(N6073), .A1(N6044), .A2(N6045) );
  NOR2_X1 NOR2_2312( .ZN(N6076), .A1(N6049), .A2(N6046) );
  NOR2_X1 NOR2_2313( .ZN(N6080), .A1(N6023), .A2(N6052) );
  NOR2_X1 NOR2_2314( .ZN(N6081), .A1(N6052), .A2(N6020) );
  NOR2_X1 NOR2_2315( .ZN(N6082), .A1(N6056), .A2(N6057) );
  NOR2_X1 NOR2_2316( .ZN(N6085), .A1(N6061), .A2(N588) );
  NOR2_X1 NOR2_2317( .ZN(N6089), .A1(N6037), .A2(N6064) );
  NOR2_X1 NOR2_2318( .ZN(N6090), .A1(N6064), .A2(N636) );
  NOR2_X1 NOR2_2319( .ZN(N6091), .A1(N5975), .A2(N6064) );
  NOR2_X1 NOR2_2320( .ZN(N6094), .A1(N6068), .A2(N6069) );
  NOR2_X1 NOR2_2321( .ZN(N6097), .A1(N6073), .A2(N6070) );
  NOR2_X1 NOR2_2322( .ZN(N6101), .A1(N6049), .A2(N6076) );
  NOR2_X1 NOR2_2323( .ZN(N6102), .A1(N6076), .A2(N6046) );
  NOR2_X1 NOR2_2324( .ZN(N6103), .A1(N6080), .A2(N6081) );
  NOR2_X1 NOR2_2325( .ZN(N6106), .A1(N6061), .A2(N6085) );
  NOR2_X1 NOR2_2326( .ZN(N6107), .A1(N6085), .A2(N588) );
  NOR2_X1 NOR2_2327( .ZN(N6108), .A1(N6005), .A2(N6085) );
  NOR2_X1 NOR2_2328( .ZN(N6111), .A1(N6089), .A2(N6090) );
  NOR2_X1 NOR2_2329( .ZN(N6114), .A1(N6094), .A2(N6091) );
  NOR2_X1 NOR2_2330( .ZN(N6118), .A1(N6073), .A2(N6097) );
  NOR2_X1 NOR2_2331( .ZN(N6119), .A1(N6097), .A2(N6070) );
  NOR2_X1 NOR2_2332( .ZN(N6120), .A1(N6101), .A2(N6102) );
  NOR2_X1 NOR2_2333( .ZN(N6123), .A1(N6106), .A2(N6107) );
  NOR2_X1 NOR2_2334( .ZN(N6124), .A1(N6111), .A2(N6108) );
  NOR2_X1 NOR2_2335( .ZN(N6128), .A1(N6094), .A2(N6114) );
  NOR2_X1 NOR2_2336( .ZN(N6129), .A1(N6114), .A2(N6091) );
  NOR2_X1 NOR2_2337( .ZN(N6130), .A1(N6118), .A2(N6119) );
  NOR2_X1 NOR2_2338( .ZN(N6133), .A1(N6111), .A2(N6124) );
  NOR2_X1 NOR2_2339( .ZN(N6134), .A1(N6124), .A2(N6108) );
  NOR2_X1 NOR2_2340( .ZN(N6135), .A1(N6128), .A2(N6129) );
  NOR2_X1 NOR2_2341( .ZN(N6138), .A1(N6133), .A2(N6134) );
  INV_X1 NOT1_2342( .ZN(N6141), .A(N6138) );
  NOR2_X1 NOR2_2343( .ZN(N6145), .A1(N6138), .A2(N6141) );
  INV_X1 NOT1_2344( .ZN(N6146), .A(N6141) );
  NOR2_X1 NOR2_2345( .ZN(N6147), .A1(N6124), .A2(N6141) );
  NOR2_X1 NOR2_2346( .ZN(N6150), .A1(N6145), .A2(N6146) );
  NOR2_X1 NOR2_2347( .ZN(N6151), .A1(N6135), .A2(N6147) );
  NOR2_X1 NOR2_2348( .ZN(N6155), .A1(N6135), .A2(N6151) );
  NOR2_X1 NOR2_2349( .ZN(N6156), .A1(N6151), .A2(N6147) );
  NOR2_X1 NOR2_2350( .ZN(N6157), .A1(N6114), .A2(N6151) );
  NOR2_X1 NOR2_2351( .ZN(N6160), .A1(N6155), .A2(N6156) );
  NOR2_X1 NOR2_2352( .ZN(N6161), .A1(N6130), .A2(N6157) );
  NOR2_X1 NOR2_2353( .ZN(N6165), .A1(N6130), .A2(N6161) );
  NOR2_X1 NOR2_2354( .ZN(N6166), .A1(N6161), .A2(N6157) );
  NOR2_X1 NOR2_2355( .ZN(N6167), .A1(N6097), .A2(N6161) );
  NOR2_X1 NOR2_2356( .ZN(N6170), .A1(N6165), .A2(N6166) );
  NOR2_X1 NOR2_2357( .ZN(N6171), .A1(N6120), .A2(N6167) );
  NOR2_X1 NOR2_2358( .ZN(N6175), .A1(N6120), .A2(N6171) );
  NOR2_X1 NOR2_2359( .ZN(N6176), .A1(N6171), .A2(N6167) );
  NOR2_X1 NOR2_2360( .ZN(N6177), .A1(N6076), .A2(N6171) );
  NOR2_X1 NOR2_2361( .ZN(N6180), .A1(N6175), .A2(N6176) );
  NOR2_X1 NOR2_2362( .ZN(N6181), .A1(N6103), .A2(N6177) );
  NOR2_X1 NOR2_2363( .ZN(N6185), .A1(N6103), .A2(N6181) );
  NOR2_X1 NOR2_2364( .ZN(N6186), .A1(N6181), .A2(N6177) );
  NOR2_X1 NOR2_2365( .ZN(N6187), .A1(N6052), .A2(N6181) );
  NOR2_X1 NOR2_2366( .ZN(N6190), .A1(N6185), .A2(N6186) );
  NOR2_X1 NOR2_2367( .ZN(N6191), .A1(N6082), .A2(N6187) );
  NOR2_X1 NOR2_2368( .ZN(N6195), .A1(N6082), .A2(N6191) );
  NOR2_X1 NOR2_2369( .ZN(N6196), .A1(N6191), .A2(N6187) );
  NOR2_X1 NOR2_2370( .ZN(N6197), .A1(N6026), .A2(N6191) );
  NOR2_X1 NOR2_2371( .ZN(N6200), .A1(N6195), .A2(N6196) );
  NOR2_X1 NOR2_2372( .ZN(N6201), .A1(N6058), .A2(N6197) );
  NOR2_X1 NOR2_2373( .ZN(N6205), .A1(N6058), .A2(N6201) );
  NOR2_X1 NOR2_2374( .ZN(N6206), .A1(N6201), .A2(N6197) );
  NOR2_X1 NOR2_2375( .ZN(N6207), .A1(N5996), .A2(N6201) );
  NOR2_X1 NOR2_2376( .ZN(N6210), .A1(N6205), .A2(N6206) );
  NOR2_X1 NOR2_2377( .ZN(N6211), .A1(N6032), .A2(N6207) );
  NOR2_X1 NOR2_2378( .ZN(N6215), .A1(N6032), .A2(N6211) );
  NOR2_X1 NOR2_2379( .ZN(N6216), .A1(N6211), .A2(N6207) );
  NOR2_X1 NOR2_2380( .ZN(N6217), .A1(N5962), .A2(N6211) );
  NOR2_X1 NOR2_2381( .ZN(N6220), .A1(N6215), .A2(N6216) );
  NOR2_X1 NOR2_2382( .ZN(N6221), .A1(N6002), .A2(N6217) );
  NOR2_X1 NOR2_2383( .ZN(N6225), .A1(N6002), .A2(N6221) );
  NOR2_X1 NOR2_2384( .ZN(N6226), .A1(N6221), .A2(N6217) );
  NOR2_X1 NOR2_2385( .ZN(N6227), .A1(N5919), .A2(N6221) );
  NOR2_X1 NOR2_2386( .ZN(N6230), .A1(N6225), .A2(N6226) );
  NOR2_X1 NOR2_2387( .ZN(N6231), .A1(N5968), .A2(N6227) );
  NOR2_X1 NOR2_2388( .ZN(N6235), .A1(N5968), .A2(N6231) );
  NOR2_X1 NOR2_2389( .ZN(N6236), .A1(N6231), .A2(N6227) );
  NOR2_X1 NOR2_2390( .ZN(N6237), .A1(N5873), .A2(N6231) );
  NOR2_X1 NOR2_2391( .ZN(N6240), .A1(N6235), .A2(N6236) );
  NOR2_X1 NOR2_2392( .ZN(N6241), .A1(N5925), .A2(N6237) );
  NOR2_X1 NOR2_2393( .ZN(N6245), .A1(N5925), .A2(N6241) );
  NOR2_X1 NOR2_2394( .ZN(N6246), .A1(N6241), .A2(N6237) );
  NOR2_X1 NOR2_2395( .ZN(N6247), .A1(N5825), .A2(N6241) );
  NOR2_X1 NOR2_2396( .ZN(N6250), .A1(N6245), .A2(N6246) );
  NOR2_X1 NOR2_2397( .ZN(N6251), .A1(N5879), .A2(N6247) );
  NOR2_X1 NOR2_2398( .ZN(N6255), .A1(N5879), .A2(N6251) );
  NOR2_X1 NOR2_2399( .ZN(N6256), .A1(N6251), .A2(N6247) );
  NOR2_X1 NOR2_2400( .ZN(N6257), .A1(N5776), .A2(N6251) );
  NOR2_X1 NOR2_2401( .ZN(N6260), .A1(N6255), .A2(N6256) );
  NOR2_X1 NOR2_2402( .ZN(N6261), .A1(N5831), .A2(N6257) );
  NOR2_X1 NOR2_2403( .ZN(N6265), .A1(N5831), .A2(N6261) );
  NOR2_X1 NOR2_2404( .ZN(N6266), .A1(N6261), .A2(N6257) );
  NOR2_X1 NOR2_2405( .ZN(N6267), .A1(N5721), .A2(N6261) );
  NOR2_X1 NOR2_2406( .ZN(N6270), .A1(N6265), .A2(N6266) );
  NOR2_X2 NOR2_2407( .ZN(N6271), .A1(N5782), .A2(N6267) );
  NOR2_X2 NOR2_2408( .ZN(N6275), .A1(N5782), .A2(N6271) );
  NOR2_X4 NOR2_2409( .ZN(N6276), .A1(N6271), .A2(N6267) );
  NOR2_X4 NOR2_2410( .ZN(N6277), .A1(N5666), .A2(N6271) );
  NOR2_X4 NOR2_2411( .ZN(N6280), .A1(N6275), .A2(N6276) );
  NOR2_X4 NOR2_2412( .ZN(N6281), .A1(N5727), .A2(N6277) );
  NOR2_X4 NOR2_2413( .ZN(N6285), .A1(N5727), .A2(N6281) );
  NOR2_X1 NOR2_2414( .ZN(N6286), .A1(N6281), .A2(N6277) );
  NOR2_X1 NOR2_2415( .ZN(N6287), .A1(N5602), .A2(N6281) );
  NOR2_X1 NOR2_2416( .ZN(N6288), .A1(N6285), .A2(N6286) );

endmodule
