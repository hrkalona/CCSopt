//# 36 inputs
//# 39 outputs
//# 211 D-type flipflops
//# 3570 inverters
//# 2027 gates (955 ANDs + 528 NANDs + 431 ORs + 113 NORs)

module s9234(CK,g102,g107,g1290,g1293,g22,g23,g2584,g301,g306,g310,g314,g319,g32,g3222,g36,
  g3600,g37,g38,g39,g40,g4098,g4099,g41,g4100,g4101,g4102,g4103,g4104,g4105,g4106,g4107,g4108,g4109,
  g4110,g4112,g4121,g42,g4307,g4321,g44,g4422,g45,g46,g47,g4809,g5137,g5468,g5469,g557,g558,g559,
  g560,g561,g562,g563,g564,g567,g5692,g6282,g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g639,
  g6728,g702,g705,g89,g94,g98);
input CK,g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,g562,g563,
  g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,g41,g22,g44,g23;
output g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,
  g6374,g6728,g1290,g4121,g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,g4104,g4107,g4098;

  wire g678,g4130,g332,g6823,g123,g6940,g207,g6102,g695,g4147,g461,g4841,g18,g6725,g292,g3232,
    g331,g4119,g689,g4141,g24,g6726,g465,g6507,g84,g6590,g291,g3231,g676,g5330,g622,g5147,
    g117,g4839,g278,g6105,g128,g5138,g598,g4122,g554,g6827,g496,g6745,g179,g6405,g48,g6729,
    g590,g6595,g551,g6826,g682,g4134,g11,g6599,g606,g4857,g188,g6406,g646,g5148,g327,g4117,
    g361,g6582,g289,g3229,g398,g5700,g684,g4136,g619,g4858,g208,g5876,g248,g3239,g390,g5698,
    g625,g5328,g681,g4133,g437,g4847,g276,g5877,g3,g6597,g323,g4120,g224,g3235,g685,g4137,
    g43,g6407,g157,g5470,g282,g6841,g697,g4149,g206,g6101,g449,g4844,g118,g4113,g528,g6504,
    g284,g3224,g426,g4855,g634,g4424,g669,g5582,g520,g6502,g281,g6107,g175,g5472,g15,g6602,
    g631,g5581,g69,g6587,g693,g4145,g337,g2585,g457,g4842,g486,g2586,g471,g1291,g328,g4118,
    g285,g3225,g418,g4853,g402,g4849,g297,g6512,g212,g3233,g410,g4851,g430,g4856,g33,g6854,
    g662,g1831,g453,g4843,g269,g6510,g574,g6591,g441,g4846,g664,g1288,g349,g5478,g211,g6840,
    g586,g6594,g571,g5580,g29,g6853,g326,g4840,g698,g4150,g654,g5490,g293,g6511,g690,g4142,
    g445,g4845,g374,g5694,g6,g6722,g687,g4139,g357,g5480,g386,g5697,g504,g6498,g665,g4126,
    g166,g5471,g541,g6505,g74,g6588,g338,g5475,g696,g4148,g516,g6501,g536,g6506,g683,g4135,
    g353,g5479,g545,g6824,g254,g3240,g341,g5476,g290,g3230,g2,g6721,g287,g3227,g336,g6925,
    g345,g5477,g628,g5489,g679,g4131,g28,g6727,g688,g4140,g283,g6842,g613,g4423,g10,g6723,
    g14,g6724,g680,g4132,g143,g6401,g672,g5491,g667,g4127,g366,g6278,g279,g6106,g492,g6744,
    g170,g6404,g686,g4138,g288,g3228,g638,g1289,g602,g4123,g642,g4658,g280,g5878,g663,g4125,
    g610,g4124,g148,g5874,g209,g6103,g675,g1294,g478,g1292,g122,g4115,g54,g6584,g594,g6596,
    g286,g3226,g489,g2587,g616,g4657,g79,g6589,g218,g3234,g242,g3238,g578,g6592,g184,g5473,
    g119,g4114,g668,g6800,g139,g5141,g422,g4854,g210,g6839,g394,g5699,g230,g3236,g25,g6601,
    g204,g5875,g658,g4425,g650,g5329,g378,g5695,g508,g6499,g548,g6825,g370,g5693,g406,g4850,
    g236,g3237,g500,g6497,g205,g6100,g197,g6509,g666,g4128,g114,g4116,g524,g6503,g260,g3241,
    g111,g6277,g131,g5139,g7,g6598,g19,g6600,g677,g4129,g582,g6593,g485,g6801,g699,g4426,
    g193,g5474,g135,g5140,g382,g5696,g414,g4852,g434,g4848,g266,g4659,g49,g6583,g152,g6402,
    g692,g4144,g277,g6104,g127,g6941,g161,g6403,g512,g6500,g532,g6508,g64,g6586,g694,g4146,
    g691,g4143,g1,g6720,g59,g6585,I8854,g6696,I2272,I9125,g6855,I6783,g4822,I4424,g2097,g6895,
    I9152,g1835,I2919,I3040,g1770,g6837,g6822,I7466,g5624,I4809,g2974,g3537,I4757,g5457,g5304,g6062,
    g5824,g4040,I5343,I6001,g4162,g5549,g5331,I4477,g3063,g3612,I7055,g5318,g2892,g1982,I5264,g3638,
    I2225,I5451,g4323,g4086,g908,I1932,I5933,g4346,I8252,g6294,I2473,g971,I7333,g5386,I8812,g6688,
    g1674,g985,I3528,g1422,I8958,g6774,I5050,g3246,I4501,I2324,g1209,g2945,I4133,g5121,I6775,g1997,
    g1398,g3128,I4375,I8005,g6110,g1541,g1094,g5670,g5527,g2738,g2327,I9047,g4528,I6096,g2244,I3379,
    g6192,g5946,g2709,I3864,g1332,I2349,g4530,I6102,g1680,g1011,g2078,g1345,I2215,I3010,g1504,g5813,
    I7612,I7509,g5587,I5379,g3940,g3800,g3388,g2907,g1914,I9085,g2035,I3144,g2959,g1861,I9236,g4010,
    g3601,I2287,g927,I4273,g2197,I8270,g6300,g5740,I7501,I5777,g3807,g2876,g1943,g873,I6525,I5882,
    g3871,g2656,I3800,I8473,g6485,I2199,g900,I1927,g6708,I8834,I2399,g729,I3278,g1695,g6520,I8476,
    g940,I6677,g4757,g3902,g3575,g5687,g5567,g2915,g1931,g847,I3235,g1807,I3343,g1623,g6431,I8295,
    g709,g6812,I8984,I6576,g4700,g749,I1847,g3090,I4331,I9107,g2214,I3349,g4618,g4246,g6376,g6267,
    I5511,I6349,g4569,g4343,g4011,I5674,g4003,I8177,g6173,g2110,g1381,I3134,g1336,I8229,I3334,g1330,
    I7197,g5431,g4566,g4198,I7397,g5561,I4534,g2858,g1714,g1110,I4961,g3597,g2663,g2308,g3456,g2640,
    I6801,g922,I1947,g4693,I6283,I5484,g5570,g5392,g5860,g5634,g4334,g3733,I3804,g2575,I2207,I5153,
    g3330,g3355,g3100,g5645,g5537,g6733,I8891,g5691,g5568,g4804,g4473,g6838,I4414,g2090,g6610,I8696,
    g2877,g2434,I4903,g3223,g6796,I4288,I3313,g1337,g5879,g5770,g3463,g2682,I4513,g2765,I2578,g5358,
    I7012,I3202,g1812,I5421,g1076,I2115,g6069,g5791,I7817,g5924,g6540,g6474,I6352,g4564,I1865,g4202,
    I5622,I6867,g5082,g3876,I7349,I8144,g6182,g1175,g1375,I2411,g3118,I4366,g3318,I4593,g2464,I3596,
    g3872,g3312,g4494,I6004,I2870,g1161,g4518,I6066,g2215,g5615,I7372,g4567,I6139,I4382,g2265,I3776,
    g2044,g3057,I4282,I5600,g3821,I3593,g1295,I2825,g1143,g1285,g852,g3457,g2653,g5174,g5099,I6386,
    g4462,I3965,g2268,I8488,g6426,g6849,I9074,I6599,g4823,I2408,g719,g3834,I5027,g2295,g1578,g1384,
    I2420,g1339,I2370,g5545,I6170,I9128,g6864,g6898,I9161,g1838,g1595,g6900,I9167,g2194,I3331,g6797,
    I8961,g2394,I3537,I3050,g1439,I3641,g1491,I2943,g1715,I5736,g4022,I8450,I6280,g4430,g4933,I6625,
    g5420,I7086,g4521,I6075,g1672,I7058,g5281,I2887,g1123,I2122,g1477,g952,I4495,I2228,g5794,I7593,
    g1643,I2608,g3022,I4437,g2108,g2705,I3858,g3813,g3258,I8650,g6529,g1647,g2242,I3373,g1205,I2033,
    I5871,g3744,g774,I1859,g6819,I8994,g6694,I8800,g4379,I5848,g5905,g5852,g3519,g2740,I7856,g5994,
    g921,g1551,g1742,I2756,I4752,g2859,g6488,g6367,g2254,I3391,I8594,g6446,g2814,I4023,g4289,I5746,
    I6247,I6756,g4775,g6701,I8821,I8972,g6795,I3271,g1748,I2845,g1193,g5300,I6952,g2350,I3502,I8806,
    g6686,I3611,g1771,I2137,I8943,I2337,I2913,g1792,g1754,I2773,g6886,g2409,g1815,g894,I1917,g1273,
    g839,I5424,g3725,I6403,g4492,g6314,I8044,g4799,g4485,I9155,g6882,g2836,g2509,g2212,I6763,g4780,
    g3860,I5081,g2967,I4166,I9008,g5440,g5266,g3710,g3029,I5523,g3840,g843,g1543,g1006,I5478,g6408,
    g6283,g4153,I5545,I6359,g6136,g2822,I4031,g6706,I8913,g6743,I2692,g1037,g946,g1729,I2731,I5551,
    g4059,g4802,I6470,g3962,I5214,I2154,I4189,g2159,I5499,g3847,g5151,I6819,g3158,I4398,g6806,I8978,
    I4706,I7637,g5530,I7270,g6878,I5926,g2921,g1950,g6065,g5784,I6315,g4446,I4371,g2555,g6887,I4429,
    g2102,g6122,I7838,g6465,I8329,g6322,I8056,g1660,g1946,I3053,g6230,g6040,g5010,I6646,g4511,I6045,
    I6874,g4861,g2895,g1894,g6033,g2837,g2512,I2979,g1263,g5884,g5864,I8342,I2218,g1513,g878,I2312,
    g897,I3714,g1852,I4297,I8255,g6292,I8815,g6689,I5998,I1868,I7608,g5605,I5862,g3863,g1679,g1378,
    I2414,g4714,I6324,I2293,g5278,I6937,g3284,g3019,I4684,g2687,I8497,g6481,I4516,I6537,g4711,g3545,
    g3085,g2788,I3983,g6137,I7859,g5667,g5524,g6891,I9140,I2907,g1335,I2358,g3380,g2831,I4791,g6337,
    I8089,I4309,g2525,I2828,g3832,I5023,I2269,g5566,I7318,g3853,I5068,I3736,g2460,I6612,g4660,I7161,
    g5465,I7361,g2842,I4050,g1805,I2854,I6417,g4617,I3623,g4262,I5713,I7051,g5219,I2221,g3559,g2603,
    g4736,I6366,g2485,I3614,I7451,g5597,I2703,g1189,I8267,g6297,g4623,g1947,I3056,I5885,g3746,I7999,
    I7146,g5231,I6330,g4560,I7346,g5531,I3871,g2145,g6305,g4375,I5840,g4871,I8761,g6563,g3204,I4441,
    g4722,I6346,g710,I4498,g2686,g829,g5113,I6753,g1632,g760,I2067,I4347,I8828,g6661,I8872,I8411,
    g1653,I2630,I3782,I8727,g6536,g2031,I3140,I5436,g3729,g2252,I3385,g5908,g5753,g2958,I7472,g5626,
    g2176,I3319,I2716,g1115,I5831,g3842,g1160,I5182,g3271,g5518,I7258,g5418,I5382,g3952,g2405,I3543,
    I2848,g1917,I3016,g2829,g2491,I3946,I7116,g5299,I4019,g1841,I5923,I6090,g4393,I4362,I3672,g1656,
    g3040,I4255,I3077,I6485,g5593,I7355,g3440,I4678,g3969,I5233,g6312,I8040,I4452,g2117,I4173,I8217,
    g895,I6456,g4633,g4523,I6081,g1233,I2231,I6649,g4643,g4293,g5264,g4943,I9158,g1054,g5160,g2796,
    I3999,I6355,g2473,I3605,I3099,g1519,I8576,g6436,I2805,I8866,I3304,g1740,I4486,g3093,g5521,I7261,
    I3499,g1450,I8716,g6518,g1725,g1113,I7596,I8875,g3875,I5106,g2324,I3478,I4504,g2726,I2119,g5450,
    g5292,I5037,g3705,g5996,I5394,I8644,g4499,I6015,I2352,I6063,g4381,g6746,I8916,I2867,I8699,g6573,
    g2177,I3322,g5179,g5379,I7035,I2893,g1236,I7646,I3044,g1257,I2196,g3839,I5040,g6932,I9217,g4273,
    I5728,g5658,g5512,g6624,I8730,I6118,g4406,I6318,g4447,g2276,g2849,g2577,I3572,g1787,I2835,I5442,
    g3731,g2670,I6057,I8524,g6496,g6526,g1461,I6989,g5307,I2614,g1675,g1101,I2125,g3343,g3571,I2821,
    g1221,g4712,g6576,g6487,I6549,g4699,I8258,g6293,I8818,g6690,I3534,g2245,I3382,I3729,g2436,I3961,
    I5454,g3874,g2291,I3434,g5997,g5854,g4534,I6114,I3927,I5532,g3861,g1684,I2668,g6699,g1639,g815,
    g1338,I2367,g1963,I3074,I8186,g6179,I6321,g4559,I4226,g1109,g1791,I8975,g6791,g2256,g889,I2306,
    g896,g3792,g4745,g2819,g2467,g4014,I5316,I8426,g6424,I5412,g4034,I6253,g4608,g2088,g2923,g1969,
    g2408,I8614,g6537,I3513,g2488,I3617,g1759,I2782,g2701,I3855,I7190,g5432,g6691,g6524,I6740,g4781,
    g4513,I6051,g6794,g5596,g1957,I3068,I3352,g6119,I7829,I2904,g1256,g6319,I8051,g1049,g5901,g2886,
    g1966,I6552,g4702,I4059,g1878,g4036,I5337,g3094,I4337,I4459,g2134,I8544,g6453,g4679,I6269,g6352,
    I8110,g6818,I8991,g6577,I3288,g1710,g3567,g3074,g1284,I5487,I7704,g5723,g848,g5092,g4753,g1498,
    I2479,I2763,g2870,g2296,I3022,g1426,I4261,g1857,I2391,g4382,I5857,g3776,g3466,g6893,I9146,g1833,
    I3422,g1641,g5574,g5407,I3749,g2484,g3593,g2997,g6211,g5992,g2650,I3794,g5714,I7475,g932,I8061,
    g6113,g4805,I5328,g1584,g743,g4111,I8665,g1539,I5109,I3546,I2159,I6570,g4719,g2136,g1395,I4664,
    g2924,I8027,g6237,I4246,g2336,I3488,I7336,g716,I1832,I3560,g1673,g736,I1841,g4770,g2768,g2367,
    I8174,g2594,I3723,g4798,I6464,g6325,g6821,g6785,g4188,g2806,g2446,I3632,g3450,I4688,I3037,g1769,
    g6939,I9230,g1052,I3653,g1305,I3102,I2315,g1222,I2811,g6083,g5809,g2887,g1858,I2047,g6544,I6607,
    g4632,g4281,g5889,g5742,I7164,g2934,g2004,g2230,I3355,g4437,I5948,I5388,g4302,g4068,I5865,g3743,
    I7814,g4579,g4206,g4869,g4662,g6306,I8030,I3752,g5375,I7029,I8107,I6337,g1730,g1114,g3289,g3034,
    I2485,g3777,I6587,g4803,I8159,g6167,I6111,g4404,g3835,I5030,I6311,g4444,I8223,g2096,I3212,I9143,
    g3882,I5119,g1070,g2550,I3665,I6615,g3042,I4671,g2928,I2880,g2845,g2565,g1897,I2992,g6622,I8724,
    I2537,I5896,g3879,g2195,g4265,I5716,g2891,g1884,g2913,g1925,I6795,I3364,g1648,g5384,g5220,I9134,
    g6904,I9179,g4786,I6448,g3799,g6514,I8462,g4364,I5825,I8447,g6410,I3770,I5019,I2417,I7683,g5702,
    I9044,g3541,g2643,I2982,g1678,I2658,I6414,I2234,g1331,I2346,g4296,I5753,I2128,I3553,I6020,g4176,
    g3332,g3079,I7167,I6420,g6695,I8803,I2330,g1122,g3209,I6507,g4644,g4532,I6108,g1682,I9113,I1856,
    g3802,g2481,I3608,g5627,g931,g2692,I3840,I4217,g2163,I3215,I4066,g2582,g5551,I7295,g5686,I3886,
    I6737,g2497,I3626,I5385,I6956,g2154,g1755,I2776,g4189,I5597,g6792,g4706,I6308,g6416,I8243,g6286,
    I8417,g6420,g3901,I6630,g5774,I3675,g6522,I8482,g6115,g1045,I3281,g1761,I7039,g5309,I7484,g5630,
    g1173,I2185,I4455,g2118,I8629,g5273,I6930,g2040,I2476,I1853,g2783,I3979,g2112,I3240,g1283,g853,
    g2312,I3462,g1369,I2405,I6750,g4771,g6654,I8758,g3714,g3041,I7583,I3684,g1733,I5006,g3604,g6684,
    g1059,I2552,g2001,I3112,I5406,g3976,g5572,g5399,I3109,I3791,g2293,g1567,g6880,I8653,I5496,g1535,
    g1088,g4639,I8527,g5543,I3808,g2125,I7276,g3881,I2355,g1177,I5409,g4309,g4074,g2828,g2830,g2494,
    g2727,g4808,I2964,g821,I1880,g6612,I8702,g5534,g5729,I7494,I6666,g4740,g6875,g1415,g1246,g4707,
    g6417,I8261,I7404,g5541,g3076,I8512,g6441,g3889,I6528,g4815,g1664,I2643,I2237,g6234,g6057,I3575,
    g5885,g5865,g6328,I8066,g1203,I5445,g6542,I8538,g6330,I8070,g1721,I2721,I5091,g3242,g6109,g2932,
    g1998,I8456,g5903,I3833,g2266,I2318,g4715,I6327,I1924,I8966,I5169,I6410,I5376,g3500,g2647,g4498,
    I6012,I2057,g1502,I5059,g3259,I5920,g4228,I2457,g1253,I3584,I5868,g3864,I2989,I2193,g5436,g3384,
    g2834,g1940,I3047,g2576,I3687,g2866,g1905,g5135,g2716,g3838,I7906,g5912,I3268,I3019,g3424,g5382,
    I7042,I5793,g3803,I3419,g1287,g6902,I9173,I6143,g4237,I6343,g4458,g846,g1671,g5805,I7604,I5415,
    g3723,I3452,I5562,g5022,g1030,I8279,g6307,I4492,g6490,g6371,I2321,g898,I9002,g3477,g6166,I7892,
    I8162,I6334,g4454,g2241,I3370,g1564,g5916,I3086,I8503,I8843,g6658,g6649,I8745,I6555,g4703,g1741,
    I2753,I6792,g5097,g3104,I4351,g1318,g2524,I3647,g2644,I3788,g6698,g1638,g754,I6621,g2119,g1391,
    I5502,g1108,I2134,I3025,g5437,I7119,g4385,I3425,g1274,I9092,g2109,g2818,g2867,g1908,g1883,g1797,
    g5579,I7478,g5628,g5150,I7517,g2893,g1985,g5752,I8232,g6332,g5917,I6567,I3678,g1690,g2975,I4176,
    g1631,I2967,I8165,g1048,I5430,g3727,g2599,g5042,I6672,g1711,I2712,I3635,g6652,I8752,g5442,g5270,
    g1055,I2570,I2860,I5475,I4743,I3105,g2170,I3301,g2370,I3522,I5913,g6193,g5957,g1333,I3255,I8552,
    g6455,g1774,I2817,g4766,I6406,I5397,g1846,I2940,g5054,g4816,g4801,g4487,g6834,I5991,I7110,g5291,
    g3534,I5910,g3750,I3755,g5296,I6946,I8687,g6568,I6933,g5124,g2544,I3662,I8662,I5609,g3893,I4474,
    g3052,g1176,g3014,g6121,I7835,I7002,g5308,g766,g3885,I5124,g4226,g4050,g2106,g2306,g1743,g1320,
    g2790,g2413,g6232,g6048,I5217,g3673,I8570,g6433,I8860,I4480,g3073,g1994,I2275,g909,g6938,I9227,
    I5466,g3787,g4173,I5577,I8710,g6517,g2461,I7590,I3602,I3007,g2756,g2353,g2622,I3764,I3059,I3578,
    g1484,I3868,g5888,g5731,g838,g6519,I6289,g4433,I9024,g6803,I5448,g3960,I3767,g5787,g5685,g2904,
    g1991,g6552,g6606,I8684,I3581,I5333,g3491,I2284,g4718,g4767,g4601,I3261,g1783,g1847,g3207,I5774,
    I9077,g6845,I8659,g6523,g4535,I4976,g1685,I2671,I8506,g6483,g2841,g2541,g4582,g4210,I4229,g2391,
    I8626,I2029,g964,g791,g2695,I3843,g2637,I3779,g4227,g5439,g3798,I9104,g5063,I3284,g6570,I5692,
    I6132,g4219,g6525,I8491,g6710,I8840,I5418,I6680,g4713,g4721,I2588,g2416,I3556,g3095,I4340,g3037,
    I4252,g845,I2204,I5493,I8180,g6176,I4220,g2164,I7966,I8591,g6448,g2315,I3465,g5866,g6879,g6607,
    I6558,g4705,g4502,g5049,I6685,g6836,I1958,I1942,g3719,g3053,I8438,g5575,g5411,I8420,g6422,I3388,
    g1324,g2874,g1849,g3752,I4935,g3932,I3028,I5594,g4388,g3724,I3428,g1825,I2973,g1687,I7254,g5458,
    g5922,I3247,g6615,I8707,I7150,g5355,I4327,g4428,g3786,g5584,g5539,g5896,I2653,I3826,g3364,g3114,
    I8515,g6492,g4192,g3054,I4279,g4002,I4303,g2612,I8300,g6299,I8002,g2243,I3376,g3770,I9014,g6820,
    I3638,g1772,I5723,g3942,g4741,I6371,I8641,g5052,I6692,g6832,I9021,g4910,I2648,g980,g2234,I3367,
    I9082,g1890,g1359,I3883,g2574,I4240,g2165,g2330,g1777,g4609,I6182,I8441,g4308,I2050,g1734,I3758,
    g2041,g5086,g4732,g6142,g951,I8969,g2800,g2430,g5730,I7497,g2554,I3669,g4758,I6382,I2839,I3861,
    g1834,g6905,I9182,I3711,g1848,I4986,g2213,I3346,g5897,g5025,g4814,g6515,g5425,I7091,I2172,I2278,
    g917,I7796,I4681,g2947,g1480,g2902,g1899,g6697,I2143,I2343,g4222,I5481,g3297,g3046,I3206,I6546,
    I2334,I6809,g5051,I5743,I6995,I5890,g3878,I3509,g3963,g3791,I8884,g6704,I5505,g1688,I2688,g4752,
    I6434,I2961,I6231,g4350,g4509,I6039,g5087,I9095,g5801,I7600,g2155,I3274,I9208,g6922,g4640,I3093,
    g965,I3493,I3816,g2580,g1326,I8235,I6099,g4398,I8282,g6309,g3049,I4270,g6528,I8500,g1760,I2785,
    g4493,g6351,I1850,g834,I8988,g6787,g6530,I4777,g5045,I8693,g6655,g5445,g5274,I4799,I8548,g6454,
    I7193,g3498,g2634,I5854,g2619,I3761,I8555,g6456,I3519,g2872,g1922,g1608,g1220,I6292,I8240,I9164,
    g6885,g4397,I9233,g1192,I7640,g5773,I7073,g6884,I9119,I2593,g5059,I6697,g5920,I7692,I9038,g2457,
    I3587,g5578,I6444,g4503,g4655,g1423,I2442,g923,g3740,I7176,g1588,g798,I8113,g6147,I7342,I2182,
    I3830,g3162,I4402,g5261,I6918,I4294,I6543,g6618,g1665,g5926,g2158,g6143,I7865,g4562,g6235,g2598,
    I3726,g1327,I2521,g1063,g5415,I7081,g3452,g2625,I7996,I5400,g6566,I8582,I8494,g6428,I6534,I8518,
    g6494,g1681,g4723,I8567,g6432,g6134,I7852,g5664,g5352,g2232,I3361,g6548,I6927,g3086,I2724,g2253,
    I2179,g3486,g2869,g2813,I2379,g1696,I2700,I6885,g4872,g4497,g3504,g2675,g1732,I2738,I5116,I3909,
    g1001,I3441,I7069,g3070,I8264,g6296,g6621,I8721,I7469,g5625,g3897,g3251,g3263,g1472,g1043,I5977,
    g4319,I8521,g6495,I6036,g4370,I2611,g893,g6412,g1739,g1116,I3531,g1593,g3967,g4249,I8470,g6567,
    I8585,g6533,g4460,g996,I2041,g3331,I3890,g4772,g5247,g4900,g4531,I6105,I5633,g3768,I8878,I2663,
    I3505,I8647,g3766,I4955,g1533,g5564,I5103,I3650,g3801,g3487,I3013,I5696,g2691,g2317,I6798,g5741,
    g5602,I2802,g1204,I3474,g5638,g6160,I5508,g3867,g6933,I9220,I5944,g4356,g2962,g2008,g6521,I8479,
    I9098,I5472,g3846,I8981,g6793,g2506,I3080,I8674,g1820,I5043,g3247,I6495,g4607,g1936,g1756,I6437,
    g4501,g3173,I4410,g4399,I6302,g4440,I8997,g6790,g1117,I8541,g6452,g1317,g2608,I6579,g5993,g3557,
    I3569,g1789,g2111,g2275,g5466,I8332,I7701,g5720,g3369,I4646,I8153,g6185,g3007,g2615,I9101,I2864,
    g5571,g5395,g5861,g5636,g3868,g2174,g3459,g2664,I1877,g1775,g5448,g835,g5711,g6835,I9028,g1581,
    g910,I6042,g4374,g1060,g2284,I3431,I6786,g4824,g1460,g3793,g6611,g2591,I3720,g3015,I2749,I6054,
    g4194,g5538,I6296,g4436,g2602,I2623,I5460,g5509,I7251,g4400,I5899,g1937,g6541,I8535,I9185,g6877,
    I8600,g6451,g2931,g1988,g4760,I8074,g5067,g1190,I2175,g6353,g5873,g2905,g4167,I8910,g6802,g2628,
    g1156,g2515,g5493,I7065,g5256,g5077,I6706,g4731,g4220,I5644,I5177,I4276,I3161,g1270,g5381,I4667,
    I9131,g6901,I9170,g3771,I8623,g3216,g1824,g5552,I8453,g6457,I2424,I1844,g862,g2973,I4170,g1954,
    I3065,g3030,I4243,g1250,I5739,g1363,g1837,I5463,g5950,g1053,g1738,I8668,g6574,g6484,g2440,g3564,
    g2618,g6714,g6670,I5520,I5668,g3828,g4284,I8285,g6310,g3732,I5391,g6580,g6491,g6032,g5631,g5536,
    g3108,g6876,I6362,I4354,g3308,g3060,I6759,g4778,g2875,I6377,g4508,I8809,g6687,g6623,g6076,g5797,
    g6889,g5751,I7506,I3316,g1344,g3589,I7481,g5629,I3034,g2410,I3550,g1627,g2777,g6375,I8189,g2884,
    I2044,g3084,g2839,g2535,I5084,I7960,g5925,g899,g6651,I8749,g3448,g4565,g4195,I3681,g1821,I5053,
    g3455,g6285,g2172,I3307,g6937,I5568,g4533,g2667,I3811,g1683,g1017,g2343,g5168,g6339,I8093,g3196,
    I4433,g4914,I5002,I5630,I7267,I5157,g3454,I9035,I9203,g6921,g1731,I3258,g1735,I2745,I8273,g6301,
    g6809,g5890,g1782,g1935,I6452,g4629,I5929,g4152,g1661,g6252,g6231,g6044,g5011,I8444,g6421,g3067,
    g784,I1838,I7077,I8485,g861,I2946,g1587,g2792,I2584,I5433,I2281,I5626,g3914,I4334,g1646,I2617,
    g5869,g4191,g1084,I7808,g854,g1039,I2449,g6778,I6425,g5573,g5403,I5056,g4619,I2831,g2518,I3644,
    g1583,g1702,g1107,I2382,I8414,g6418,I8946,g1919,I2916,g2776,g2378,g4784,g1276,g2283,I3294,g1720,
    g3852,g6572,I4762,g2862,g5532,I6635,g2264,I3405,g6712,g6676,g851,I6766,g4783,I6087,g4392,g6543,
    I6305,g4441,g2360,g1793,g2933,I4123,I2620,g4190,I5526,g3848,g4157,I8335,g6308,I8831,g6665,g6931,
    g1546,I2873,I2037,g6534,I8881,g3605,I4802,I5603,g2996,I3942,g1503,I5439,g3730,g6742,g6560,g2179,
    I3328,g6014,I9122,g4704,g6414,I5702,g3845,I4258,g5383,I7045,g4903,g5303,g6903,I9176,g3441,g2835,
    g1407,g4250,g6513,I8459,g913,g4613,I5952,g4367,g4810,I6488,g2882,g1854,I7352,g5533,g3075,g872,
    g6036,I8632,I2364,g6531,I2808,g3772,I6582,g4765,I6689,g2981,I8579,g6438,I8869,I4489,g3458,g865,
    I2296,g3890,I4192,g4170,I3659,I4471,I7170,g5435,I8276,g4929,g2744,I1935,g2802,g2437,g949,I8564,
    I5320,g4626,g4270,g1340,I2373,g3480,g2986,g6653,I8755,I7802,I7061,I7187,g5387,g6579,g5116,I5987,
    g4224,g5316,I6976,I2635,g5434,g2864,g1887,I6430,g855,g4894,g4813,g1249,g4620,I5252,I2791,I7514,
    g5590,I2309,I2140,I8888,I3691,g5210,g6786,I6564,I8171,g6170,I8429,g6425,I7358,g6164,I8156,g6233,
    g6052,I2707,g4292,I7695,g2968,I5078,I2890,g4526,g3859,I7107,g5277,I5907,g3883,g1762,g2889,g1975,
    g4403,g4603,g6532,g4443,I5517,I9041,g4439,g5117,g6553,I5876,g3870,g2175,g2871,I2604,g3183,I4420,
    g2722,I4462,g2135,I8309,g6304,g1556,g3779,I8246,g3023,g1928,I3031,I7811,g5921,I7698,g1064,g6888,
    I2998,I6048,g4376,I7339,g4276,I5731,I4249,I3004,I1825,g4561,g2838,g1747,g3451,I2162,g1563,I9011,
    g2809,g1586,g4527,I6093,I2290,g4647,g3346,I4623,I5236,g2672,g2231,I3358,g4764,I6400,g5995,g6844,
    I7173,I3785,I6780,g4825,g1394,g1206,I6023,I2735,I2728,g1232,g1557,g4046,I5556,g2104,g1372,g2099,
    g1366,I4519,I2385,g6707,g1471,I2464,g4320,I3906,g4394,g6189,g3043,I4264,g3748,I6816,g5111,I3516,
    g2754,g2347,g4242,g1254,g1814,g6575,g6486,g4516,I6060,g6715,g6673,g4716,g5250,g6604,I8678,g1038,
    I6397,g1773,I2814,I2131,I7104,g4299,I5756,g6833,g6535,g5453,g2712,g2320,g6711,g4016,I8620,g6539,
    I8531,g6896,g1836,I2922,g5423,g6116,g6461,I8897,g1918,I3244,I7490,g5583,I4980,g3546,g5853,I4324,
    g2961,I5071,I3340,g1282,I5705,g6162,I8150,g6419,I6723,g4761,g2927,g1979,g4360,g6930,g2885,g5535,
    g6565,I2445,g2660,g2946,g938,g4435,g4517,g5717,I3656,I4794,I2491,g2903,g1902,I8635,g6363,I2169,
    g942,g6730,g3775,I8432,g3922,I7463,g5622,g6385,g6271,g6881,I9110,g3980,g2036,g1764,g706,I6441,
    g4624,g4915,g4669,g2178,I3325,g2679,I3823,g6070,I3525,I4285,I3310,g1640,g6897,I2925,g6561,g3460,
    I8226,I4510,g2753,g6890,g5452,I4291,g5894,g2805,g2443,I1938,g1788,g2422,I6772,g4788,g6480,I4312,
    I6531,g4402,g4017,I1862,I2240,g4615,g837,g5661,I1835,I3590,g1781,I7686,g5705,g1842,g1612,g1219,
    g6427,g6087,I6942,I8767,g6619,g6365,g3501,I3222,g1790,g6447,I6244,g6439,I2958,I9116,g6298,g5084,
    g4727,I5654,I3797,I6992,g2346,I5837,g3850,g2433,I2388,I6573,I3563,g6290,I2601,g2752,g6373,I8183,
    g3363,g3110,g5919,I7689,I2428,g4563,I2190,I3408,g3453,g6369,g2042,I3155,I5249,g6578,g6489,I6540,
    I3291,g1286,g2364,g2233,I5612,g1911,g5136,g3912,g3505,I2741,I8940,g6783,I2910,g1645,I3071,g5647,
    I3705,g2316,I3471,I2638,g844,g5546,g5388,g3857,I4465,g6015,g5857,g6415,I6126,g4240,I5686,I2883,
    I8671,I7707,g6239,g2103,I2327,I5708,I8857,I5640,g5120,g6429,g2706,I3773,I2165,I2212,g2888,g1972,
    g5565,I4195,g2173,g2029,g2171,g1934,g2787,g2956,g4151,I8638,I3819,I3836,g1832,g1806,I7587,g4769,
    g4606,I2949,g3778,g6188,I6949,g4185,g1898,I2995,g3782,g6562,g6114,g5892,g4451,I8290,I4306,g4229,
    I7284,g4614,g6564,I5324,I7832,g5943,I5469,g1953,g3267,I4321,g1819,I2877,g2957,g6685,I2952,I6072,
    g6609,I7113,I8034,I3062,g1776,g2449,I3620,g6450,g2865,g6883,g4837,I8509,g6437,g2604,I4267,g2098,
    g4251,g945,g6466,g5915,I7679,g4622,I8467,g6789,g6291,I2150,g6165,g6571,I8597,g5110,I5699,g5310,
    I3298,g1650,I2627,I3485,g3527,g809,I1874,g849,I5606,I5879,I2361,g3970,g1594,g6538,g6469,I3083,
    I2857,I7643,I3708,g2086,I3198,g2728,I4468,g2583,g3320,g6067,g5788,g1275,g6467,g1322,g4520,g1328,
    g4431,I5938,g4252,g1321,g3906,g2470,g3789,g5064,g2025,g6493,g5899,g4790,I5843,g4405,I4964,g1550,
    g4380,g4286,I4198,g3299,g5563,g4911,I3733,g6700,g1891,I2986,g5237,g5083,g3892,g2678,I3225,g1813,
    g6442,g4225,g2766,g2361,g2087,g1352,g2105,I7143,g5323,g2801,I4003,g5089,I5065,g714,I3540,g1670,
    g4980,g4678,g2748,I3923,g1823,g3478,g1142,g2755,g2169,g5242,g5085,I8168,I8863,g1255,I5033,I7799,
    g6817,g3728,g3082,I4315,g3482,g2713,g6444,g1692,I2696,g6605,I8681,g1726,g2091,g1355,g1960,g5295,
    g3751,g2061,g2007,g1411,I6250,g4514,g2059,g1402,g2920,g2157,g6118,g2767,I4358,I4821,I3090,g1112,
    g1267,g4510,g1319,g5918,g3002,I8573,g6435,I4483,I5514,I8713,I4507,g1329,I2340,I3694,g1811,I2788,
    g857,g5872,g2581,I2760,g3866,I8907,I9137,g1830,I7264,I8435,g6411,g6734,I8894,g1703,g4215,I5637,
    I2779,g6074,g3064,g3785,g1624,I2581,g5895,g4314,g4080,g6080,g1075,I8603,I4391,g6713,g6679,g1644,
    g6569,g2030,I3137,I5490,I4223,I8220,g4768,g2826,g1699,g4386,g2861,g4806,I8423,g6423,g5050,g1724,
    I8588,g6443,I4522,g1174,g842,g4434,g3083,g4322,I3232,g2609,g4687,g6527,g6108,I7153,g2883,I6084,
    g4391,g4182,I3096,I3496,g715,g5708,g1119,g2066,g1341,g3150,g1315,I8103,I3395,I3337,g4496,I6008,
    g1577,g4550,g3773,I4537,g5958,g5818,I2147,g6608,I8690,I5615,g830,g3769,g3622,g2827,g3856,g3836,
    g3212,g1853,g2333,g6287,g3844,g4807,I5223,I6561,I2596,g6161,g856,g6361,I8147,g2196,g2803,g4159,
    I6986,g5230,g6051,g804,I1871,g2538,g1325,I3481,g6242,g4248,g4692,I7805,I3599,g4726,g4154,I5548,
    g1636,g3921,g3512,g5540,g1106,g6732,I2842,I5893,g3747,I2460,g3462,g2381,I6789,g6043,I7871,g6097,
    I3001,g4218,g4267,I5720,g2390,g2397,g5199,g1046,g2505,g3788,g6034,g6434,I6299,g4438,I5750,I2929,
    g6347,g1191,g3192,I3746,g5947,g3485,g1637,g2631,I8656,g3854,g6445,g2817,g4519,g6413,I8249,I5790,
    I6078,g4387,I6340,g5923,I3468,g1802,I6959,g3219,I4318,I7634,g5727,I5427,g3726,g3031,g6117,g5880,
    g1642,g6482,I5904,g3749,g5886,g6657,I3152,g1334,I2053,g5114,I5403,g5314,I6972,I2453,g1654,I5529,
    g3975,g3911,I5148,g6581,g1880,g1603,I5618,g2772,g2743,g6784,g2890,g1875,I4300,g1978,g1387,g3796,
    g1659,I3629,g3124,g2856,g2010,g2734,I3902,g4524,g836,g3540,g5887,g1542,g3177,I3717,I6895,I5542,
    g4577,g4717,g4465,g5433,g3742,g5017,g2863,g3199,g5550,g3781,g5891,g3898,g3900,g1118,g3797,g6850,
    g6163,g5726,g3510,g3910,I5457,g2688,g2857,g3291,g2976,I2402,I6923,g1056,g3502,g1529,g3984,g1649,
    g1348,g5248,g4636,I2394,g5255,I9031,g2760,g3488,g6709,I4587,I6733,I7487,g4187,I5591,I9005,g3886,
    g2779,g4904,g4812,g1279,g1111,g5112,g2588,g6449,I6769,g4763,g3136,g2739,g1549,g947,g6894,I9149,
    I5851,g3739,g4536,g6735,I2970,g858,I3115,I3251,g6303,g3465,g3322,g3783,g4522,g6440,g2043,I3158,
    g6039,I8764,g3096,I4343,g3851,g1552,I8617,g850,g5576,g4537,g4410,g5149,g6276,g4612,g2914,g6616,
    I2376,g3342,g4328,g4092,g4351,I7963,g3481,g2820,g2936,g2026,g3354,I5204,g5119,g5701,g1358,g5577,
    g4213,g6120,g2922,I6812,g6788,g5893,g2908,g6095,g2060,g6617,g6906,g5975,g5821,g4512,g6702,g3001,
    g4166,g6516,g6409,I3148,g3761,g4529,g4773,g3830,g2079,g4155,g6892,g6936,I2955,g2840,g3745,g5544,
    g4450,g1559,I6069,g4463,g943,I8837,g6078,g5061,I6701,g6478,g866,g6035,g4720,g3677,g3140,g2954,
    g2966,g5046,g6656,g4193,g2032,g1749,g3814,g5391,g2568,g2912,g5467,g2357,g1323,g4625,g4232,g1666,
    g4938,g5019,g6236,g6295,g5684,g1528,g1351,g5115,g5251,g5069,g5315,I5094,g1655,g1410,g5167,g6899,
    g929,g5385,g2778,g3370,g2894,I7007,g4163,g4525,g3483,g6194,g1829,g5542,g3306,g2998,g4158,g1555,
    g3790,g2039,g3187,g3387,g3461,g4587,I6033,g4179,g5554,g5455,g3904,g3200,g2919,g2952,g4455,g3599,
    g4545,g4416,g5090,g4020,g6212,I7910,g5456,g5649,g4507,g2764,g6430,g5155,g3016,g6229,g5260,g6289,
    g4628,g4515,g2120,g6479,g2906,g2789,g5118,g2771,g6620,g5193,g4967,I5360,g3532,g3536,g3539,g3544,
    g5598,g6249,g4666,g4630,g4627,g3629,g3328,g6085,g4648,g4407,g5232,g2340,g5938,g5909,g3554,g2941,
    g3903,g1474,g6640,g6549,g4172,g3930,g4372,g3490,g4667,g4653,g4651,g3166,g3366,g6829,g3649,g6911,
    g3155,g3698,g6270,g4792,g1417,g4471,g6473,g6397,g1628,g4621,g3953,g5158,g4993,g6124,g6324,g3880,
    g2121,g6394,g3279,g3619,g3167,g5311,g5013,g4468,g3367,g3652,g3843,g3533,g4593,g4277,g3686,g5180,
    g4950,g5380,g4160,g3923,g3321,g2089,g6245,g3670,g3625,I5359,g5559,g5024,g6144,g6344,g6272,g2948,
    g2137,g6259,g2955,g6088,g6852,g6847,g6923,g6918,g6917,g5515,g5364,g1499,g4835,g3687,g4271,g4004,
    g4611,g3985,g4300,g3341,g6650,g4541,g4199,g3645,g5123,g4670,g3691,g4209,g3816,g4353,g3989,g6336,
    g6246,g6768,g6750,g4744,g3434,g3659,g5351,g5326,g3358,g5648,g6934,g3275,g3311,g5410,g3615,g2062,
    g3374,g4600,g4054,g6096,g1436,g5172,g4877,g3180,g5618,g5506,g5143,g6913,g5235,g4580,g2085,g6266,
    g5555,g5014,g2166,g6248,g6342,g6264,g5621,g5508,g3628,g6255,g6081,g3630,g6692,g3300,g6154,g6354,
    g4184,g3934,g5494,g5443,g4384,g4339,g3971,g4838,g3123,g3323,g4672,g4635,g4631,g2733,g3666,g6129,
    g6329,g3888,g2073,g5360,g6828,g4285,g3351,g6830,g3648,g3655,g1706,g6068,g4044,g6468,g1609,g3172,
    g3278,g3372,g2781,g3618,g3667,g3143,g3282,g6716,g6682,g6149,g3693,g3134,g3334,g6848,g3741,g6843,
    g5153,g5209,g5353,g5327,g6241,g1808,g3113,g5558,g5018,g6644,g6152,g6258,g4178,g3959,g1575,g4378,
    g4831,g5492,g5441,g5600,g5502,g6614,g6556,g4947,g3360,g6125,g1419,g918,g3641,g4873,g4037,g2896,
    g4495,g3913,g3379,g5175,g5094,g3658,g6061,g5500,g5430,g5074,g3611,g4042,g5184,g4442,g4239,g4164,
    g3958,g2807,g5424,g6145,g3997,g3425,g3694,g6345,g6273,g3132,g3680,g6637,g3353,g2142,g2255,g6159,
    g2081,g3558,g5499,g5451,g4389,g4171,g3956,g6315,g3849,g4371,g4429,g4253,g4787,g2937,g6047,g6874,
    g6873,g2267,g1716,g5444,g1574,g5269,g4684,g4584,g4791,g3936,g6243,g6935,g2746,g4759,g4500,g6128,
    g5414,g6130,g5660,g3375,g4449,g4266,g3651,g4865,g4776,g2953,g2068,g3285,g4833,g5178,g5679,g5378,
    g3339,g1689,g5182,g2699,g2747,g6090,g4362,g3996,g3672,g4052,g3643,g4452,g3820,g6056,g1826,g6148,
    g6348,g5560,g5044,g3634,g6155,g6851,g6846,g3551,g3099,g3304,g4486,g3499,g4730,g5632,g5095,g4794,
    g6260,g5495,g1138,g3613,g6318,g3865,g901,g5164,g5194,g5233,g2821,g5454,g4549,g5553,g5012,g6321,
    g3873,g3660,g6625,g4045,g4445,g4235,g6253,g4373,g4001,g5189,g4491,g6909,g4169,g3966,g5171,g4369,
    g3999,g3679,g4602,g5371,g3378,g5429,g5956,g5783,g4868,g4774,g5675,g3135,g4459,g4245,g3335,g3831,
    g3182,g3288,g3382,g4793,g4015,g2107,g6141,g6341,g6261,g6645,g3632,g3437,g2853,g3653,g5201,g4859,
    g3208,g2551,g3302,g6158,g5449,g5246,g5604,g5098,g4021,g5498,g1585,g6275,g6311,g3837,g4671,g4645,
    g4641,g4247,g4007,g4826,g5162,g5088,g5362,g3296,g5419,g2935,g6559,g5728,g5623,g5486,g5185,g3171,
    g3371,g6628,g2138,g4165,g3927,g4048,g4448,g3815,g3281,g4827,g4333,g3964,I2566,g1633,g3684,g4396,
    g3338,g2056,g5406,g3309,g5635,g5682,g5487,g6123,g6323,g3877,g3759,g5226,g6151,g3449,g6648,g5173,
    g5373,g4181,g3939,g2720,g4685,g4591,g5169,g5093,g5369,I4040,g3362,g6343,g6268,g6693,g6334,g3858,
    g6555,g2909,g2092,g4041,g6313,g3841,g5940,g4673,g4656,g4654,g5188,g6908,g6907,g5216,g6094,g4168,
    g3925,g4368,g3998,g5671,g3678,g5428,g4058,g3635,g2860,g3682,g3305,g2960,g5910,g5816,g3755,g2659,
    g1686,g5883,g3373,g5217,g4866,g4863,g4777,g3283,g3602,I2574,g5165,g6777,g6762,g3718,g1157,g3767,
    g4688,g4568,g1784,g2021,g6799,g4948,g6782,g2794,g3203,g6132,g6238,g6153,g4183,g3965,g4383,g6558,
    g5181,g3689,g4588,g2419,g5197,g4161,g3931,g4361,g3995,g3671,g4051,g6092,g2323,g5562,g5228,g3609,
    g6262,g6736,g3758,g4043,g3365,g1558,g5673,g4347,g3986,g3133,g3333,g3774,g4697,g4589,g3780,g6737,
    g6077,g3662,g6643,g3290,g6634,g6545,g2113,g1576,g6099,g3181,g3381,g3685,g3700,g3421,g2846,g5569,
    g5348,g4597,g6613,g6554,g4739,g2850,g6269,g4937,g4668,g4642,g4638,g3631,g2160,g4390,g3301,g4156,
    g3926,g4942,g5183,g5023,g3935,g4363,g4032,g4053,g4453,g4238,g5161,g3669,g5361,g3368,g6135,g5665,
    g6831,g4544,g6288,g4357,g3990,g5146,g6916,g5633,g6749,g6798,g4946,g6781,g5944,g5778,g5240,g5043,
    g3941,g2307,g6302,g6719,g1570,g4683,g4585,g5681,g3688,g4735,g2018,g6265,g4782,g4661,g4637,g4634,
    g4949,g3326,g6770,g6754,g3760,g5936,g4039,g5317,g3383,g5601,g3608,g3924,g4583,g3161,g2339,g3361,
    g4616,g4231,g3665,g3127,g3327,g3146,g3633,g5937,g5775,g3103,g3303,g5668,g6338,g6251,g5190,g5501,
    g5156,g5356,g5265,g5942,g4789,g3316,g5954,g5163,g6098,g3147,g5363,g3681,g5053,g4599,g3697,g5157,
    g5357,g4244,g4340,g3972,g3117,g3317,g4035,g6086,g4214,g1822,g1620,g3784,g2916,g3479,g6131,g3668,
    g6331,g3891,g4236,g3907,g3294,g5949,g3190,g6766,g3156,g3356,g5646,g2873,g1845,g6748,g5603,g5504,
    g5484,g4928,g3704,g4464,g4272,g4785,g6091,g3810,g5952,g5616,g5505,g6718,g6767,g3157,g3357,g4489,
    g2770,g5503,g3626,g4038,g5617,g3683,g4836,g3661,g6247,g3627,g5945,g2808,g2009,g3292,g3646,g2759,
    g6910,g3603,g3484,g5482,g3702,g6066,g5214,g3616,g6055,g6133,g5663,g6333,g3896,g3764,g5402,g5236,
    g4708,g5556,g5015,g3277,g3617,g6093,g2897,g6256,g6816,g4829,g6263,g4874,g3709,g5557,g5016,g3340,
    g6631,g3522,g4177,g3933,g5948,g5779,g4377,g3690,g5955,g5782,g5350,g5325,g5438,g5224,g2868,g1316,
    g3310,g4797,g5212,g3663,g2793,g2015,g4344,g3981,g5229,g6772,g3762,g4694,g1481,g4578,g3657,g2721,
    g4488,g4701,g4596,g3928,g3899,g3464,g5620,g5507,g4870,g4779,g3295,g2671,g2263,g3089,g3489,g2607,
    g5192,g5485,g5941,g5777,g4230,g3756,g6126,g6326,g3833,g4033,g2758,g3350,g6924,g6920,g6919,g5176,
    g4395,g5376,g5911,g5817,g6127,g6327,g3884,g5225,g4342,g3978,g6146,g6346,g6274,g4354,I5352,g3529,
    g3531,g3535,g3538,g5177,g6240,g4205,g3620,g1027,g2685,g2700,g6316,g3855,g5898,g5800,g4401,g1514,
    g5900,g5804,g2950,g2156,g5245,g1763,g4828,g3298,g4830,g5144,g4592,g6914,g2101,g5488,g4932,g1416,
    g5683,g6317,g3862,g5215,g4864,g5951,g5780,g4677,g4652,g4646,g3176,g3376,g3286,g3765,g4349,g6060,
    g3518,g3521,g3526,g3530,g3610,g6739,g3324,g6079,g5122,g3377,g4352,g3988,g4867,g4811,g6156,g3287,
    g5096,g4186,g3973,g5496,g5446,g6250,g4280,g3144,g3344,g5142,g3819,g6912,g6157,g5481,g3701,g5497,
    g5447,g5154,g5354,g5249,g4461,g4241,g4756,I5351,g5218,g3650,g4345,g3982,g3336,g4359,g3806,g2024,
    g3905,g3887,g3276,g3122,g2435,g2732,g4047,g6646,g3433,g905,g5953,g5781,g6084,g6603,g5677,g3195,
    g3337,g5349,g5324,g5198,g5398,g6647,g1691,g3692,g3154,g4800,g5152,g6320,g3869,g5211,g4860,g5186,
    g5599,g4490,g3293,g6771,g6758,g3329,g5170,g5091,g4456,g3829,g4348,g3987,g4355,g5939,g5776,g2294,
    g4698,g4586,g5483,g3703,g6738,g6244,g2356,g6140,g6340,g6257,g5187,g6082,g4057,g5904,g5812,g5200,
    g4457,g4261,g5241,g3349,g2053,g5145,g6915,g4834,g4686,g4590,g5191,g3699,g4598,g5637,g5159,g5359,
    g3644,g3319,g3352,g5047,g3954,g2311,g3186,g3170,g3614,g3325,g4341,g3977,g2782,g3280,g4691,g4581,
    g5935,g2949,g3511,g3517,g3520,g3525,g5234,g3636,g2292,g6089,g6731,g6717,g4427,g6557,g4358,g3991,
    g2084,g5213,g4862,g6254,g6150,g5902,g5808,g3145,g3345,g6773,g3763,g3191,g4180,g3929,g5166,g3637,
    g4832,g6769,g3307,g3359,g3757,g3315,g3642,g3654,g5619,I8376,I8393,I8394,I8395,I8377,g5659,g2100,
    g1582,g5374,g3598,I8136,g5666,I8137,g6280,I9057,I8081,I9064,I9065,I9066,g5372,I8129,I8367,I8368,
    I8369,I8370,g4243,g5202,g4000,I8349,I8345,I8346,I8347,I8348,g6703,I8119,g5674,g6747,I8211,I8386,
    g5680,g6358,I8387,g6281,I8385,I8359,g4233,g5672,g5048,I8128,I7970,I7987,I8118,g1589,I8358,g6659,
    g6073,g6741,g6929,g3992,g5678,g2080,I7980,I8360,I8356,I8357,I8379,g6357,g5066,I8209,g5662,I7972,
    I9059,g6279,g5669,g5368,I7979,g4936,g6926,I8378,I8135,g3012,g6400,g6927,g6660,I8208,g3028,I8138,
    I9058,g5060,g4819,I7978,I7989,I7971,g3215,I8774,g3503,I7969,g4941,I7988,I8080,g6669,I8126,g5062,
    g6359,I8779,I7981,I8127,I8778,I8210,g5377,I8117,I8079,g6335,g5065,g2995,g2095,g1573,g6683,g5676,
    I8773,g4432,g5068,I7990,I8120,g2067,g4234,g5227,I8082,g5370,g3013,g6740,g6928,g2951,g6705,g6075,
    g5367,I7217,I7216,I7571,I7569,I2073,I2072,I2796,I2795,g948,I2014,I2015,I4205,I4203,I3875,I3874,
    g3109,I5536,I5537,I5658,g3983,I5657,I2527,I2528,I4444,I5271,I5269,I2898,I2897,I2797,I2245,I2244,
    I3988,I2543,I2544,I1963,I1961,I5209,I5207,I7562,I7231,I7232,I6744,I6745,I4182,I6186,g4301,I6185,
    I7441,I7439,I6026,g4223,g4221,I2768,I2766,I3933,g2731,I3894,I3895,I7238,I7239,I4160,I4161,I2934,
    I2933,I3179,I3177,I6187,g3955,I6027,I4233,g2769,I3953,I3954,g1044,I2081,I2082,g4674,I6391,g4504,
    I6390,g4680,I2080,I8195,I8194,g1534,I2498,I2499,I2497,g1042,g1036,g939,I1987,I1988,I2061,I2062,
    I2676,I2674,I2767,I7528,I7529,I7434,I7432,I2074,I7210,I7208,I6964,I6962,I5208,I5302,I5300,I7535,
    I7536,I6195,I6196,I2542,I1994,I4445,I2060,I5189,I5187,I3178,I4920,I4919,I2003,I3916,I3914,I5309,
    I5307,I5759,I6659,g4762,I4940,I4939,I2935,I3412,I3413,I3411,I3189,I3188,I3990,I4151,I4152,I2090,
    I2089,g5862,I9050,I5766,g3961,g3957,g3968,I5227,I5228,I7527,I5226,g4049,I7224,I7223,I5767,I5535,
    g2944,I4921,I6028,I7244,I5188,I5270,I9051,I9052,I5308,I2506,g1047,I3445,I3169,I3170,g1540,I3168,
    I7556,I7555,I5196,I5195,I7563,I7440,I2507,I1995,I3446,I3447,I7237,g2757,I3934,I3935,I6743,I4183,
    I7557,I2300,I2299,I5197,I4159,I3741,I3739,I6660,I6661,I5257,I2526,I5301,I4204,I7218,I6175,I3455,
    I6500,I6499,I3846,I4210,I6474,I6475,g2698,I3847,I3848,g1518,I7520,I4784,I4782,I1952,I1951,I8202,
    I8201,I1986,I5760,I5768,I1970,I1969,I7225,I7209,I2301,I7245,I3740,I6963,I3456,I3457,I3126,I3125,
    I3400,I3398,I4526,I4527,I4528,g2795,I6176,I6177,I7230,I7433,I3127,I4234,I4235,I5784,I5782,I7550,
    I7548,I4546,I4545,I5294,I5292,g937,I1979,I1980,g4472,g1473,g1470,g1459,g928,I1962,I7097,I4547,
    I3697,I7312,I7311,I2109,I2110,I2013,g2804,I4009,I4010,g5863,I2022,I2021,I7576,g5688,I3190,I3952,
    I7549,I7577,I5647,g3974,I1978,I7246,I4150,g3621,I4008,I2675,g926,I1953,I3893,I4212,I7313,I2108,
    I5244,I5242,I7534,I7522,I7521,I6194,I3970,I4941,g3979,I7542,I7541,I2682,I2681,I4211,I3876,I2091,
    I3915,I4783,I7543,g930,I1971,I7570,I5293,I2246,I6392,g944,I2004,I2005,I6473,g2719,I8203,I2899,
    g941,I1996,I2508,g2745,g2791,I3989,I8196,I5259,g1560,g4610,I6501,I3399,I3698,I3699,g950,I2023,
    I4446,I5783,g2940,I5761,I3972,I7098,I7099,g2780,I3971,I5258,I7564,I5648,I5649,I5243,I2683,I7578,
    I5659,I4184,g3528,g3664,g3656,g3647,g1449,g1418,g1879,extra0,extra1,extra2,extra3,extra4,extra5,extra6,
    extra7,extra8,extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,extra17,extra18,extra19,extra20,extra21,extra22,
    extra23,extra24;

  DFF_X2 DFF_0( .CK(CK), .Q(g678), .D(g4130) );
  DFF_X2 DFF_1( .CK(CK), .Q(g332), .D(g6823) );
  DFF_X2 DFF_2( .CK(CK), .Q(g123), .D(g6940) );
  DFF_X1 DFF_3( .CK(CK), .Q(g207), .D(g6102) );
  DFF_X1 DFF_4( .CK(CK), .Q(g695), .D(g4147) );
  DFF_X1 DFF_5( .CK(CK), .Q(g461), .D(g4841) );
  DFF_X1 DFF_6( .CK(CK), .Q(g18), .D(g6725) );
  DFF_X1 DFF_7( .CK(CK), .Q(g292), .D(g3232) );
  DFF_X1 DFF_8( .CK(CK), .Q(g331), .D(g4119) );
  DFF_X1 DFF_9( .CK(CK), .Q(g689), .D(g4141) );
  DFF_X1 DFF_10( .CK(CK), .Q(g24), .D(g6726) );
  DFF_X1 DFF_11( .CK(CK), .Q(g465), .D(g6507) );
  DFF_X1 DFF_12( .CK(CK), .Q(g84), .D(g6590) );
  DFF_X1 DFF_13( .CK(CK), .Q(g291), .D(g3231) );
  DFF_X1 DFF_14( .CK(CK), .Q(g676), .D(g5330) );
  DFF_X1 DFF_15( .CK(CK), .Q(g622), .D(g5147) );
  DFF_X1 DFF_16( .CK(CK), .Q(g117), .D(g4839) );
  DFF_X1 DFF_17( .CK(CK), .Q(g278), .D(g6105) );
  DFF_X1 DFF_18( .CK(CK), .Q(g128), .D(g5138) );
  DFF_X1 DFF_19( .CK(CK), .Q(g598), .D(g4122) );
  DFF_X1 DFF_20( .CK(CK), .Q(g554), .D(g6827) );
  DFF_X1 DFF_21( .CK(CK), .Q(g496), .D(g6745) );
  DFF_X1 DFF_22( .CK(CK), .Q(g179), .D(g6405) );
  DFF_X1 DFF_23( .CK(CK), .Q(g48), .D(g6729) );
  DFF_X1 DFF_24( .CK(CK), .Q(g590), .D(g6595) );
  DFF_X1 DFF_25( .CK(CK), .Q(g551), .D(g6826) );
  DFF_X1 DFF_26( .CK(CK), .Q(g682), .D(g4134) );
  DFF_X1 DFF_27( .CK(CK), .Q(g11), .D(g6599) );
  DFF_X1 DFF_28( .CK(CK), .Q(g606), .D(g4857) );
  DFF_X1 DFF_29( .CK(CK), .Q(g188), .D(g6406) );
  DFF_X1 DFF_30( .CK(CK), .Q(g646), .D(g5148) );
  DFF_X1 DFF_31( .CK(CK), .Q(g327), .D(g4117) );
  DFF_X1 DFF_32( .CK(CK), .Q(g361), .D(g6582) );
  DFF_X1 DFF_33( .CK(CK), .Q(g289), .D(g3229) );
  DFF_X1 DFF_34( .CK(CK), .Q(g398), .D(g5700) );
  DFF_X1 DFF_35( .CK(CK), .Q(g684), .D(g4136) );
  DFF_X1 DFF_36( .CK(CK), .Q(g619), .D(g4858) );
  DFF_X1 DFF_37( .CK(CK), .Q(g208), .D(g5876) );
  DFF_X1 DFF_38( .CK(CK), .Q(g248), .D(g3239) );
  DFF_X1 DFF_39( .CK(CK), .Q(g390), .D(g5698) );
  DFF_X1 DFF_40( .CK(CK), .Q(g625), .D(g5328) );
  DFF_X1 DFF_41( .CK(CK), .Q(g681), .D(g4133) );
  DFF_X1 DFF_42( .CK(CK), .Q(g437), .D(g4847) );
  DFF_X1 DFF_43( .CK(CK), .Q(g276), .D(g5877) );
  DFF_X1 DFF_44( .CK(CK), .Q(g3), .D(g6597) );
  DFF_X1 DFF_45( .CK(CK), .Q(g323), .D(g4120) );
  DFF_X1 DFF_46( .CK(CK), .Q(g224), .D(g3235) );
  DFF_X1 DFF_47( .CK(CK), .Q(g685), .D(g4137) );
  DFF_X1 DFF_48( .CK(CK), .Q(g43), .D(g6407) );
  DFF_X1 DFF_49( .CK(CK), .Q(g157), .D(g5470) );
  DFF_X1 DFF_50( .CK(CK), .Q(g282), .D(g6841) );
  DFF_X1 DFF_51( .CK(CK), .Q(g697), .D(g4149) );
  DFF_X1 DFF_52( .CK(CK), .Q(g206), .D(g6101) );
  DFF_X1 DFF_53( .CK(CK), .Q(g449), .D(g4844) );
  DFF_X1 DFF_54( .CK(CK), .Q(g118), .D(g4113) );
  DFF_X1 DFF_55( .CK(CK), .Q(g528), .D(g6504) );
  DFF_X1 DFF_56( .CK(CK), .Q(g284), .D(g3224) );
  DFF_X1 DFF_57( .CK(CK), .Q(g426), .D(g4855) );
  DFF_X1 DFF_58( .CK(CK), .Q(g634), .D(g4424) );
  DFF_X1 DFF_59( .CK(CK), .Q(g669), .D(g5582) );
  DFF_X1 DFF_60( .CK(CK), .Q(g520), .D(g6502) );
  DFF_X1 DFF_61( .CK(CK), .Q(g281), .D(g6107) );
  DFF_X1 DFF_62( .CK(CK), .Q(g175), .D(g5472) );
  DFF_X1 DFF_63( .CK(CK), .Q(g15), .D(g6602) );
  DFF_X1 DFF_64( .CK(CK), .Q(g631), .D(g5581) );
  DFF_X1 DFF_65( .CK(CK), .Q(g69), .D(g6587) );
  DFF_X1 DFF_66( .CK(CK), .Q(g693), .D(g4145) );
  DFF_X1 DFF_67( .CK(CK), .Q(g337), .D(g2585) );
  DFF_X1 DFF_68( .CK(CK), .Q(g457), .D(g4842) );
  DFF_X1 DFF_69( .CK(CK), .Q(g486), .D(g2586) );
  DFF_X1 DFF_70( .CK(CK), .Q(g471), .D(g1291) );
  DFF_X1 DFF_71( .CK(CK), .Q(g328), .D(g4118) );
  DFF_X1 DFF_72( .CK(CK), .Q(g285), .D(g3225) );
  DFF_X1 DFF_73( .CK(CK), .Q(g418), .D(g4853) );
  DFF_X1 DFF_74( .CK(CK), .Q(g402), .D(g4849) );
  DFF_X2 DFF_75( .CK(CK), .Q(g297), .D(g6512) );
  DFF_X2 DFF_76( .CK(CK), .Q(g212), .D(g3233) );
  DFF_X2 DFF_77( .CK(CK), .Q(g410), .D(g4851) );
  DFF_X1 DFF_78( .CK(CK), .Q(g430), .D(g4856) );
  DFF_X1 DFF_79( .CK(CK), .Q(g33), .D(g6854) );
  DFF_X1 DFF_80( .CK(CK), .Q(g662), .D(g1831) );
  DFF_X1 DFF_81( .CK(CK), .Q(g453), .D(g4843) );
  DFF_X1 DFF_82( .CK(CK), .Q(g269), .D(g6510) );
  DFF_X1 DFF_83( .CK(CK), .Q(g574), .D(g6591) );
  DFF_X1 DFF_84( .CK(CK), .Q(g441), .D(g4846) );
  DFF_X1 DFF_85( .CK(CK), .Q(g664), .D(g1288) );
  DFF_X1 DFF_86( .CK(CK), .Q(g349), .D(g5478) );
  DFF_X1 DFF_87( .CK(CK), .Q(g211), .D(g6840) );
  DFF_X1 DFF_88( .CK(CK), .Q(g586), .D(g6594) );
  DFF_X1 DFF_89( .CK(CK), .Q(g571), .D(g5580) );
  DFF_X1 DFF_90( .CK(CK), .Q(g29), .D(g6853) );
  DFF_X1 DFF_91( .CK(CK), .Q(g326), .D(g4840) );
  DFF_X1 DFF_92( .CK(CK), .Q(g698), .D(g4150) );
  DFF_X1 DFF_93( .CK(CK), .Q(g654), .D(g5490) );
  DFF_X1 DFF_94( .CK(CK), .Q(g293), .D(g6511) );
  DFF_X1 DFF_95( .CK(CK), .Q(g690), .D(g4142) );
  DFF_X1 DFF_96( .CK(CK), .Q(g445), .D(g4845) );
  DFF_X1 DFF_97( .CK(CK), .Q(g374), .D(g5694) );
  DFF_X1 DFF_98( .CK(CK), .Q(g6), .D(g6722) );
  DFF_X1 DFF_99( .CK(CK), .Q(g687), .D(g4139) );
  DFF_X1 DFF_100( .CK(CK), .Q(g357), .D(g5480) );
  DFF_X1 DFF_101( .CK(CK), .Q(g386), .D(g5697) );
  DFF_X1 DFF_102( .CK(CK), .Q(g504), .D(g6498) );
  DFF_X1 DFF_103( .CK(CK), .Q(g665), .D(g4126) );
  DFF_X1 DFF_104( .CK(CK), .Q(g166), .D(g5471) );
  DFF_X1 DFF_105( .CK(CK), .Q(g541), .D(g6505) );
  DFF_X1 DFF_106( .CK(CK), .Q(g74), .D(g6588) );
  DFF_X1 DFF_107( .CK(CK), .Q(g338), .D(g5475) );
  DFF_X1 DFF_108( .CK(CK), .Q(g696), .D(g4148) );
  DFF_X1 DFF_109( .CK(CK), .Q(g516), .D(g6501) );
  DFF_X1 DFF_110( .CK(CK), .Q(g536), .D(g6506) );
  DFF_X1 DFF_111( .CK(CK), .Q(g683), .D(g4135) );
  DFF_X1 DFF_112( .CK(CK), .Q(g353), .D(g5479) );
  DFF_X1 DFF_113( .CK(CK), .Q(g545), .D(g6824) );
  DFF_X1 DFF_114( .CK(CK), .Q(g254), .D(g3240) );
  DFF_X1 DFF_115( .CK(CK), .Q(g341), .D(g5476) );
  DFF_X1 DFF_116( .CK(CK), .Q(g290), .D(g3230) );
  DFF_X1 DFF_117( .CK(CK), .Q(g2), .D(g6721) );
  DFF_X1 DFF_118( .CK(CK), .Q(g287), .D(g3227) );
  DFF_X1 DFF_119( .CK(CK), .Q(g336), .D(g6925) );
  DFF_X1 DFF_120( .CK(CK), .Q(g345), .D(g5477) );
  DFF_X1 DFF_121( .CK(CK), .Q(g628), .D(g5489) );
  DFF_X1 DFF_122( .CK(CK), .Q(g679), .D(g4131) );
  DFF_X1 DFF_123( .CK(CK), .Q(g28), .D(g6727) );
  DFF_X1 DFF_124( .CK(CK), .Q(g688), .D(g4140) );
  DFF_X1 DFF_125( .CK(CK), .Q(g283), .D(g6842) );
  DFF_X1 DFF_126( .CK(CK), .Q(g613), .D(g4423) );
  DFF_X1 DFF_127( .CK(CK), .Q(g10), .D(g6723) );
  DFF_X1 DFF_128( .CK(CK), .Q(g14), .D(g6724) );
  DFF_X1 DFF_129( .CK(CK), .Q(g680), .D(g4132) );
  DFF_X1 DFF_130( .CK(CK), .Q(g143), .D(g6401) );
  DFF_X1 DFF_131( .CK(CK), .Q(g672), .D(g5491) );
  DFF_X1 DFF_132( .CK(CK), .Q(g667), .D(g4127) );
  DFF_X1 DFF_133( .CK(CK), .Q(g366), .D(g6278) );
  DFF_X1 DFF_134( .CK(CK), .Q(g279), .D(g6106) );
  DFF_X1 DFF_135( .CK(CK), .Q(g492), .D(g6744) );
  DFF_X1 DFF_136( .CK(CK), .Q(g170), .D(g6404) );
  DFF_X1 DFF_137( .CK(CK), .Q(g686), .D(g4138) );
  DFF_X1 DFF_138( .CK(CK), .Q(g288), .D(g3228) );
  DFF_X1 DFF_139( .CK(CK), .Q(g638), .D(g1289) );
  DFF_X1 DFF_140( .CK(CK), .Q(g602), .D(g4123) );
  DFF_X1 DFF_141( .CK(CK), .Q(g642), .D(g4658) );
  DFF_X1 DFF_142( .CK(CK), .Q(g280), .D(g5878) );
  DFF_X1 DFF_143( .CK(CK), .Q(g663), .D(g4125) );
  DFF_X1 DFF_144( .CK(CK), .Q(g610), .D(g4124) );
  DFF_X1 DFF_145( .CK(CK), .Q(g148), .D(g5874) );
  DFF_X1 DFF_146( .CK(CK), .Q(g209), .D(g6103) );
  DFF_X1 DFF_147( .CK(CK), .Q(g675), .D(g1294) );
  DFF_X1 DFF_148( .CK(CK), .Q(g478), .D(g1292) );
  DFF_X1 DFF_149( .CK(CK), .Q(g122), .D(g4115) );
  DFF_X1 DFF_150( .CK(CK), .Q(g54), .D(g6584) );
  DFF_X1 DFF_151( .CK(CK), .Q(g594), .D(g6596) );
  DFF_X1 DFF_152( .CK(CK), .Q(g286), .D(g3226) );
  DFF_X1 DFF_153( .CK(CK), .Q(g489), .D(g2587) );
  DFF_X1 DFF_154( .CK(CK), .Q(g616), .D(g4657) );
  DFF_X1 DFF_155( .CK(CK), .Q(g79), .D(g6589) );
  DFF_X1 DFF_156( .CK(CK), .Q(g218), .D(g3234) );
  DFF_X1 DFF_157( .CK(CK), .Q(g242), .D(g3238) );
  DFF_X1 DFF_158( .CK(CK), .Q(g578), .D(g6592) );
  DFF_X1 DFF_159( .CK(CK), .Q(g184), .D(g5473) );
  DFF_X1 DFF_160( .CK(CK), .Q(g119), .D(g4114) );
  DFF_X1 DFF_161( .CK(CK), .Q(g668), .D(g6800) );
  DFF_X1 DFF_162( .CK(CK), .Q(g139), .D(g5141) );
  DFF_X1 DFF_163( .CK(CK), .Q(g422), .D(g4854) );
  DFF_X1 DFF_164( .CK(CK), .Q(g210), .D(g6839) );
  DFF_X1 DFF_165( .CK(CK), .Q(g394), .D(g5699) );
  DFF_X1 DFF_166( .CK(CK), .Q(g230), .D(g3236) );
  DFF_X1 DFF_167( .CK(CK), .Q(g25), .D(g6601) );
  DFF_X1 DFF_168( .CK(CK), .Q(g204), .D(g5875) );
  DFF_X1 DFF_169( .CK(CK), .Q(g658), .D(g4425) );
  DFF_X1 DFF_170( .CK(CK), .Q(g650), .D(g5329) );
  DFF_X1 DFF_171( .CK(CK), .Q(g378), .D(g5695) );
  DFF_X1 DFF_172( .CK(CK), .Q(g508), .D(g6499) );
  DFF_X1 DFF_173( .CK(CK), .Q(g548), .D(g6825) );
  DFF_X1 DFF_174( .CK(CK), .Q(g370), .D(g5693) );
  DFF_X1 DFF_175( .CK(CK), .Q(g406), .D(g4850) );
  DFF_X1 DFF_176( .CK(CK), .Q(g236), .D(g3237) );
  DFF_X1 DFF_177( .CK(CK), .Q(g500), .D(g6497) );
  DFF_X1 DFF_178( .CK(CK), .Q(g205), .D(g6100) );
  DFF_X1 DFF_179( .CK(CK), .Q(g197), .D(g6509) );
  DFF_X1 DFF_180( .CK(CK), .Q(g666), .D(g4128) );
  DFF_X1 DFF_181( .CK(CK), .Q(g114), .D(g4116) );
  DFF_X1 DFF_182( .CK(CK), .Q(g524), .D(g6503) );
  DFF_X1 DFF_183( .CK(CK), .Q(g260), .D(g3241) );
  DFF_X1 DFF_184( .CK(CK), .Q(g111), .D(g6277) );
  DFF_X1 DFF_185( .CK(CK), .Q(g131), .D(g5139) );
  DFF_X1 DFF_186( .CK(CK), .Q(g7), .D(g6598) );
  DFF_X1 DFF_187( .CK(CK), .Q(g19), .D(g6600) );
  DFF_X2 DFF_188( .CK(CK), .Q(g677), .D(g4129) );
  DFF_X2 DFF_189( .CK(CK), .Q(g582), .D(g6593) );
  DFF_X2 DFF_190( .CK(CK), .Q(g485), .D(g6801) );
  DFF_X2 DFF_191( .CK(CK), .Q(g699), .D(g4426) );
  DFF_X2 DFF_192( .CK(CK), .Q(g193), .D(g5474) );
  DFF_X2 DFF_193( .CK(CK), .Q(g135), .D(g5140) );
  DFF_X2 DFF_194( .CK(CK), .Q(g382), .D(g5696) );
  DFF_X1 DFF_195( .CK(CK), .Q(g414), .D(g4852) );
  DFF_X1 DFF_196( .CK(CK), .Q(g434), .D(g4848) );
  DFF_X1 DFF_197( .CK(CK), .Q(g266), .D(g4659) );
  DFF_X1 DFF_198( .CK(CK), .Q(g49), .D(g6583) );
  DFF_X1 DFF_199( .CK(CK), .Q(g152), .D(g6402) );
  DFF_X1 DFF_200( .CK(CK), .Q(g692), .D(g4144) );
  DFF_X1 DFF_201( .CK(CK), .Q(g277), .D(g6104) );
  DFF_X1 DFF_202( .CK(CK), .Q(g127), .D(g6941) );
  DFF_X1 DFF_203( .CK(CK), .Q(g161), .D(g6403) );
  DFF_X1 DFF_204( .CK(CK), .Q(g512), .D(g6500) );
  DFF_X1 DFF_205( .CK(CK), .Q(g532), .D(g6508) );
  DFF_X1 DFF_206( .CK(CK), .Q(g64), .D(g6586) );
  DFF_X1 DFF_207( .CK(CK), .Q(g694), .D(g4146) );
  DFF_X1 DFF_208( .CK(CK), .Q(g691), .D(g4143) );
  DFF_X1 DFF_209( .CK(CK), .Q(g1), .D(g6720) );
  DFF_X1 DFF_210( .CK(CK), .Q(g59), .D(g6585) );
  INV_X1 NOT_0( .ZN(I8854), .A(g6696) );
  INV_X1 NOT_1( .ZN(g1289), .A(I2272) );
  INV_X1 NOT_2( .ZN(I9125), .A(g6855) );
  INV_X1 NOT_3( .ZN(I6783), .A(g4822) );
  INV_X1 NOT_4( .ZN(I4424), .A(g2097) );
  INV_X1 NOT_5( .ZN(g6895), .A(I9152) );
  INV_X1 NOT_6( .ZN(g1835), .A(I2919) );
  INV_X1 NOT_7( .ZN(I3040), .A(g1770) );
  INV_X1 NOT_8( .ZN(g6837), .A(g6822) );
  INV_X1 NOT_9( .ZN(I7466), .A(g5624) );
  INV_X1 NOT_10( .ZN(I4809), .A(g2974) );
  INV_X1 NOT_11( .ZN(g3537), .A(I4757) );
  INV_X1 NOT_12( .ZN(g5457), .A(g5304) );
  INV_X1 NOT_13( .ZN(g6062), .A(g5824) );
  INV_X1 NOT_14( .ZN(g4040), .A(I5343) );
  INV_X1 NOT_15( .ZN(I6001), .A(g4162) );
  INV_X1 NOT_16( .ZN(g5549), .A(g5331) );
  INV_X1 NOT_17( .ZN(I4477), .A(g3063) );
  INV_X1 NOT_18( .ZN(g3612), .A(I4809) );
  INV_X1 NOT_19( .ZN(I7055), .A(g5318) );
  INV_X1 NOT_20( .ZN(g2892), .A(g1982) );
  INV_X1 NOT_21( .ZN(I5264), .A(g3638) );
  INV_X1 NOT_22( .ZN(I2225), .A(g696) );
  INV_X1 NOT_23( .ZN(g4123), .A(I5451) );
  INV_X1 NOT_24( .ZN(g4323), .A(g4086) );
  INV_X1 NOT_25( .ZN(g908), .A(I1932) );
  INV_X1 NOT_26( .ZN(I5933), .A(g4346) );
  INV_X1 NOT_27( .ZN(I8252), .A(g6294) );
  INV_X1 NOT_28( .ZN(I2473), .A(g971) );
  INV_X1 NOT_29( .ZN(I7333), .A(g5386) );
  INV_X1 NOT_30( .ZN(I8812), .A(g6688) );
  INV_X1 NOT_31( .ZN(g1674), .A(g985) );
  INV_X1 NOT_32( .ZN(I3528), .A(g1422) );
  INV_X1 NOT_33( .ZN(I8958), .A(g6774) );
  INV_X1 NOT_34( .ZN(I5050), .A(g3246) );
  INV_X1 NOT_35( .ZN(g3234), .A(I4501) );
  INV_X1 NOT_36( .ZN(I2324), .A(g1209) );
  INV_X1 NOT_37( .ZN(g2945), .A(I4133) );
  INV_X1 NOT_38( .ZN(g5121), .A(I6775) );
  INV_X1 NOT_39( .ZN(g1997), .A(g1398) );
  INV_X1 NOT_40( .ZN(g3128), .A(I4375) );
  INV_X1 NOT_41( .ZN(I8005), .A(g6110) );
  INV_X1 NOT_42( .ZN(g1541), .A(g1094) );
  INV_X1 NOT_43( .ZN(g5670), .A(g5527) );
  INV_X1 NOT_44( .ZN(g2738), .A(g2327) );
  INV_X8 NOT_45( .ZN(g6842), .A(I9047) );
  INV_X8 NOT_46( .ZN(g4528), .A(I6096) );
  INV_X8 NOT_47( .ZN(g2244), .A(I3379) );
  INV_X8 NOT_48( .ZN(g6192), .A(g5946) );
  INV_X1 NOT_49( .ZN(g2709), .A(I3864) );
  INV_X1 NOT_50( .ZN(g1332), .A(I2349) );
  INV_X1 NOT_51( .ZN(g4530), .A(I6102) );
  INV_X1 NOT_52( .ZN(g1680), .A(g1011) );
  INV_X1 NOT_53( .ZN(g2078), .A(g1345) );
  INV_X1 NOT_54( .ZN(g1209), .A(I2215) );
  INV_X1 NOT_55( .ZN(I3010), .A(g1504) );
  INV_X1 NOT_56( .ZN(g5813), .A(I7612) );
  INV_X1 NOT_57( .ZN(I7509), .A(g5587) );
  INV_X1 NOT_58( .ZN(I5379), .A(g3940) );
  INV_X1 NOT_59( .ZN(g3800), .A(g3388) );
  INV_X1 NOT_60( .ZN(g2907), .A(g1914) );
  INV_X1 NOT_61( .ZN(g6854), .A(I9085) );
  INV_X1 NOT_62( .ZN(g2035), .A(I3144) );
  INV_X1 NOT_63( .ZN(g2959), .A(g1861) );
  INV_X1 NOT_64( .ZN(g6941), .A(I9236) );
  INV_X1 NOT_65( .ZN(g4010), .A(g3601) );
  INV_X1 NOT_66( .ZN(I2287), .A(g927) );
  INV_X1 NOT_67( .ZN(I4273), .A(g2197) );
  INV_X1 NOT_68( .ZN(I8270), .A(g6300) );
  INV_X1 NOT_69( .ZN(g5740), .A(I7501) );
  INV_X1 NOT_70( .ZN(I5777), .A(g3807) );
  INV_X1 NOT_71( .ZN(g2876), .A(g1943) );
  INV_X1 NOT_72( .ZN(g873), .A(g306) );
  INV_X1 NOT_73( .ZN(g4839), .A(I6525) );
  INV_X1 NOT_74( .ZN(I5882), .A(g3871) );
  INV_X1 NOT_75( .ZN(g2656), .A(I3800) );
  INV_X1 NOT_76( .ZN(I8473), .A(g6485) );
  INV_X1 NOT_77( .ZN(I2199), .A(g33) );
  INV_X1 NOT_78( .ZN(g900), .A(I1927) );
  INV_X1 NOT_79( .ZN(g6708), .A(I8834) );
  INV_X1 NOT_80( .ZN(I2399), .A(g729) );
  INV_X1 NOT_81( .ZN(I3278), .A(g1695) );
  INV_X1 NOT_82( .ZN(g6520), .A(I8476) );
  INV_X1 NOT_83( .ZN(g940), .A(g64) );
  INV_X1 NOT_84( .ZN(I6677), .A(g4757) );
  INV_X1 NOT_85( .ZN(g3902), .A(g3575) );
  INV_X1 NOT_86( .ZN(g5687), .A(g5567) );
  INV_X1 NOT_87( .ZN(g2915), .A(g1931) );
  INV_X1 NOT_88( .ZN(g847), .A(g590) );
  INV_X1 NOT_89( .ZN(I3235), .A(g1807) );
  INV_X1 NOT_90( .ZN(I3343), .A(g1623) );
  INV_X1 NOT_91( .ZN(g6431), .A(I8295) );
  INV_X4 NOT_92( .ZN(g709), .A(g114) );
  INV_X4 NOT_93( .ZN(g6812), .A(I8984) );
  INV_X1 NOT_94( .ZN(I6576), .A(g4700) );
  INV_X1 NOT_95( .ZN(g749), .A(I1847) );
  INV_X1 NOT_96( .ZN(g3090), .A(I4331) );
  INV_X1 NOT_97( .ZN(I9107), .A(g6855) );
  INV_X1 NOT_98( .ZN(g2214), .A(I3349) );
  INV_X1 NOT_99( .ZN(g4618), .A(g4246) );
  INV_X1 NOT_100( .ZN(g6376), .A(g6267) );
  INV_X1 NOT_101( .ZN(g4143), .A(I5511) );
  INV_X1 NOT_102( .ZN(I6349), .A(g4569) );
  INV_X1 NOT_103( .ZN(g4343), .A(g4011) );
  INV_X1 NOT_104( .ZN(I5674), .A(g4003) );
  INV_X1 NOT_105( .ZN(I8177), .A(g6173) );
  INV_X1 NOT_106( .ZN(g2110), .A(g1381) );
  INV_X1 NOT_107( .ZN(I3134), .A(g1336) );
  INV_X1 NOT_108( .ZN(g6405), .A(I8229) );
  INV_X1 NOT_109( .ZN(I3334), .A(g1330) );
  INV_X1 NOT_110( .ZN(I7197), .A(g5431) );
  INV_X1 NOT_111( .ZN(g4566), .A(g4198) );
  INV_X1 NOT_112( .ZN(I7397), .A(g5561) );
  INV_X1 NOT_113( .ZN(I4534), .A(g2858) );
  INV_X1 NOT_114( .ZN(g1714), .A(g1110) );
  INV_X2 NOT_115( .ZN(I4961), .A(g3597) );
  INV_X2 NOT_116( .ZN(g2663), .A(g2308) );
  INV_X2 NOT_117( .ZN(g3456), .A(g2640) );
  INV_X1 NOT_118( .ZN(g5141), .A(I6801) );
  INV_X1 NOT_119( .ZN(g922), .A(I1947) );
  INV_X1 NOT_120( .ZN(g4693), .A(I6283) );
  INV_X1 NOT_121( .ZN(g4134), .A(I5484) );
  INV_X1 NOT_122( .ZN(g5570), .A(g5392) );
  INV_X1 NOT_123( .ZN(g5860), .A(g5634) );
  INV_X1 NOT_124( .ZN(g4334), .A(g3733) );
  INV_X1 NOT_125( .ZN(I3804), .A(g2575) );
  INV_X1 NOT_126( .ZN(I2207), .A(g7) );
  INV_X1 NOT_127( .ZN(I5153), .A(g3330) );
  INV_X1 NOT_128( .ZN(g3355), .A(g3100) );
  INV_X1 NOT_129( .ZN(g5645), .A(g5537) );
  INV_X1 NOT_130( .ZN(g6733), .A(I8891) );
  INV_X1 NOT_131( .ZN(g5691), .A(g5568) );
  INV_X1 NOT_132( .ZN(g4804), .A(g4473) );
  INV_X1 NOT_133( .ZN(I9047), .A(g6838) );
  INV_X1 NOT_134( .ZN(I4414), .A(g2090) );
  INV_X1 NOT_135( .ZN(g6610), .A(I8696) );
  INV_X1 NOT_136( .ZN(g2877), .A(g2434) );
  INV_X1 NOT_137( .ZN(I4903), .A(g3223) );
  INV_X1 NOT_138( .ZN(g6796), .A(I8958) );
  INV_X1 NOT_139( .ZN(g3063), .A(I4288) );
  INV_X1 NOT_140( .ZN(I3313), .A(g1337) );
  INV_X1 NOT_141( .ZN(g5879), .A(g5770) );
  INV_X1 NOT_142( .ZN(g3463), .A(g2682) );
  INV_X1 NOT_143( .ZN(I4513), .A(g2765) );
  INV_X1 NOT_144( .ZN(g1623), .A(I2578) );
  INV_X1 NOT_145( .ZN(g5358), .A(I7012) );
  INV_X1 NOT_146( .ZN(I3202), .A(g1812) );
  INV_X1 NOT_147( .ZN(I2215), .A(g695) );
  INV_X1 NOT_148( .ZN(g4113), .A(I5421) );
  INV_X1 NOT_149( .ZN(g1076), .A(I2115) );
  INV_X1 NOT_150( .ZN(g6069), .A(g5791) );
  INV_X1 NOT_151( .ZN(I7817), .A(g5924) );
  INV_X1 NOT_152( .ZN(g6540), .A(g6474) );
  INV_X1 NOT_153( .ZN(I6352), .A(g4564) );
  INV_X1 NOT_154( .ZN(I1865), .A(g279) );
  INV_X1 NOT_155( .ZN(g4202), .A(I5622) );
  INV_X1 NOT_156( .ZN(I6867), .A(g5082) );
  INV_X1 NOT_157( .ZN(I5511), .A(g3876) );
  INV_X2 NOT_158( .ZN(g5587), .A(I7349) );
  INV_X2 NOT_159( .ZN(I8144), .A(g6182) );
  INV_X2 NOT_160( .ZN(g1175), .A(g42) );
  INV_X1 NOT_161( .ZN(g1375), .A(I2411) );
  INV_X1 NOT_162( .ZN(g3118), .A(I4366) );
  INV_X1 NOT_163( .ZN(g3318), .A(I4593) );
  INV_X1 NOT_164( .ZN(g2464), .A(I3596) );
  INV_X1 NOT_165( .ZN(g3872), .A(g3312) );
  INV_X1 NOT_166( .ZN(g4494), .A(I6004) );
  INV_X1 NOT_167( .ZN(I2870), .A(g1161) );
  INV_X1 NOT_168( .ZN(g4518), .A(I6066) );
  INV_X1 NOT_169( .ZN(I4288), .A(g2215) );
  INV_X1 NOT_170( .ZN(g5615), .A(I7372) );
  INV_X1 NOT_171( .ZN(g4567), .A(I6139) );
  INV_X1 NOT_172( .ZN(I4382), .A(g2265) );
  INV_X1 NOT_173( .ZN(I3776), .A(g2044) );
  INV_X1 NOT_174( .ZN(g3057), .A(I4282) );
  INV_X1 NOT_175( .ZN(I5600), .A(g3821) );
  INV_X1 NOT_176( .ZN(I3593), .A(g1295) );
  INV_X1 NOT_177( .ZN(I2825), .A(g1143) );
  INV_X1 NOT_178( .ZN(g1285), .A(g852) );
  INV_X1 NOT_179( .ZN(g3457), .A(g2653) );
  INV_X2 NOT_180( .ZN(g5174), .A(g5099) );
  INV_X2 NOT_181( .ZN(I6386), .A(g4462) );
  INV_X1 NOT_182( .ZN(I3965), .A(g2268) );
  INV_X1 NOT_183( .ZN(I8488), .A(g6426) );
  INV_X1 NOT_184( .ZN(g6849), .A(I9074) );
  INV_X1 NOT_185( .ZN(I6599), .A(g4823) );
  INV_X1 NOT_186( .ZN(I2408), .A(g719) );
  INV_X1 NOT_187( .ZN(g3834), .A(I5027) );
  INV_X1 NOT_188( .ZN(g2295), .A(g1578) );
  INV_X1 NOT_189( .ZN(g1384), .A(I2420) );
  INV_X1 NOT_190( .ZN(g1339), .A(I2370) );
  INV_X1 NOT_191( .ZN(g5545), .A(g5331) );
  INV_X1 NOT_192( .ZN(I6170), .A(g4343) );
  INV_X1 NOT_193( .ZN(I9128), .A(g6864) );
  INV_X1 NOT_194( .ZN(g6898), .A(I9161) );
  INV_X1 NOT_195( .ZN(g1838), .A(g1595) );
  INV_X1 NOT_196( .ZN(g6900), .A(I9167) );
  INV_X1 NOT_197( .ZN(g2194), .A(I3331) );
  INV_X1 NOT_198( .ZN(g6797), .A(I8961) );
  INV_X1 NOT_199( .ZN(g2394), .A(I3537) );
  INV_X1 NOT_200( .ZN(I3050), .A(g1439) );
  INV_X1 NOT_201( .ZN(I3641), .A(g1491) );
  INV_X1 NOT_202( .ZN(I2943), .A(g1715) );
  INV_X1 NOT_203( .ZN(I5736), .A(g4022) );
  INV_X1 NOT_204( .ZN(g6510), .A(I8450) );
  INV_X1 NOT_205( .ZN(I6280), .A(g4430) );
  INV_X2 NOT_206( .ZN(g4933), .A(I6625) );
  INV_X2 NOT_207( .ZN(g5420), .A(I7086) );
  INV_X1 NOT_208( .ZN(g4521), .A(I6075) );
  INV_X1 NOT_209( .ZN(g1672), .A(g1094) );
  INV_X1 NOT_210( .ZN(I7058), .A(g5281) );
  INV_X1 NOT_211( .ZN(I2887), .A(g1123) );
  INV_X1 NOT_212( .ZN(I2122), .A(g689) );
  INV_X1 NOT_213( .ZN(g1477), .A(g952) );
  INV_X1 NOT_214( .ZN(g3232), .A(I4495) );
  INV_X1 NOT_215( .ZN(I2228), .A(g15) );
  INV_X1 NOT_216( .ZN(g5794), .A(I7593) );
  INV_X1 NOT_217( .ZN(g1643), .A(I2608) );
  INV_X1 NOT_218( .ZN(I4495), .A(g3022) );
  INV_X1 NOT_219( .ZN(I4437), .A(g2108) );
  INV_X1 NOT_220( .ZN(g2705), .A(I3858) );
  INV_X1 NOT_221( .ZN(g3813), .A(g3258) );
  INV_X1 NOT_222( .ZN(I8650), .A(g6529) );
  INV_X1 NOT_223( .ZN(I3379), .A(g1647) );
  INV_X1 NOT_224( .ZN(g2242), .A(I3373) );
  INV_X1 NOT_225( .ZN(g1205), .A(g45) );
  INV_X1 NOT_226( .ZN(I2033), .A(g678) );
  INV_X1 NOT_227( .ZN(I5871), .A(g3744) );
  INV_X1 NOT_228( .ZN(g774), .A(I1859) );
  INV_X1 NOT_229( .ZN(g6819), .A(I8994) );
  INV_X1 NOT_230( .ZN(g6694), .A(I8800) );
  INV_X1 NOT_231( .ZN(g4379), .A(I5848) );
  INV_X1 NOT_232( .ZN(g5905), .A(g5852) );
  INV_X1 NOT_233( .ZN(g3519), .A(g2740) );
  INV_X1 NOT_234( .ZN(I7856), .A(g5994) );
  INV_X2 NOT_235( .ZN(g921), .A(g111) );
  INV_X2 NOT_236( .ZN(g1551), .A(g1011) );
  INV_X1 NOT_237( .ZN(g1742), .A(I2756) );
  INV_X1 NOT_238( .ZN(I4752), .A(g2859) );
  INV_X1 NOT_239( .ZN(g6488), .A(g6367) );
  INV_X1 NOT_240( .ZN(g2254), .A(I3391) );
  INV_X1 NOT_241( .ZN(I8594), .A(g6446) );
  INV_X1 NOT_242( .ZN(g2814), .A(I4023) );
  INV_X1 NOT_243( .ZN(g4289), .A(I5746) );
  INV_X1 NOT_244( .ZN(g4658), .A(I6247) );
  INV_X1 NOT_245( .ZN(I6756), .A(g4775) );
  INV_X1 NOT_246( .ZN(g6701), .A(I8821) );
  INV_X1 NOT_247( .ZN(I8972), .A(g6795) );
  INV_X1 NOT_248( .ZN(I3271), .A(g1748) );
  INV_X1 NOT_249( .ZN(I2845), .A(g1193) );
  INV_X1 NOT_250( .ZN(g5300), .A(I6952) );
  INV_X1 NOT_251( .ZN(g2350), .A(I3502) );
  INV_X1 NOT_252( .ZN(I8806), .A(g6686) );
  INV_X1 NOT_253( .ZN(I3611), .A(g1771) );
  INV_X1 NOT_254( .ZN(I2137), .A(g1) );
  INV_X1 NOT_255( .ZN(I8943), .A(g6774) );
  INV_X1 NOT_256( .ZN(I2337), .A(g1209) );
  INV_X1 NOT_257( .ZN(I2913), .A(g1792) );
  INV_X1 NOT_258( .ZN(g1754), .A(I2773) );
  INV_X1 NOT_259( .ZN(g6886), .A(I9125) );
  INV_X1 NOT_260( .ZN(g2409), .A(g1815) );
  INV_X1 NOT_261( .ZN(g894), .A(I1917) );
  INV_X1 NOT_262( .ZN(g1273), .A(g839) );
  INV_X2 NOT_263( .ZN(I5424), .A(g3725) );
  INV_X2 NOT_264( .ZN(I6403), .A(g4492) );
  INV_X1 NOT_265( .ZN(g6314), .A(I8044) );
  INV_X1 NOT_266( .ZN(g4799), .A(g4485) );
  INV_X1 NOT_267( .ZN(I9155), .A(g6882) );
  INV_X1 NOT_268( .ZN(g2836), .A(g2509) );
  INV_X1 NOT_269( .ZN(g2212), .A(I3343) );
  INV_X1 NOT_270( .ZN(I6763), .A(g4780) );
  INV_X1 NOT_271( .ZN(g3860), .A(I5081) );
  INV_X1 NOT_272( .ZN(g2967), .A(I4166) );
  INV_X1 NOT_273( .ZN(g6825), .A(I9008) );
  INV_X1 NOT_274( .ZN(g5440), .A(g5266) );
  INV_X1 NOT_275( .ZN(g3710), .A(g3029) );
  INV_X1 NOT_276( .ZN(I5523), .A(g3840) );
  INV_X1 NOT_277( .ZN(g843), .A(g574) );
  INV_X1 NOT_278( .ZN(g1543), .A(g1006) );
  INV_X1 NOT_279( .ZN(g4132), .A(I5478) );
  INV_X1 NOT_280( .ZN(g6408), .A(g6283) );
  INV_X1 NOT_281( .ZN(g4153), .A(I5545) );
  INV_X1 NOT_282( .ZN(I6359), .A(g4566) );
  INV_X1 NOT_283( .ZN(g6136), .A(I7856) );
  INV_X1 NOT_284( .ZN(g2822), .A(I4031) );
  INV_X1 NOT_285( .ZN(I8891), .A(g6706) );
  INV_X1 NOT_286( .ZN(I8913), .A(g6743) );
  INV_X1 NOT_287( .ZN(I2692), .A(g1037) );
  INV_X1 NOT_288( .ZN(g6594), .A(I8650) );
  INV_X1 NOT_289( .ZN(g946), .A(g361) );
  INV_X1 NOT_290( .ZN(g1729), .A(I2731) );
  INV_X4 NOT_291( .ZN(I5551), .A(g4059) );
  INV_X4 NOT_292( .ZN(g4802), .A(I6470) );
  INV_X1 NOT_293( .ZN(g3962), .A(I5214) );
  INV_X1 NOT_294( .ZN(I2154), .A(g14) );
  INV_X1 NOT_295( .ZN(I4189), .A(g2159) );
  INV_X1 NOT_296( .ZN(I5499), .A(g3847) );
  INV_X1 NOT_297( .ZN(g5151), .A(I6819) );
  INV_X1 NOT_298( .ZN(g3158), .A(I4398) );
  INV_X1 NOT_299( .ZN(g6806), .A(I8978) );
  INV_X1 NOT_300( .ZN(I4706), .A(g2877) );
  INV_X1 NOT_301( .ZN(g5875), .A(I7637) );
  INV_X1 NOT_302( .ZN(g5530), .A(I7270) );
  INV_X1 NOT_303( .ZN(I9167), .A(g6878) );
  INV_X1 NOT_304( .ZN(I5926), .A(g4153) );
  INV_X1 NOT_305( .ZN(g2921), .A(g1950) );
  INV_X1 NOT_306( .ZN(g6065), .A(g5784) );
  INV_X1 NOT_307( .ZN(I6315), .A(g4446) );
  INV_X1 NOT_308( .ZN(I4371), .A(g2555) );
  INV_X1 NOT_309( .ZN(g6887), .A(I9128) );
  INV_X1 NOT_310( .ZN(I4429), .A(g2102) );
  INV_X1 NOT_311( .ZN(g6122), .A(I7838) );
  INV_X1 NOT_312( .ZN(g6465), .A(I8329) );
  INV_X1 NOT_313( .ZN(g6322), .A(I8056) );
  INV_X1 NOT_314( .ZN(g1660), .A(g985) );
  INV_X1 NOT_315( .ZN(g1946), .A(I3053) );
  INV_X4 NOT_316( .ZN(g6230), .A(g6040) );
  INV_X4 NOT_317( .ZN(g5010), .A(I6646) );
  INV_X4 NOT_318( .ZN(g4511), .A(I6045) );
  INV_X1 NOT_319( .ZN(I6874), .A(g4861) );
  INV_X1 NOT_320( .ZN(g2895), .A(g1894) );
  INV_X1 NOT_321( .ZN(g6033), .A(g5824) );
  INV_X1 NOT_322( .ZN(g2837), .A(g2512) );
  INV_X1 NOT_323( .ZN(I2979), .A(g1263) );
  INV_X1 NOT_324( .ZN(I3864), .A(g2044) );
  INV_X1 NOT_325( .ZN(g5884), .A(g5864) );
  INV_X1 NOT_326( .ZN(I8342), .A(g6314) );
  INV_X1 NOT_327( .ZN(I2218), .A(g11) );
  INV_X1 NOT_328( .ZN(g1513), .A(g878) );
  INV_X1 NOT_329( .ZN(I2312), .A(g897) );
  INV_X1 NOT_330( .ZN(I3714), .A(g1852) );
  INV_X1 NOT_331( .ZN(I4297), .A(g2555) );
  INV_X1 NOT_332( .ZN(I8255), .A(g6292) );
  INV_X1 NOT_333( .ZN(I8815), .A(g6689) );
  INV_X1 NOT_334( .ZN(g4492), .A(I5998) );
  INV_X1 NOT_335( .ZN(I1868), .A(g280) );
  INV_X1 NOT_336( .ZN(I7608), .A(g5605) );
  INV_X1 NOT_337( .ZN(I5862), .A(g3863) );
  INV_X1 NOT_338( .ZN(g1679), .A(g985) );
  INV_X1 NOT_339( .ZN(g1378), .A(I2414) );
  INV_X1 NOT_340( .ZN(g4714), .A(I6324) );
  INV_X1 NOT_341( .ZN(I2293), .A(g971) );
  INV_X1 NOT_342( .ZN(g5278), .A(I6937) );
  INV_X1 NOT_343( .ZN(g3284), .A(g3019) );
  INV_X1 NOT_344( .ZN(I4684), .A(g2687) );
  INV_X1 NOT_345( .ZN(I8497), .A(g6481) );
  INV_X1 NOT_346( .ZN(g3239), .A(I4516) );
  INV_X1 NOT_347( .ZN(I6537), .A(g4711) );
  INV_X1 NOT_348( .ZN(g3545), .A(g3085) );
  INV_X1 NOT_349( .ZN(g2788), .A(I3983) );
  INV_X8 NOT_350( .ZN(g6137), .A(I7859) );
  INV_X1 NOT_351( .ZN(g5667), .A(g5524) );
  INV_X1 NOT_352( .ZN(g6891), .A(I9140) );
  INV_X1 NOT_353( .ZN(g1831), .A(I2907) );
  INV_X1 NOT_354( .ZN(g1335), .A(I2358) );
  INV_X1 NOT_355( .ZN(g3380), .A(g2831) );
  INV_X1 NOT_356( .ZN(I4791), .A(g2814) );
  INV_X1 NOT_357( .ZN(g6337), .A(I8089) );
  INV_X1 NOT_358( .ZN(I4309), .A(g2525) );
  INV_X1 NOT_359( .ZN(I2828), .A(g1193) );
  INV_X1 NOT_360( .ZN(g3832), .A(I5023) );
  INV_X1 NOT_361( .ZN(g1288), .A(I2269) );
  INV_X1 NOT_362( .ZN(g5566), .A(I7318) );
  INV_X1 NOT_363( .ZN(g3853), .A(I5068) );
  INV_X1 NOT_364( .ZN(I3736), .A(g2460) );
  INV_X1 NOT_365( .ZN(I6612), .A(g4660) );
  INV_X1 NOT_366( .ZN(I7161), .A(g5465) );
  INV_X1 NOT_367( .ZN(I7361), .A(g5566) );
  INV_X1 NOT_368( .ZN(g2842), .A(I4050) );
  INV_X1 NOT_369( .ZN(g1805), .A(I2854) );
  INV_X1 NOT_370( .ZN(I6417), .A(g4617) );
  INV_X1 NOT_371( .ZN(I3623), .A(g1491) );
  INV_X8 NOT_372( .ZN(g4262), .A(I5713) );
  INV_X8 NOT_373( .ZN(I7051), .A(g5219) );
  INV_X8 NOT_374( .ZN(I2221), .A(g43) );
  INV_X1 NOT_375( .ZN(g3559), .A(g2603) );
  INV_X1 NOT_376( .ZN(g4736), .A(I6366) );
  INV_X1 NOT_377( .ZN(g2485), .A(I3614) );
  INV_X1 NOT_378( .ZN(I7451), .A(g5597) );
  INV_X1 NOT_379( .ZN(I2703), .A(g1189) );
  INV_X1 NOT_380( .ZN(I8267), .A(g6297) );
  INV_X1 NOT_381( .ZN(g4623), .A(g4262) );
  INV_X1 NOT_382( .ZN(g1947), .A(I3056) );
  INV_X1 NOT_383( .ZN(I5885), .A(g3746) );
  INV_X1 NOT_384( .ZN(I7999), .A(g6137) );
  INV_X1 NOT_385( .ZN(g878), .A(g639) );
  INV_X1 NOT_386( .ZN(I7146), .A(g5231) );
  INV_X1 NOT_387( .ZN(I6330), .A(g4560) );
  INV_X1 NOT_388( .ZN(I7346), .A(g5531) );
  INV_X1 NOT_389( .ZN(I3871), .A(g2145) );
  INV_X1 NOT_390( .ZN(I8329), .A(g6305) );
  INV_X1 NOT_391( .ZN(g4375), .A(I5840) );
  INV_X1 NOT_392( .ZN(g4871), .A(I6599) );
  INV_X1 NOT_393( .ZN(I8761), .A(g6563) );
  INV_X1 NOT_394( .ZN(g3204), .A(I4441) );
  INV_X1 NOT_395( .ZN(g4722), .A(I6346) );
  INV_X1 NOT_396( .ZN(g710), .A(g128) );
  INV_X1 NOT_397( .ZN(I4498), .A(g2686) );
  INV_X1 NOT_398( .ZN(g829), .A(g323) );
  INV_X1 NOT_399( .ZN(g5113), .A(I6753) );
  INV_X1 NOT_400( .ZN(g1632), .A(g760) );
  INV_X1 NOT_401( .ZN(g1037), .A(I2067) );
  INV_X1 NOT_402( .ZN(g3100), .A(I4347) );
  INV_X1 NOT_403( .ZN(I8828), .A(g6661) );
  INV_X1 NOT_404( .ZN(g6726), .A(I8872) );
  INV_X8 NOT_405( .ZN(g6497), .A(I8411) );
  INV_X1 NOT_406( .ZN(g1653), .A(I2630) );
  INV_X1 NOT_407( .ZN(g2640), .A(I3782) );
  INV_X1 NOT_408( .ZN(I8727), .A(g6536) );
  INV_X1 NOT_409( .ZN(g2031), .A(I3140) );
  INV_X1 NOT_410( .ZN(I5436), .A(g3729) );
  INV_X1 NOT_411( .ZN(g2252), .A(I3385) );
  INV_X1 NOT_412( .ZN(g5908), .A(g5753) );
  INV_X1 NOT_413( .ZN(g2958), .A(g1861) );
  INV_X1 NOT_414( .ZN(I7472), .A(g5626) );
  INV_X1 NOT_415( .ZN(g2176), .A(I3319) );
  INV_X1 NOT_416( .ZN(I2716), .A(g1115) );
  INV_X1 NOT_417( .ZN(I5831), .A(g3842) );
  INV_X1 NOT_418( .ZN(I2349), .A(g1160) );
  INV_X1 NOT_419( .ZN(g4139), .A(I5499) );
  INV_X1 NOT_420( .ZN(I5182), .A(g3271) );
  INV_X1 NOT_421( .ZN(g5518), .A(I7258) );
  INV_X1 NOT_422( .ZN(g5567), .A(g5418) );
  INV_X1 NOT_423( .ZN(I5382), .A(g3952) );
  INV_X1 NOT_424( .ZN(g2405), .A(I3543) );
  INV_X1 NOT_425( .ZN(I2848), .A(g1193) );
  INV_X1 NOT_426( .ZN(g1917), .A(I3016) );
  INV_X1 NOT_427( .ZN(g2829), .A(g2491) );
  INV_X1 NOT_428( .ZN(g2765), .A(I3946) );
  INV_X1 NOT_429( .ZN(I7116), .A(g5299) );
  INV_X8 NOT_430( .ZN(I4019), .A(g1841) );
  INV_X8 NOT_431( .ZN(g4424), .A(I5923) );
  INV_X8 NOT_432( .ZN(I6090), .A(g4393) );
  INV_X1 NOT_433( .ZN(I4362), .A(g2555) );
  INV_X1 NOT_434( .ZN(I3672), .A(g1656) );
  INV_X1 NOT_435( .ZN(g3040), .A(I4255) );
  INV_X1 NOT_436( .ZN(I3077), .A(g1439) );
  INV_X1 NOT_437( .ZN(g4809), .A(I6485) );
  INV_X1 NOT_438( .ZN(g5593), .A(I7355) );
  INV_X1 NOT_439( .ZN(g3440), .A(I4678) );
  INV_X1 NOT_440( .ZN(g3969), .A(I5233) );
  INV_X1 NOT_441( .ZN(g6312), .A(I8040) );
  INV_X1 NOT_442( .ZN(I6366), .A(g4569) );
  INV_X1 NOT_443( .ZN(I4452), .A(g2117) );
  INV_X1 NOT_444( .ZN(g2974), .A(I4173) );
  INV_X1 NOT_445( .ZN(g6401), .A(I8217) );
  INV_X1 NOT_446( .ZN(g895), .A(g139) );
  INV_X1 NOT_447( .ZN(I6456), .A(g4633) );
  INV_X1 NOT_448( .ZN(g4523), .A(I6081) );
  INV_X1 NOT_449( .ZN(g1233), .A(I2231) );
  INV_X1 NOT_450( .ZN(I6649), .A(g4693) );
  INV_X1 NOT_451( .ZN(g4643), .A(g4293) );
  INV_X1 NOT_452( .ZN(g5264), .A(g4943) );
  INV_X1 NOT_453( .ZN(I9158), .A(g6887) );
  INV_X1 NOT_454( .ZN(g1054), .A(g485) );
  INV_X1 NOT_455( .ZN(g5160), .A(g5099) );
  INV_X1 NOT_456( .ZN(g2796), .A(I3999) );
  INV_X1 NOT_457( .ZN(I6355), .A(g4569) );
  INV_X1 NOT_458( .ZN(g2473), .A(I3605) );
  INV_X1 NOT_459( .ZN(I3099), .A(g1519) );
  INV_X1 NOT_460( .ZN(I8576), .A(g6436) );
  INV_X1 NOT_461( .ZN(g1770), .A(I2805) );
  INV_X1 NOT_462( .ZN(I8866), .A(g6701) );
  INV_X1 NOT_463( .ZN(I3304), .A(g1740) );
  INV_X1 NOT_464( .ZN(I4486), .A(g3093) );
  INV_X1 NOT_465( .ZN(g5521), .A(I7261) );
  INV_X1 NOT_466( .ZN(I3499), .A(g1450) );
  INV_X1 NOT_467( .ZN(I8716), .A(g6518) );
  INV_X1 NOT_468( .ZN(g1725), .A(g1113) );
  INV_X1 NOT_469( .ZN(I7596), .A(g5605) );
  INV_X1 NOT_470( .ZN(g6727), .A(I8875) );
  INV_X1 NOT_471( .ZN(g3875), .A(I5106) );
  INV_X1 NOT_472( .ZN(g2324), .A(I3478) );
  INV_X1 NOT_473( .ZN(I4504), .A(g2726) );
  INV_X1 NOT_474( .ZN(I2119), .A(g688) );
  INV_X1 NOT_475( .ZN(g5450), .A(g5292) );
  INV_X1 NOT_476( .ZN(I5037), .A(g3705) );
  INV_X1 NOT_477( .ZN(g5996), .A(g5824) );
  INV_X1 NOT_478( .ZN(g4104), .A(I5394) );
  INV_X1 NOT_479( .ZN(g6592), .A(I8644) );
  INV_X1 NOT_480( .ZN(g4099), .A(I5379) );
  INV_X1 NOT_481( .ZN(g4499), .A(I6015) );
  INV_X1 NOT_482( .ZN(I2352), .A(g1161) );
  INV_X1 NOT_483( .ZN(I6063), .A(g4381) );
  INV_X1 NOT_484( .ZN(g6746), .A(I8916) );
  INV_X1 NOT_485( .ZN(I2867), .A(g1143) );
  INV_X1 NOT_486( .ZN(I8699), .A(g6573) );
  INV_X1 NOT_487( .ZN(g2177), .A(I3322) );
  INV_X1 NOT_488( .ZN(g5179), .A(g5099) );
  INV_X1 NOT_489( .ZN(g5379), .A(I7035) );
  INV_X1 NOT_490( .ZN(I2893), .A(g1236) );
  INV_X1 NOT_491( .ZN(g5878), .A(I7646) );
  INV_X1 NOT_492( .ZN(I3044), .A(g1257) );
  INV_X1 NOT_493( .ZN(g1189), .A(I2196) );
  INV_X1 NOT_494( .ZN(g3839), .A(I5040) );
  INV_X1 NOT_495( .ZN(g6932), .A(I9217) );
  INV_X1 NOT_496( .ZN(g4273), .A(I5728) );
  INV_X1 NOT_497( .ZN(g5658), .A(g5512) );
  INV_X1 NOT_498( .ZN(g6624), .A(I8730) );
  INV_X1 NOT_499( .ZN(I6118), .A(g4406) );
  INV_X1 NOT_500( .ZN(I6318), .A(g4447) );
  INV_X32 NOT_501( .ZN(I3983), .A(g2276) );
  INV_X32 NOT_502( .ZN(g2849), .A(g2577) );
  INV_X1 NOT_503( .ZN(I3572), .A(g1295) );
  INV_X1 NOT_504( .ZN(g1787), .A(I2835) );
  INV_X1 NOT_505( .ZN(I5442), .A(g3731) );
  INV_X1 NOT_506( .ZN(I4678), .A(g2670) );
  INV_X1 NOT_507( .ZN(I6057), .A(g4379) );
  INV_X1 NOT_508( .ZN(I8524), .A(g6496) );
  INV_X1 NOT_509( .ZN(I4331), .A(g2555) );
  INV_X1 NOT_510( .ZN(I8644), .A(g6526) );
  INV_X1 NOT_511( .ZN(I3543), .A(g1461) );
  INV_X1 NOT_512( .ZN(I6989), .A(g5307) );
  INV_X1 NOT_513( .ZN(I2614), .A(g1123) );
  INV_X1 NOT_514( .ZN(g1675), .A(g1101) );
  INV_X1 NOT_515( .ZN(I2370), .A(g1123) );
  INV_X1 NOT_516( .ZN(I2125), .A(g698) );
  INV_X1 NOT_517( .ZN(g3235), .A(I4504) );
  INV_X1 NOT_518( .ZN(g3343), .A(g3090) );
  INV_X1 NOT_519( .ZN(I5233), .A(g3571) );
  INV_X1 NOT_520( .ZN(I2821), .A(g1221) );
  INV_X1 NOT_521( .ZN(g4712), .A(I6318) );
  INV_X1 NOT_522( .ZN(g985), .A(g638) );
  INV_X1 NOT_523( .ZN(g6576), .A(g6487) );
  INV_X1 NOT_524( .ZN(I6549), .A(g4699) );
  INV_X16 NOT_525( .ZN(I8258), .A(g6293) );
  INV_X1 NOT_526( .ZN(I8818), .A(g6690) );
  INV_X1 NOT_527( .ZN(I3534), .A(g1295) );
  INV_X1 NOT_528( .ZN(g2245), .A(I3382) );
  INV_X1 NOT_529( .ZN(I3729), .A(g2436) );
  INV_X1 NOT_530( .ZN(I3961), .A(g1835) );
  INV_X1 NOT_531( .ZN(I5454), .A(g3874) );
  INV_X1 NOT_532( .ZN(g2291), .A(I3434) );
  INV_X1 NOT_533( .ZN(g5997), .A(g5854) );
  INV_X1 NOT_534( .ZN(g4534), .A(I6114) );
  INV_X1 NOT_535( .ZN(I3927), .A(g2245) );
  INV_X1 NOT_536( .ZN(I5532), .A(g3861) );
  INV_X1 NOT_537( .ZN(g1684), .A(I2668) );
  INV_X1 NOT_538( .ZN(g6699), .A(I8815) );
  INV_X1 NOT_539( .ZN(g1639), .A(g815) );
  INV_X1 NOT_540( .ZN(g1338), .A(I2367) );
  INV_X1 NOT_541( .ZN(g1963), .A(I3074) );
  INV_X1 NOT_542( .ZN(I8186), .A(g6179) );
  INV_X1 NOT_543( .ZN(I6321), .A(g4559) );
  INV_X1 NOT_544( .ZN(I4226), .A(g2525) );
  INV_X1 NOT_545( .ZN(g1109), .A(I2137) );
  INV_X1 NOT_546( .ZN(g1791), .A(I2845) );
  INV_X1 NOT_547( .ZN(I8975), .A(g6791) );
  INV_X1 NOT_548( .ZN(I3946), .A(g2256) );
  INV_X1 NOT_549( .ZN(g889), .A(g310) );
  INV_X1 NOT_550( .ZN(I2306), .A(g896) );
  INV_X1 NOT_551( .ZN(g3792), .A(g3388) );
  INV_X1 NOT_552( .ZN(I6625), .A(g4745) );
  INV_X1 NOT_553( .ZN(g2819), .A(g2467) );
  INV_X1 NOT_554( .ZN(g4014), .A(I5316) );
  INV_X1 NOT_555( .ZN(I8426), .A(g6424) );
  INV_X1 NOT_556( .ZN(I5412), .A(g4034) );
  INV_X32 NOT_557( .ZN(g4660), .A(I6253) );
  INV_X32 NOT_558( .ZN(I6253), .A(g4608) );
  INV_X1 NOT_559( .ZN(g2088), .A(I3202) );
  INV_X1 NOT_560( .ZN(g2923), .A(g1969) );
  INV_X1 NOT_561( .ZN(I4173), .A(g2408) );
  INV_X1 NOT_562( .ZN(I8614), .A(g6537) );
  INV_X1 NOT_563( .ZN(I3513), .A(g1450) );
  INV_X1 NOT_564( .ZN(g2488), .A(I3617) );
  INV_X1 NOT_565( .ZN(g1759), .A(I2782) );
  INV_X1 NOT_566( .ZN(I2756), .A(g1175) );
  INV_X1 NOT_567( .ZN(g2701), .A(I3855) );
  INV_X1 NOT_568( .ZN(I7190), .A(g5432) );
  INV_X1 NOT_569( .ZN(I8821), .A(g6691) );
  INV_X1 NOT_570( .ZN(g6524), .A(I8488) );
  INV_X1 NOT_571( .ZN(I6740), .A(g4781) );
  INV_X1 NOT_572( .ZN(g4513), .A(I6051) );
  INV_X1 NOT_573( .ZN(I8984), .A(g6794) );
  INV_X1 NOT_574( .ZN(I7501), .A(g5596) );
  INV_X1 NOT_575( .ZN(g1957), .A(I3068) );
  INV_X1 NOT_576( .ZN(g2215), .A(I3352) );
  INV_X1 NOT_577( .ZN(g6119), .A(I7829) );
  INV_X1 NOT_578( .ZN(I2904), .A(g1256) );
  INV_X1 NOT_579( .ZN(g6319), .A(I8051) );
  INV_X1 NOT_580( .ZN(g1049), .A(g266) );
  INV_X1 NOT_581( .ZN(g5901), .A(g5753) );
  INV_X1 NOT_582( .ZN(g2886), .A(g1966) );
  INV_X2 NOT_583( .ZN(I6552), .A(g4702) );
  INV_X1 NOT_584( .ZN(I4059), .A(g1878) );
  INV_X1 NOT_585( .ZN(g4036), .A(I5337) );
  INV_X1 NOT_586( .ZN(g3094), .A(I4337) );
  INV_X1 NOT_587( .ZN(I4459), .A(g2134) );
  INV_X1 NOT_588( .ZN(I8544), .A(g6453) );
  INV_X1 NOT_589( .ZN(g4679), .A(I6269) );
  INV_X1 NOT_590( .ZN(g6352), .A(I8110) );
  INV_X1 NOT_591( .ZN(g6818), .A(I8991) );
  INV_X1 NOT_592( .ZN(g6577), .A(g6488) );
  INV_X1 NOT_593( .ZN(I1847), .A(g209) );
  INV_X1 NOT_594( .ZN(I3288), .A(g1710) );
  INV_X1 NOT_595( .ZN(g3567), .A(g3074) );
  INV_X1 NOT_596( .ZN(I3382), .A(g1284) );
  INV_X1 NOT_597( .ZN(g1715), .A(I2716) );
  INV_X1 NOT_598( .ZN(g4135), .A(I5487) );
  INV_X1 NOT_599( .ZN(I7704), .A(g5723) );
  INV_X1 NOT_600( .ZN(g848), .A(g594) );
  INV_X1 NOT_601( .ZN(g5092), .A(g4753) );
  INV_X1 NOT_602( .ZN(g1498), .A(I2479) );
  INV_X1 NOT_603( .ZN(I2763), .A(g1236) );
  INV_X1 NOT_604( .ZN(g2870), .A(g2296) );
  INV_X1 NOT_605( .ZN(I3022), .A(g1426) );
  INV_X1 NOT_606( .ZN(I4261), .A(g1857) );
  INV_X1 NOT_607( .ZN(I2391), .A(g774) );
  INV_X1 NOT_608( .ZN(g4382), .A(I5857) );
  INV_X1 NOT_609( .ZN(g3776), .A(g3466) );
  INV_X1 NOT_610( .ZN(g6893), .A(I9146) );
  INV_X1 NOT_611( .ZN(g1833), .A(I2913) );
  INV_X4 NOT_612( .ZN(I3422), .A(g1641) );
  INV_X4 NOT_613( .ZN(g5574), .A(g5407) );
  INV_X1 NOT_614( .ZN(I3749), .A(g2484) );
  INV_X1 NOT_615( .ZN(g3593), .A(g2997) );
  INV_X1 NOT_616( .ZN(g6211), .A(g5992) );
  INV_X1 NOT_617( .ZN(g2650), .A(I3794) );
  INV_X1 NOT_618( .ZN(g5714), .A(I7475) );
  INV_X1 NOT_619( .ZN(g932), .A(g337) );
  INV_X1 NOT_620( .ZN(I8061), .A(g6113) );
  INV_X1 NOT_621( .ZN(g4805), .A(g4473) );
  INV_X1 NOT_622( .ZN(g4022), .A(I5328) );
  INV_X1 NOT_623( .ZN(g1584), .A(g743) );
  INV_X1 NOT_624( .ZN(g4422), .A(g4111) );
  INV_X1 NOT_625( .ZN(g6599), .A(I8665) );
  INV_X1 NOT_626( .ZN(g1539), .A(g878) );
  INV_X1 NOT_627( .ZN(I5109), .A(g3710) );
  INV_X1 NOT_628( .ZN(g2408), .A(I3546) );
  INV_X1 NOT_629( .ZN(I2159), .A(g465) );
  INV_X1 NOT_630( .ZN(I6570), .A(g4719) );
  INV_X1 NOT_631( .ZN(g2136), .A(g1395) );
  INV_X1 NOT_632( .ZN(I4664), .A(g2924) );
  INV_X1 NOT_633( .ZN(I8027), .A(g6237) );
  INV_X1 NOT_634( .ZN(I4246), .A(g2194) );
  INV_X1 NOT_635( .ZN(g2336), .A(I3488) );
  INV_X1 NOT_636( .ZN(g5580), .A(I7336) );
  INV_X1 NOT_637( .ZN(g716), .A(I1832) );
  INV_X1 NOT_638( .ZN(I3560), .A(g1673) );
  INV_X1 NOT_639( .ZN(g736), .A(I1841) );
  INV_X4 NOT_640( .ZN(I6525), .A(g4770) );
  INV_X1 NOT_641( .ZN(g2768), .A(g2367) );
  INV_X1 NOT_642( .ZN(g6370), .A(I8174) );
  INV_X1 NOT_643( .ZN(g2594), .A(I3723) );
  INV_X1 NOT_644( .ZN(g4798), .A(I6464) );
  INV_X1 NOT_645( .ZN(g6325), .A(I8061) );
  INV_X1 NOT_646( .ZN(g6821), .A(g6785) );
  INV_X1 NOT_647( .ZN(g4560), .A(g4188) );
  INV_X1 NOT_648( .ZN(g2806), .A(g2446) );
  INV_X1 NOT_649( .ZN(I3632), .A(g1295) );
  INV_X1 NOT_650( .ZN(g3450), .A(I4688) );
  INV_X1 NOT_651( .ZN(I3037), .A(g1769) );
  INV_X1 NOT_652( .ZN(g6939), .A(I9230) );
  INV_X1 NOT_653( .ZN(g1052), .A(g668) );
  INV_X1 NOT_654( .ZN(I3653), .A(g1305) );
  INV_X1 NOT_655( .ZN(I3102), .A(g1426) );
  INV_X1 NOT_656( .ZN(I2115), .A(g687) );
  INV_X1 NOT_657( .ZN(I2315), .A(g1222) );
  INV_X1 NOT_658( .ZN(I2811), .A(g1209) );
  INV_X1 NOT_659( .ZN(g6083), .A(g5809) );
  INV_X1 NOT_660( .ZN(g2887), .A(g1858) );
  INV_X1 NOT_661( .ZN(I2047), .A(g682) );
  INV_X1 NOT_662( .ZN(g6544), .A(I8544) );
  INV_X1 NOT_663( .ZN(I6607), .A(g4745) );
  INV_X1 NOT_664( .ZN(g4632), .A(g4281) );
  INV_X1 NOT_665( .ZN(g5889), .A(g5742) );
  INV_X1 NOT_666( .ZN(g5476), .A(I7164) );
  INV_X1 NOT_667( .ZN(g2934), .A(g2004) );
  INV_X4 NOT_668( .ZN(g2230), .A(I3355) );
  INV_X4 NOT_669( .ZN(g4437), .A(I5948) );
  INV_X1 NOT_670( .ZN(g4102), .A(I5388) );
  INV_X1 NOT_671( .ZN(g4302), .A(g4068) );
  INV_X1 NOT_672( .ZN(I5865), .A(g3743) );
  INV_X1 NOT_673( .ZN(g6106), .A(I7814) );
  INV_X1 NOT_674( .ZN(g4579), .A(g4206) );
  INV_X1 NOT_675( .ZN(g4869), .A(g4662) );
  INV_X1 NOT_676( .ZN(g6306), .A(I8030) );
  INV_X1 NOT_677( .ZN(I3752), .A(g2044) );
  INV_X1 NOT_678( .ZN(g5375), .A(I7029) );
  INV_X1 NOT_679( .ZN(I8107), .A(g6136) );
  INV_X1 NOT_680( .ZN(g4719), .A(I6337) );
  INV_X1 NOT_681( .ZN(g1730), .A(g1114) );
  INV_X1 NOT_682( .ZN(g3289), .A(g3034) );
  INV_X1 NOT_683( .ZN(g1504), .A(I2485) );
  INV_X1 NOT_684( .ZN(g3777), .A(g3388) );
  INV_X1 NOT_685( .ZN(I6587), .A(g4803) );
  INV_X1 NOT_686( .ZN(I8159), .A(g6167) );
  INV_X1 NOT_687( .ZN(I6111), .A(g4404) );
  INV_X1 NOT_688( .ZN(g3835), .A(I5030) );
  INV_X1 NOT_689( .ZN(I6311), .A(g4444) );
  INV_X1 NOT_690( .ZN(I8223), .A(g6325) );
  INV_X1 NOT_691( .ZN(g2096), .A(I3212) );
  INV_X1 NOT_692( .ZN(I9143), .A(g6886) );
  INV_X1 NOT_693( .ZN(g3882), .A(I5119) );
  INV_X1 NOT_694( .ZN(g1070), .A(g94) );
  INV_X1 NOT_695( .ZN(g2550), .A(I3665) );
  INV_X2 NOT_696( .ZN(I6615), .A(g4745) );
  INV_X2 NOT_697( .ZN(g3271), .A(g3042) );
  INV_X1 NOT_698( .ZN(I4671), .A(g2928) );
  INV_X1 NOT_699( .ZN(I2880), .A(g1143) );
  INV_X1 NOT_700( .ZN(g2845), .A(g2565) );
  INV_X1 NOT_701( .ZN(g1897), .A(I2992) );
  INV_X1 NOT_702( .ZN(g6622), .A(I8724) );
  INV_X1 NOT_703( .ZN(I2537), .A(g971) );
  INV_X1 NOT_704( .ZN(I5896), .A(g3879) );
  INV_X1 NOT_705( .ZN(g2195), .A(I3334) );
  INV_X1 NOT_706( .ZN(g4265), .A(I5716) );
  INV_X1 NOT_707( .ZN(g2891), .A(g1884) );
  INV_X1 NOT_708( .ZN(g2913), .A(g1925) );
  INV_X1 NOT_709( .ZN(g5139), .A(I6795) );
  INV_X1 NOT_710( .ZN(I3364), .A(g1648) );
  INV_X1 NOT_711( .ZN(g5384), .A(g5220) );
  INV_X1 NOT_712( .ZN(I9134), .A(g6864) );
  INV_X1 NOT_713( .ZN(I2272), .A(g908) );
  INV_X1 NOT_714( .ZN(g6904), .A(I9179) );
  INV_X1 NOT_715( .ZN(g4786), .A(I6448) );
  INV_X1 NOT_716( .ZN(g3799), .A(g3388) );
  INV_X4 NOT_717( .ZN(g6514), .A(I8462) );
  INV_X4 NOT_718( .ZN(g4364), .A(I5825) );
  INV_X1 NOT_719( .ZN(I8447), .A(g6410) );
  INV_X1 NOT_720( .ZN(I3770), .A(g2145) );
  INV_X1 NOT_721( .ZN(I5019), .A(g3318) );
  INV_X1 NOT_722( .ZN(I2417), .A(g774) );
  INV_X1 NOT_723( .ZN(g6403), .A(I8223) );
  INV_X1 NOT_724( .ZN(g5809), .A(I7608) );
  INV_X1 NOT_725( .ZN(I7683), .A(g5702) );
  INV_X1 NOT_726( .ZN(g6841), .A(I9044) );
  INV_X1 NOT_727( .ZN(g3541), .A(g2643) );
  INV_X1 NOT_728( .ZN(I2982), .A(g1426) );
  INV_X1 NOT_729( .ZN(g1678), .A(I2658) );
  INV_X1 NOT_730( .ZN(g4770), .A(I6414) );
  INV_X1 NOT_731( .ZN(g1006), .A(I2047) );
  INV_X1 NOT_732( .ZN(I2234), .A(g697) );
  INV_X1 NOT_733( .ZN(g1331), .A(I2346) );
  INV_X1 NOT_734( .ZN(g4296), .A(I5753) );
  INV_X1 NOT_735( .ZN(I2128), .A(g18) );
  INV_X1 NOT_736( .ZN(g3238), .A(I4513) );
  INV_X1 NOT_737( .ZN(I3553), .A(g1305) );
  INV_X1 NOT_738( .ZN(I6020), .A(g4176) );
  INV_X1 NOT_739( .ZN(g3332), .A(g3079) );
  INV_X1 NOT_740( .ZN(g5477), .A(I7167) );
  INV_X1 NOT_741( .ZN(I6420), .A(g4618) );
  INV_X1 NOT_742( .ZN(g6695), .A(I8803) );
  INV_X1 NOT_743( .ZN(I2330), .A(g1122) );
  INV_X1 NOT_744( .ZN(g3209), .A(I4452) );
  INV_X1 NOT_745( .ZN(I6507), .A(g4644) );
  INV_X1 NOT_746( .ZN(g4532), .A(I6108) );
  INV_X1 NOT_747( .ZN(g1682), .A(g829) );
  INV_X1 NOT_748( .ZN(g6107), .A(I7817) );
  INV_X1 NOT_749( .ZN(I9113), .A(g6855) );
  INV_X1 NOT_750( .ZN(I1856), .A(g204) );
  INV_X1 NOT_751( .ZN(g1305), .A(I2293) );
  INV_X1 NOT_752( .ZN(g6536), .A(I8524) );
  INV_X1 NOT_753( .ZN(g3802), .A(g3388) );
  INV_X4 NOT_754( .ZN(I5728), .A(g4022) );
  INV_X2 NOT_755( .ZN(g2481), .A(I3608) );
  INV_X1 NOT_756( .ZN(I7475), .A(g5627) );
  INV_X1 NOT_757( .ZN(g931), .A(g54) );
  INV_X1 NOT_758( .ZN(g1748), .A(I2763) );
  INV_X1 NOT_759( .ZN(g2692), .A(I3840) );
  INV_X1 NOT_760( .ZN(I4217), .A(g2163) );
  INV_X1 NOT_761( .ZN(g2097), .A(I3215) );
  INV_X1 NOT_762( .ZN(I4066), .A(g2582) );
  INV_X1 NOT_763( .ZN(g5551), .A(I7295) );
  INV_X1 NOT_764( .ZN(g5742), .A(g5686) );
  INV_X1 NOT_765( .ZN(g2726), .A(I3886) );
  INV_X1 NOT_766( .ZN(g5099), .A(I6737) );
  INV_X1 NOT_767( .ZN(g2497), .A(I3626) );
  INV_X1 NOT_768( .ZN(I5385), .A(g3962) );
  INV_X1 NOT_769( .ZN(g5304), .A(I6956) );
  INV_X1 NOT_770( .ZN(g2154), .A(I3271) );
  INV_X1 NOT_771( .ZN(g1755), .A(I2776) );
  INV_X1 NOT_772( .ZN(g4189), .A(I5597) );
  INV_X1 NOT_773( .ZN(I8978), .A(g6792) );
  INV_X1 NOT_774( .ZN(g4706), .A(I6308) );
  INV_X1 NOT_775( .ZN(g6416), .A(I8258) );
  INV_X1 NOT_776( .ZN(I8243), .A(g6286) );
  INV_X1 NOT_777( .ZN(I8417), .A(g6420) );
  INV_X1 NOT_778( .ZN(g3901), .A(g3575) );
  INV_X1 NOT_779( .ZN(I6630), .A(g4745) );
  INV_X1 NOT_780( .ZN(I7646), .A(g5774) );
  INV_X1 NOT_781( .ZN(I3675), .A(g1491) );
  INV_X1 NOT_782( .ZN(g6522), .A(I8482) );
  INV_X1 NOT_783( .ZN(g6115), .A(g5879) );
  INV_X1 NOT_784( .ZN(g1045), .A(g699) );
  INV_X1 NOT_785( .ZN(I3281), .A(g1761) );
  INV_X1 NOT_786( .ZN(I7039), .A(g5309) );
  INV_X1 NOT_787( .ZN(I7484), .A(g5630) );
  INV_X1 NOT_788( .ZN(g1173), .A(I2185) );
  INV_X2 NOT_789( .ZN(I4455), .A(g2118) );
  INV_X2 NOT_790( .ZN(I8629), .A(g6544) );
  INV_X2 NOT_791( .ZN(g5273), .A(I6930) );
  INV_X1 NOT_792( .ZN(I4133), .A(g2040) );
  INV_X1 NOT_793( .ZN(g1491), .A(I2476) );
  INV_X1 NOT_794( .ZN(g760), .A(I1853) );
  INV_X1 NOT_795( .ZN(g2783), .A(I3979) );
  INV_X1 NOT_796( .ZN(g4281), .A(I5736) );
  INV_X1 NOT_797( .ZN(g3600), .A(I4791) );
  INV_X1 NOT_798( .ZN(g2112), .A(I3240) );
  INV_X1 NOT_799( .ZN(g1283), .A(g853) );
  INV_X1 NOT_800( .ZN(g2312), .A(I3462) );
  INV_X1 NOT_801( .ZN(g1369), .A(I2405) );
  INV_X1 NOT_802( .ZN(I6750), .A(g4771) );
  INV_X1 NOT_803( .ZN(g6654), .A(I8758) );
  INV_X1 NOT_804( .ZN(g3714), .A(g3041) );
  INV_X1 NOT_805( .ZN(I7583), .A(g5605) );
  INV_X1 NOT_806( .ZN(I3684), .A(g1733) );
  INV_X1 NOT_807( .ZN(I5006), .A(g3604) );
  INV_X1 NOT_808( .ZN(I8800), .A(g6684) );
  INV_X1 NOT_809( .ZN(g1059), .A(g702) );
  INV_X4 NOT_810( .ZN(g1578), .A(I2552) );
  INV_X4 NOT_811( .ZN(g2001), .A(I3112) );
  INV_X1 NOT_812( .ZN(I5406), .A(g3976) );
  INV_X1 NOT_813( .ZN(g5572), .A(g5399) );
  INV_X1 NOT_814( .ZN(I3109), .A(g1504) );
  INV_X1 NOT_815( .ZN(I3791), .A(g2044) );
  INV_X1 NOT_816( .ZN(g2293), .A(g1567) );
  INV_X1 NOT_817( .ZN(g6880), .A(I9107) );
  INV_X1 NOT_818( .ZN(g6595), .A(I8653) );
  INV_X1 NOT_819( .ZN(g4138), .A(I5496) );
  INV_X1 NOT_820( .ZN(g1535), .A(g1088) );
  INV_X1 NOT_821( .ZN(g4639), .A(g4289) );
  INV_X1 NOT_822( .ZN(g6537), .A(I8527) );
  INV_X1 NOT_823( .ZN(g5543), .A(g5331) );
  INV_X1 NOT_824( .ZN(I3808), .A(g2125) );
  INV_X1 NOT_825( .ZN(I7276), .A(g5375) );
  INV_X1 NOT_826( .ZN(I5487), .A(g3881) );
  INV_X1 NOT_827( .ZN(I2355), .A(g1177) );
  INV_X1 NOT_828( .ZN(g4109), .A(I5409) );
  INV_X1 NOT_829( .ZN(g4309), .A(g4074) );
  INV_X1 NOT_830( .ZN(g2828), .A(g2488) );
  INV_X1 NOT_831( .ZN(g2830), .A(g2494) );
  INV_X1 NOT_832( .ZN(g2727), .A(g2324) );
  INV_X1 NOT_833( .ZN(g4808), .A(g4473) );
  INV_X1 NOT_834( .ZN(I2964), .A(g1257) );
  INV_X1 NOT_835( .ZN(g821), .A(I1880) );
  INV_X1 NOT_836( .ZN(g6612), .A(I8702) );
  INV_X1 NOT_837( .ZN(g5534), .A(I7276) );
  INV_X1 NOT_838( .ZN(g5729), .A(I7494) );
  INV_X1 NOT_839( .ZN(I6666), .A(g4740) );
  INV_X1 NOT_840( .ZN(I9179), .A(g6875) );
  INV_X1 NOT_841( .ZN(g1415), .A(g1246) );
  INV_X4 NOT_842( .ZN(g4707), .A(I6311) );
  INV_X4 NOT_843( .ZN(g6417), .A(I8261) );
  INV_X1 NOT_844( .ZN(I7404), .A(g5541) );
  INV_X1 NOT_845( .ZN(g3076), .A(I4309) );
  INV_X1 NOT_846( .ZN(I8512), .A(g6441) );
  INV_X1 NOT_847( .ZN(g3889), .A(g3575) );
  INV_X1 NOT_848( .ZN(I6528), .A(g4815) );
  INV_X1 NOT_849( .ZN(g1664), .A(I2643) );
  INV_X1 NOT_850( .ZN(g1246), .A(I2237) );
  INV_X1 NOT_851( .ZN(g6234), .A(g6057) );
  INV_X1 NOT_852( .ZN(I3575), .A(g1305) );
  INV_X1 NOT_853( .ZN(g5885), .A(g5865) );
  INV_X1 NOT_854( .ZN(g6328), .A(I8066) );
  INV_X1 NOT_855( .ZN(g1203), .A(I2207) );
  INV_X1 NOT_856( .ZN(I5445), .A(g4040) );
  INV_X1 NOT_857( .ZN(g5946), .A(g5729) );
  INV_X1 NOT_858( .ZN(g6542), .A(I8538) );
  INV_X1 NOT_859( .ZN(g6330), .A(I8070) );
  INV_X1 NOT_860( .ZN(g1721), .A(I2721) );
  INV_X1 NOT_861( .ZN(I5091), .A(g3242) );
  INV_X1 NOT_862( .ZN(I8056), .A(g6109) );
  INV_X1 NOT_863( .ZN(g2932), .A(g1998) );
  INV_X1 NOT_864( .ZN(I8456), .A(g6417) );
  INV_X1 NOT_865( .ZN(g5903), .A(g5753) );
  INV_X1 NOT_866( .ZN(I3833), .A(g2266) );
  INV_X1 NOT_867( .ZN(I2318), .A(g1236) );
  INV_X1 NOT_868( .ZN(g4715), .A(I6327) );
  INV_X1 NOT_869( .ZN(I2367), .A(g1161) );
  INV_X1 NOT_870( .ZN(I1924), .A(g663) );
  INV_X1 NOT_871( .ZN(g6800), .A(I8966) );
  INV_X1 NOT_872( .ZN(I5169), .A(g3593) );
  INV_X1 NOT_873( .ZN(I6410), .A(g4473) );
  INV_X1 NOT_874( .ZN(g4098), .A(I5376) );
  INV_X1 NOT_875( .ZN(g3500), .A(g2647) );
  INV_X1 NOT_876( .ZN(g4498), .A(I6012) );
  INV_X1 NOT_877( .ZN(I2057), .A(g685) );
  INV_X1 NOT_878( .ZN(g1502), .A(g709) );
  INV_X1 NOT_879( .ZN(I5059), .A(g3259) );
  INV_X1 NOT_880( .ZN(I5920), .A(g4228) );
  INV_X1 NOT_881( .ZN(I2457), .A(g1253) );
  INV_X1 NOT_882( .ZN(I3584), .A(g1678) );
  INV_X1 NOT_883( .ZN(I5868), .A(g3864) );
  INV_X1 NOT_884( .ZN(I2989), .A(g1519) );
  INV_X1 NOT_885( .ZN(I2193), .A(g693) );
  INV_X1 NOT_886( .ZN(g5436), .A(I7116) );
  INV_X1 NOT_887( .ZN(g3384), .A(g2834) );
  INV_X1 NOT_888( .ZN(g1940), .A(I3047) );
  INV_X1 NOT_889( .ZN(g2576), .A(I3687) );
  INV_X1 NOT_890( .ZN(g2866), .A(g1905) );
  INV_X1 NOT_891( .ZN(g5135), .A(I6783) );
  INV_X1 NOT_892( .ZN(g2716), .A(I3871) );
  INV_X1 NOT_893( .ZN(g3838), .A(I5037) );
  INV_X1 NOT_894( .ZN(I7906), .A(g5912) );
  INV_X1 NOT_895( .ZN(I3268), .A(g1656) );
  INV_X1 NOT_896( .ZN(I3019), .A(g1755) );
  INV_X1 NOT_897( .ZN(g3424), .A(I4671) );
  INV_X1 NOT_898( .ZN(g5382), .A(I7042) );
  INV_X1 NOT_899( .ZN(I5793), .A(g3803) );
  INV_X1 NOT_900( .ZN(I3419), .A(g1287) );
  INV_X1 NOT_901( .ZN(g6902), .A(I9173) );
  INV_X1 NOT_902( .ZN(I6143), .A(g4237) );
  INV_X1 NOT_903( .ZN(I6343), .A(g4458) );
  INV_X1 NOT_904( .ZN(g846), .A(g586) );
  INV_X1 NOT_905( .ZN(g1671), .A(g985) );
  INV_X1 NOT_906( .ZN(g5805), .A(I7604) );
  INV_X1 NOT_907( .ZN(I5415), .A(g3723) );
  INV_X1 NOT_908( .ZN(g6512), .A(I8456) );
  INV_X1 NOT_909( .ZN(I3452), .A(g1450) );
  INV_X1 NOT_910( .ZN(g4162), .A(I5562) );
  INV_X1 NOT_911( .ZN(g5022), .A(I6666) );
  INV_X1 NOT_912( .ZN(g1030), .A(I2057) );
  INV_X1 NOT_913( .ZN(I8279), .A(g6307) );
  INV_X1 NOT_914( .ZN(g3231), .A(I4492) );
  INV_X1 NOT_915( .ZN(g6490), .A(g6371) );
  INV_X1 NOT_916( .ZN(I2321), .A(g898) );
  INV_X1 NOT_917( .ZN(g6823), .A(I9002) );
  INV_X1 NOT_918( .ZN(g3477), .A(g2692) );
  INV_X1 NOT_919( .ZN(g6166), .A(I7892) );
  INV_X1 NOT_920( .ZN(g6366), .A(I8162) );
  INV_X1 NOT_921( .ZN(I6334), .A(g4454) );
  INV_X1 NOT_922( .ZN(I8872), .A(g6695) );
  INV_X1 NOT_923( .ZN(g2241), .A(I3370) );
  INV_X1 NOT_924( .ZN(g1564), .A(g1030) );
  INV_X1 NOT_925( .ZN(I7892), .A(g5916) );
  INV_X4 NOT_926( .ZN(I3086), .A(g1439) );
  INV_X4 NOT_927( .ZN(g6529), .A(I8503) );
  INV_X1 NOT_928( .ZN(I8843), .A(g6658) );
  INV_X1 NOT_929( .ZN(g6649), .A(I8745) );
  INV_X1 NOT_930( .ZN(I6555), .A(g4703) );
  INV_X1 NOT_931( .ZN(g1741), .A(I2753) );
  INV_X1 NOT_932( .ZN(I6792), .A(g5097) );
  INV_X1 NOT_933( .ZN(g3104), .A(I4351) );
  INV_X1 NOT_934( .ZN(I3385), .A(g1318) );
  INV_X1 NOT_935( .ZN(g2524), .A(I3647) );
  INV_X1 NOT_936( .ZN(g2644), .A(I3788) );
  INV_X1 NOT_937( .ZN(I8834), .A(g6661) );
  INV_X1 NOT_938( .ZN(g6698), .A(I8812) );
  INV_X1 NOT_939( .ZN(g1638), .A(g754) );
  INV_X1 NOT_940( .ZN(g839), .A(g567) );
  INV_X1 NOT_941( .ZN(I6621), .A(g4745) );
  INV_X1 NOT_942( .ZN(g2119), .A(g1391) );
  INV_X1 NOT_943( .ZN(I5502), .A(g3853) );
  INV_X1 NOT_944( .ZN(g1108), .A(I2134) );
  INV_X1 NOT_945( .ZN(I3025), .A(g1439) );
  INV_X1 NOT_946( .ZN(I2552), .A(g971) );
  INV_X1 NOT_947( .ZN(g5437), .A(I7119) );
  INV_X1 NOT_948( .ZN(g4385), .A(I5862) );
  INV_X1 NOT_949( .ZN(I3425), .A(g1274) );
  INV_X1 NOT_950( .ZN(I9092), .A(g6855) );
  INV_X1 NOT_951( .ZN(I4441), .A(g2109) );
  INV_X1 NOT_952( .ZN(g2818), .A(g2464) );
  INV_X1 NOT_953( .ZN(g2867), .A(g1908) );
  INV_X1 NOT_954( .ZN(g1883), .A(g1797) );
  INV_X1 NOT_955( .ZN(g5579), .A(I7333) );
  INV_X1 NOT_956( .ZN(I7478), .A(g5628) );
  INV_X1 NOT_957( .ZN(g4425), .A(I5926) );
  INV_X4 NOT_958( .ZN(I7035), .A(g5150) );
  INV_X4 NOT_959( .ZN(I5388), .A(g3969) );
  INV_X1 NOT_960( .ZN(I7517), .A(g5593) );
  INV_X1 NOT_961( .ZN(g2893), .A(g1985) );
  INV_X1 NOT_962( .ZN(g5752), .A(I7509) );
  INV_X1 NOT_963( .ZN(I8232), .A(g6332) );
  INV_X1 NOT_964( .ZN(g5917), .A(I7683) );
  INV_X1 NOT_965( .ZN(I6567), .A(g4715) );
  INV_X1 NOT_966( .ZN(g6720), .A(I8854) );
  INV_X1 NOT_967( .ZN(I3678), .A(g1690) );
  INV_X1 NOT_968( .ZN(g2975), .A(I4176) );
  INV_X1 NOT_969( .ZN(I5030), .A(g3242) );
  INV_X1 NOT_970( .ZN(I3331), .A(g1631) );
  INV_X1 NOT_971( .ZN(g1861), .A(I2967) );
  INV_X1 NOT_972( .ZN(g6367), .A(I8165) );
  INV_X1 NOT_973( .ZN(g1048), .A(g492) );
  INV_X1 NOT_974( .ZN(I5430), .A(g3727) );
  INV_X1 NOT_975( .ZN(g2599), .A(I3729) );
  INV_X1 NOT_976( .ZN(g5042), .A(I6672) );
  INV_X1 NOT_977( .ZN(g1711), .A(I2712) );
  INV_X1 NOT_978( .ZN(I3635), .A(g1305) );
  INV_X1 NOT_979( .ZN(g6652), .A(I8752) );
  INV_X1 NOT_980( .ZN(g5442), .A(g5270) );
  INV_X1 NOT_981( .ZN(g1055), .A(g269) );
  INV_X1 NOT_982( .ZN(I2570), .A(g1222) );
  INV_X1 NOT_983( .ZN(I2860), .A(g1177) );
  INV_X1 NOT_984( .ZN(g6057), .A(g5824) );
  INV_X1 NOT_985( .ZN(g4131), .A(I5475) );
  INV_X1 NOT_986( .ZN(I4743), .A(g2594) );
  INV_X1 NOT_987( .ZN(I3105), .A(g1439) );
  INV_X1 NOT_988( .ZN(g2170), .A(I3301) );
  INV_X1 NOT_989( .ZN(g2370), .A(I3522) );
  INV_X1 NOT_990( .ZN(g4406), .A(I5913) );
  INV_X4 NOT_991( .ZN(g6193), .A(g5957) );
  INV_X1 NOT_992( .ZN(g1333), .A(I2352) );
  INV_X1 NOT_993( .ZN(g2125), .A(I3255) );
  INV_X1 NOT_994( .ZN(I8552), .A(g6455) );
  INV_X1 NOT_995( .ZN(g1774), .A(I2817) );
  INV_X1 NOT_996( .ZN(g4766), .A(I6406) );
  INV_X1 NOT_997( .ZN(g4105), .A(I5397) );
  INV_X1 NOT_998( .ZN(g1846), .A(I2940) );
  INV_X1 NOT_999( .ZN(g5054), .A(g4816) );
  INV_X1 NOT_1000( .ZN(g4801), .A(g4487) );
  INV_X1 NOT_1001( .ZN(g6834), .A(g6821) );
  INV_X1 NOT_1002( .ZN(g4487), .A(I5991) );
  INV_X1 NOT_1003( .ZN(I7110), .A(g5291) );
  INV_X1 NOT_1004( .ZN(g3534), .A(I4752) );
  INV_X1 NOT_1005( .ZN(I5910), .A(g3750) );
  INV_X1 NOT_1006( .ZN(g5770), .A(g5645) );
  INV_X1 NOT_1007( .ZN(I3755), .A(g2125) );
  INV_X4 NOT_1008( .ZN(g5296), .A(I6946) );
  INV_X4 NOT_1009( .ZN(I8687), .A(g6568) );
  INV_X1 NOT_1010( .ZN(I6933), .A(g5124) );
  INV_X1 NOT_1011( .ZN(g2544), .A(I3662) );
  INV_X1 NOT_1012( .ZN(g6598), .A(I8662) );
  INV_X1 NOT_1013( .ZN(I5609), .A(g3893) );
  INV_X1 NOT_1014( .ZN(I4474), .A(g3052) );
  INV_X1 NOT_1015( .ZN(I2358), .A(g1176) );
  INV_X1 NOT_1016( .ZN(g3014), .A(I4217) );
  INV_X1 NOT_1017( .ZN(g6121), .A(I7835) );
  INV_X1 NOT_1018( .ZN(I7002), .A(g5308) );
  INV_X1 NOT_1019( .ZN(g766), .A(I1856) );
  INV_X1 NOT_1020( .ZN(g3885), .A(I5124) );
  INV_X1 NOT_1021( .ZN(g4226), .A(g4050) );
  INV_X1 NOT_1022( .ZN(g2106), .A(g1378) );
  INV_X1 NOT_1023( .ZN(g2306), .A(g1743) );
  INV_X1 NOT_1024( .ZN(I3373), .A(g1320) );
  INV_X1 NOT_1025( .ZN(g2790), .A(g2413) );
  INV_X1 NOT_1026( .ZN(g6232), .A(g6048) );
  INV_X1 NOT_1027( .ZN(I5217), .A(g3673) );
  INV_X1 NOT_1028( .ZN(I8570), .A(g6433) );
  INV_X1 NOT_1029( .ZN(I8860), .A(g6699) );
  INV_X1 NOT_1030( .ZN(I4480), .A(g3073) );
  INV_X1 NOT_1031( .ZN(g1994), .A(I3105) );
  INV_X1 NOT_1032( .ZN(g1290), .A(I2275) );
  INV_X1 NOT_1033( .ZN(I2275), .A(g909) );
  INV_X1 NOT_1034( .ZN(g6938), .A(I9227) );
  INV_X1 NOT_1035( .ZN(I5466), .A(g3787) );
  INV_X1 NOT_1036( .ZN(g4173), .A(I5577) );
  INV_X1 NOT_1037( .ZN(I8710), .A(g6517) );
  INV_X1 NOT_1038( .ZN(g2461), .A(I3593) );
  INV_X1 NOT_1039( .ZN(I7590), .A(g5605) );
  INV_X1 NOT_1040( .ZN(I3602), .A(g1491) );
  INV_X1 NOT_1041( .ZN(I3007), .A(g1439) );
  INV_X1 NOT_1042( .ZN(g2756), .A(g2353) );
  INV_X1 NOT_1043( .ZN(g2622), .A(I3764) );
  INV_X1 NOT_1044( .ZN(I3059), .A(g1519) );
  INV_X1 NOT_1045( .ZN(I3578), .A(g1484) );
  INV_X1 NOT_1046( .ZN(I3868), .A(g2125) );
  INV_X1 NOT_1047( .ZN(g5888), .A(g5731) );
  INV_X1 NOT_1048( .ZN(g1256), .A(g838) );
  INV_X4 NOT_1049( .ZN(g6519), .A(I8473) );
  INV_X1 NOT_1050( .ZN(I6289), .A(g4433) );
  INV_X1 NOT_1051( .ZN(I9024), .A(g6803) );
  INV_X1 NOT_1052( .ZN(I5448), .A(g3960) );
  INV_X1 NOT_1053( .ZN(I3767), .A(g2125) );
  INV_X1 NOT_1054( .ZN(g5787), .A(g5685) );
  INV_X1 NOT_1055( .ZN(g2904), .A(g1991) );
  INV_X1 NOT_1056( .ZN(g6552), .A(I8552) );
  INV_X1 NOT_1057( .ZN(g6606), .A(I8684) );
  INV_X1 NOT_1058( .ZN(g2446), .A(I3581) );
  INV_X1 NOT_1059( .ZN(I5333), .A(g3491) );
  INV_X1 NOT_1060( .ZN(I2284), .A(g922) );
  INV_X1 NOT_1061( .ZN(g1381), .A(I2417) );
  INV_X1 NOT_1062( .ZN(g4718), .A(I6334) );
  INV_X1 NOT_1063( .ZN(g4767), .A(g4601) );
  INV_X1 NOT_1064( .ZN(I3261), .A(g1783) );
  INV_X1 NOT_1065( .ZN(g1847), .A(I2943) );
  INV_X1 NOT_1066( .ZN(I4688), .A(g3207) );
  INV_X1 NOT_1067( .ZN(I5774), .A(g3807) );
  INV_X1 NOT_1068( .ZN(I9077), .A(g6845) );
  INV_X1 NOT_1069( .ZN(I8659), .A(g6523) );
  INV_X1 NOT_1070( .ZN(g4535), .A(g4173) );
  INV_X1 NOT_1071( .ZN(I4976), .A(g3575) );
  INV_X1 NOT_1072( .ZN(g1685), .A(I2671) );
  INV_X1 NOT_1073( .ZN(g2145), .A(I3268) );
  INV_X1 NOT_1074( .ZN(I8506), .A(g6483) );
  INV_X1 NOT_1075( .ZN(g2841), .A(g2541) );
  INV_X1 NOT_1076( .ZN(g4582), .A(g4210) );
  INV_X1 NOT_1077( .ZN(g3022), .A(I4229) );
  INV_X1 NOT_1078( .ZN(g2391), .A(I3534) );
  INV_X1 NOT_1079( .ZN(g6586), .A(I8626) );
  INV_X1 NOT_1080( .ZN(g952), .A(I2029) );
  INV_X1 NOT_1081( .ZN(g1263), .A(g846) );
  INV_X1 NOT_1082( .ZN(g964), .A(g357) );
  INV_X1 NOT_1083( .ZN(I2420), .A(g791) );
  INV_X1 NOT_1084( .ZN(g2695), .A(I3843) );
  INV_X4 NOT_1085( .ZN(g2637), .A(I3779) );
  INV_X4 NOT_1086( .ZN(g1950), .A(I3059) );
  INV_X4 NOT_1087( .ZN(g5138), .A(I6792) );
  INV_X1 NOT_1088( .ZN(g4227), .A(g4059) );
  INV_X1 NOT_1089( .ZN(I7295), .A(g5439) );
  INV_X1 NOT_1090( .ZN(g5791), .A(I7590) );
  INV_X1 NOT_1091( .ZN(g3798), .A(g3388) );
  INV_X1 NOT_1092( .ZN(I9104), .A(g6864) );
  INV_X1 NOT_1093( .ZN(g5309), .A(g5063) );
  INV_X1 NOT_1094( .ZN(g2159), .A(I3284) );
  INV_X1 NOT_1095( .ZN(g6570), .A(I8594) );
  INV_X1 NOT_1096( .ZN(g4246), .A(I5692) );
  INV_X1 NOT_1097( .ZN(I6132), .A(g4219) );
  INV_X1 NOT_1098( .ZN(I8174), .A(g6173) );
  INV_X1 NOT_1099( .ZN(g6525), .A(I8491) );
  INV_X1 NOT_1100( .ZN(g6710), .A(I8840) );
  INV_X1 NOT_1101( .ZN(I5418), .A(g4036) );
  INV_X1 NOT_1102( .ZN(I6680), .A(g4713) );
  INV_X1 NOT_1103( .ZN(g4721), .A(I6343) );
  INV_X1 NOT_1104( .ZN(g1631), .A(I2588) );
  INV_X1 NOT_1105( .ZN(g2416), .A(I3556) );
  INV_X1 NOT_1106( .ZN(g3095), .A(I4340) );
  INV_X1 NOT_1107( .ZN(g3037), .A(I4252) );
  INV_X1 NOT_1108( .ZN(I3502), .A(g1295) );
  INV_X1 NOT_1109( .ZN(g1257), .A(g845) );
  INV_X1 NOT_1110( .ZN(g1101), .A(I2125) );
  INV_X1 NOT_1111( .ZN(I2204), .A(g694) );
  INV_X1 NOT_1112( .ZN(I2630), .A(g1143) );
  INV_X1 NOT_1113( .ZN(I5493), .A(g3834) );
  INV_X1 NOT_1114( .ZN(I8180), .A(g6176) );
  INV_X1 NOT_1115( .ZN(I4220), .A(g2164) );
  INV_X1 NOT_1116( .ZN(I7966), .A(g6166) );
  INV_X1 NOT_1117( .ZN(I8591), .A(g6448) );
  INV_X1 NOT_1118( .ZN(g2315), .A(I3465) );
  INV_X1 NOT_1119( .ZN(g5957), .A(g5866) );
  INV_X1 NOT_1120( .ZN(g6879), .A(I9104) );
  INV_X1 NOT_1121( .ZN(g6607), .A(I8687) );
  INV_X1 NOT_1122( .ZN(I6558), .A(g4705) );
  INV_X1 NOT_1123( .ZN(g4502), .A(I6020) );
  INV_X1 NOT_1124( .ZN(g5049), .A(I6685) );
  INV_X1 NOT_1125( .ZN(I9044), .A(g6836) );
  INV_X1 NOT_1126( .ZN(g927), .A(I1958) );
  INV_X1 NOT_1127( .ZN(I1942), .A(g664) );
  INV_X1 NOT_1128( .ZN(I4023), .A(g2315) );
  INV_X1 NOT_1129( .ZN(g3719), .A(g3053) );
  INV_X1 NOT_1130( .ZN(g6506), .A(I8438) );
  INV_X1 NOT_1131( .ZN(g5575), .A(g5411) );
  INV_X1 NOT_1132( .ZN(I8420), .A(g6422) );
  INV_X1 NOT_1133( .ZN(I3388), .A(g1324) );
  INV_X1 NOT_1134( .ZN(g2874), .A(g1849) );
  INV_X1 NOT_1135( .ZN(g3752), .A(I4935) );
  INV_X1 NOT_1136( .ZN(I5397), .A(g3932) );
  INV_X1 NOT_1137( .ZN(I3028), .A(g1504) );
  INV_X1 NOT_1138( .ZN(g4188), .A(I5594) );
  INV_X1 NOT_1139( .ZN(g6587), .A(I8629) );
  INV_X1 NOT_1140( .ZN(g4388), .A(I5871) );
  INV_X1 NOT_1141( .ZN(I5421), .A(g3724) );
  INV_X1 NOT_1142( .ZN(I3428), .A(g1825) );
  INV_X1 NOT_1143( .ZN(I2973), .A(g1687) );
  INV_X1 NOT_1144( .ZN(I7254), .A(g5458) );
  INV_X1 NOT_1145( .ZN(I7814), .A(g5922) );
  INV_X1 NOT_1146( .ZN(I3247), .A(g1791) );
  INV_X2 NOT_1147( .ZN(g3042), .A(I4261) );
  INV_X2 NOT_1148( .ZN(g6615), .A(I8707) );
  INV_X2 NOT_1149( .ZN(I7150), .A(g5355) );
  INV_X1 NOT_1150( .ZN(I4327), .A(g2525) );
  INV_X1 NOT_1151( .ZN(g4428), .A(I5933) );
  INV_X1 NOT_1152( .ZN(g3786), .A(g3388) );
  INV_X1 NOT_1153( .ZN(g5584), .A(I7346) );
  INV_X1 NOT_1154( .ZN(g5539), .A(g5331) );
  INV_X1 NOT_1155( .ZN(g5896), .A(g5753) );
  INV_X1 NOT_1156( .ZN(g1673), .A(I2653) );
  INV_X1 NOT_1157( .ZN(g6374), .A(I8186) );
  INV_X1 NOT_1158( .ZN(I3826), .A(g2145) );
  INV_X1 NOT_1159( .ZN(g3364), .A(g3114) );
  INV_X1 NOT_1160( .ZN(g3233), .A(I4498) );
  INV_X1 NOT_1161( .ZN(I8515), .A(g6492) );
  INV_X1 NOT_1162( .ZN(g4564), .A(g4192) );
  INV_X1 NOT_1163( .ZN(g3054), .A(I4279) );
  INV_X1 NOT_1164( .ZN(I5562), .A(g4002) );
  INV_X1 NOT_1165( .ZN(I4303), .A(g1897) );
  INV_X1 NOT_1166( .ZN(g2612), .A(I3752) );
  INV_X1 NOT_1167( .ZN(I8300), .A(g6299) );
  INV_X1 NOT_1168( .ZN(g6284), .A(I8002) );
  INV_X1 NOT_1169( .ZN(g2243), .A(I3376) );
  INV_X1 NOT_1170( .ZN(g3770), .A(I4961) );
  INV_X1 NOT_1171( .ZN(I9014), .A(g6820) );
  INV_X1 NOT_1172( .ZN(I3638), .A(g1484) );
  INV_X1 NOT_1173( .ZN(g1772), .A(I2811) );
  INV_X1 NOT_1174( .ZN(I5723), .A(g3942) );
  INV_X1 NOT_1175( .ZN(g4741), .A(I6371) );
  INV_X1 NOT_1176( .ZN(g6591), .A(I8641) );
  INV_X1 NOT_1177( .ZN(g5052), .A(I6692) );
  INV_X1 NOT_1178( .ZN(g6832), .A(I9021) );
  INV_X1 NOT_1179( .ZN(g4910), .A(I6612) );
  INV_X1 NOT_1180( .ZN(I2648), .A(g980) );
  INV_X1 NOT_1181( .ZN(g2234), .A(I3367) );
  INV_X1 NOT_1182( .ZN(g6853), .A(I9082) );
  INV_X1 NOT_1183( .ZN(g1890), .A(g1359) );
  INV_X1 NOT_1184( .ZN(I3883), .A(g2574) );
  INV_X1 NOT_1185( .ZN(g6420), .A(I8270) );
  INV_X1 NOT_1186( .ZN(I4240), .A(g2165) );
  INV_X1 NOT_1187( .ZN(g2330), .A(g1777) );
  INV_X1 NOT_1188( .ZN(g4108), .A(I5406) );
  INV_X1 NOT_1189( .ZN(g4609), .A(I6182) );
  INV_X1 NOT_1190( .ZN(g6507), .A(I8441) );
  INV_X1 NOT_1191( .ZN(g4308), .A(I5777) );
  INV_X1 NOT_1192( .ZN(g1011), .A(I2050) );
  INV_X1 NOT_1193( .ZN(g1734), .A(g952) );
  INV_X1 NOT_1194( .ZN(I3758), .A(g2041) );
  INV_X1 NOT_1195( .ZN(g5086), .A(g4732) );
  INV_X1 NOT_1196( .ZN(g897), .A(g41) );
  INV_X1 NOT_1197( .ZN(I8040), .A(g6142) );
  INV_X1 NOT_1198( .ZN(g951), .A(g84) );
  INV_X1 NOT_1199( .ZN(I8969), .A(g6797) );
  INV_X1 NOT_1200( .ZN(g2800), .A(g2430) );
  INV_X1 NOT_1201( .ZN(g5730), .A(I7497) );
  INV_X1 NOT_1202( .ZN(g2554), .A(I3669) );
  INV_X1 NOT_1203( .ZN(g4758), .A(I6382) );
  INV_X1 NOT_1204( .ZN(I2839), .A(g1123) );
  INV_X1 NOT_1205( .ZN(I3861), .A(g1834) );
  INV_X1 NOT_1206( .ZN(g6905), .A(I9182) );
  INV_X1 NOT_1207( .ZN(g3029), .A(I4240) );
  INV_X1 NOT_1208( .ZN(I3711), .A(g1848) );
  INV_X1 NOT_1209( .ZN(I9182), .A(g6879) );
  INV_X1 NOT_1210( .ZN(g3787), .A(I4986) );
  INV_X1 NOT_1211( .ZN(g2213), .A(I3346) );
  INV_X2 NOT_1212( .ZN(g5897), .A(g5731) );
  INV_X2 NOT_1213( .ZN(g5025), .A(g4814) );
  INV_X2 NOT_1214( .ZN(g6515), .A(g6408) );
  INV_X1 NOT_1215( .ZN(g4861), .A(I6587) );
  INV_X1 NOT_1216( .ZN(g5425), .A(I7091) );
  INV_X1 NOT_1217( .ZN(I4347), .A(g2555) );
  INV_X1 NOT_1218( .ZN(I2172), .A(g691) );
  INV_X1 NOT_1219( .ZN(I2278), .A(g917) );
  INV_X1 NOT_1220( .ZN(g4711), .A(I6315) );
  INV_X1 NOT_1221( .ZN(g6100), .A(I7796) );
  INV_X1 NOT_1222( .ZN(I4681), .A(g2947) );
  INV_X1 NOT_1223( .ZN(g1480), .A(g985) );
  INV_X1 NOT_1224( .ZN(g2902), .A(g1899) );
  INV_X1 NOT_1225( .ZN(I8875), .A(g6697) );
  INV_X1 NOT_1226( .ZN(I2143), .A(g2) );
  INV_X1 NOT_1227( .ZN(I2343), .A(g1177) );
  INV_X1 NOT_1228( .ZN(I6139), .A(g4222) );
  INV_X1 NOT_1229( .ZN(g4133), .A(I5481) );
  INV_X1 NOT_1230( .ZN(g3297), .A(g3046) );
  INV_X1 NOT_1231( .ZN(g2512), .A(I3638) );
  INV_X1 NOT_1232( .ZN(g2090), .A(I3206) );
  INV_X1 NOT_1233( .ZN(g4846), .A(I6546) );
  INV_X1 NOT_1234( .ZN(I2134), .A(g705) );
  INV_X1 NOT_1235( .ZN(I6795), .A(g5022) );
  INV_X1 NOT_1236( .ZN(I6737), .A(g4662) );
  INV_X1 NOT_1237( .ZN(I2334), .A(g1193) );
  INV_X1 NOT_1238( .ZN(I6809), .A(g5051) );
  INV_X1 NOT_1239( .ZN(I5743), .A(g4022) );
  INV_X1 NOT_1240( .ZN(g5331), .A(I6995) );
  INV_X1 NOT_1241( .ZN(I5890), .A(g3878) );
  INV_X1 NOT_1242( .ZN(I3509), .A(g1461) );
  INV_X1 NOT_1243( .ZN(g3963), .A(I5217) );
  INV_X1 NOT_1244( .ZN(g3791), .A(g3388) );
  INV_X1 NOT_1245( .ZN(I8884), .A(g6704) );
  INV_X1 NOT_1246( .ZN(I5505), .A(g3860) );
  INV_X1 NOT_1247( .ZN(g1688), .A(I2688) );
  INV_X1 NOT_1248( .ZN(I6672), .A(g4752) );
  INV_X1 NOT_1249( .ZN(g4780), .A(I6434) );
  INV_X1 NOT_1250( .ZN(g6040), .A(g5824) );
  INV_X1 NOT_1251( .ZN(g1857), .A(I2961) );
  INV_X1 NOT_1252( .ZN(I6231), .A(g4350) );
  INV_X1 NOT_1253( .ZN(I3662), .A(g1688) );
  INV_X1 NOT_1254( .ZN(g4509), .A(I6039) );
  INV_X1 NOT_1255( .ZN(g5087), .A(g4736) );
  INV_X1 NOT_1256( .ZN(I9095), .A(g6855) );
  INV_X1 NOT_1257( .ZN(g5801), .A(I7600) );
  INV_X1 NOT_1258( .ZN(g2155), .A(I3274) );
  INV_X1 NOT_1259( .ZN(I9208), .A(g6922) );
  INV_X1 NOT_1260( .ZN(g4662), .A(g4640) );
  INV_X1 NOT_1261( .ZN(I3093), .A(g1426) );
  INV_X1 NOT_1262( .ZN(g965), .A(I2033) );
  INV_X1 NOT_1263( .ZN(I3493), .A(g1461) );
  INV_X1 NOT_1264( .ZN(I3816), .A(g2580) );
  INV_X1 NOT_1265( .ZN(g1326), .A(g894) );
  INV_X1 NOT_1266( .ZN(I8235), .A(g6312) );
  INV_X1 NOT_1267( .ZN(I6099), .A(g4398) );
  INV_X1 NOT_1268( .ZN(I8282), .A(g6309) );
  INV_X2 NOT_1269( .ZN(g3049), .A(I4270) );
  INV_X2 NOT_1270( .ZN(g6528), .A(I8500) );
  INV_X2 NOT_1271( .ZN(g1760), .A(I2785) );
  INV_X2 NOT_1272( .ZN(g4493), .A(I6001) );
  INV_X1 NOT_1273( .ZN(g6351), .A(I8107) );
  INV_X1 NOT_1274( .ZN(I1850), .A(g210) );
  INV_X1 NOT_1275( .ZN(g6875), .A(I9092) );
  INV_X1 NOT_1276( .ZN(g834), .A(g341) );
  INV_X1 NOT_1277( .ZN(I8988), .A(g6787) );
  INV_X1 NOT_1278( .ZN(g6530), .A(I8506) );
  INV_X1 NOT_1279( .ZN(g3575), .A(I4777) );
  INV_X1 NOT_1280( .ZN(g5045), .A(I6677) );
  INV_X1 NOT_1281( .ZN(I8693), .A(g6570) );
  INV_X1 NOT_1282( .ZN(g6655), .A(I8761) );
  INV_X1 NOT_1283( .ZN(g5445), .A(g5274) );
  INV_X1 NOT_1284( .ZN(I5713), .A(g4022) );
  INV_X1 NOT_1285( .ZN(g3604), .A(I4799) );
  INV_X1 NOT_1286( .ZN(I8548), .A(g6454) );
  INV_X1 NOT_1287( .ZN(g5491), .A(I7193) );
  INV_X1 NOT_1288( .ZN(g3498), .A(g2634) );
  INV_X1 NOT_1289( .ZN(g4381), .A(I5854) );
  INV_X1 NOT_1290( .ZN(g4847), .A(I6549) );
  INV_X1 NOT_1291( .ZN(g2118), .A(I3247) );
  INV_X1 NOT_1292( .ZN(g2619), .A(I3761) );
  INV_X1 NOT_1293( .ZN(I8555), .A(g6456) );
  INV_X1 NOT_1294( .ZN(g2367), .A(I3519) );
  INV_X1 NOT_1295( .ZN(g2872), .A(g1922) );
  INV_X1 NOT_1296( .ZN(g1608), .A(I2570) );
  INV_X1 NOT_1297( .ZN(g1220), .A(I2221) );
  INV_X1 NOT_1298( .ZN(g4700), .A(I6292) );
  INV_X1 NOT_1299( .ZN(g6410), .A(I8240) );
  INV_X1 NOT_1300( .ZN(I9164), .A(g6885) );
  INV_X1 NOT_1301( .ZN(g4397), .A(I5890) );
  INV_X1 NOT_1302( .ZN(I9233), .A(g6938) );
  INV_X1 NOT_1303( .ZN(I2776), .A(g1192) );
  INV_X1 NOT_1304( .ZN(I7640), .A(g5773) );
  INV_X1 NOT_1305( .ZN(g5407), .A(I7073) );
  INV_X1 NOT_1306( .ZN(g6884), .A(I9119) );
  INV_X1 NOT_1307( .ZN(I2593), .A(g1177) );
  INV_X1 NOT_1308( .ZN(g5059), .A(I6697) );
  INV_X1 NOT_1309( .ZN(g5920), .A(I7692) );
  INV_X1 NOT_1310( .ZN(g6839), .A(I9038) );
  INV_X1 NOT_1311( .ZN(g2457), .A(I3587) );
  INV_X1 NOT_1312( .ZN(g5578), .A(g5425) );
  INV_X1 NOT_1313( .ZN(I6444), .A(g4503) );
  INV_X1 NOT_1314( .ZN(I6269), .A(g4655) );
  INV_X1 NOT_1315( .ZN(g1423), .A(I2442) );
  INV_X1 NOT_1316( .ZN(g923), .A(g332) );
  INV_X1 NOT_1317( .ZN(I5857), .A(g3740) );
  INV_X1 NOT_1318( .ZN(I7176), .A(g5437) );
  INV_X2 NOT_1319( .ZN(g1588), .A(g798) );
  INV_X2 NOT_1320( .ZN(I8113), .A(g6147) );
  INV_X2 NOT_1321( .ZN(g5582), .A(I7342) );
  INV_X2 NOT_1322( .ZN(g1161), .A(I2182) );
  INV_X1 NOT_1323( .ZN(g6278), .A(I7966) );
  INV_X1 NOT_1324( .ZN(g2686), .A(I3830) );
  INV_X1 NOT_1325( .ZN(g6372), .A(I8180) );
  INV_X1 NOT_1326( .ZN(g3162), .A(I4402) );
  INV_X1 NOT_1327( .ZN(g5261), .A(I6918) );
  INV_X1 NOT_1328( .ZN(g3019), .A(I4226) );
  INV_X1 NOT_1329( .ZN(I4294), .A(g2525) );
  INV_X1 NOT_1330( .ZN(I6543), .A(g4718) );
  INV_X1 NOT_1331( .ZN(g6618), .A(I8716) );
  INV_X1 NOT_1332( .ZN(g1665), .A(g985) );
  INV_X1 NOT_1333( .ZN(I7829), .A(g5926) );
  INV_X1 NOT_1334( .ZN(I3723), .A(g2158) );
  INV_X1 NOT_1335( .ZN(g6143), .A(I7865) );
  INV_X1 NOT_1336( .ZN(g4562), .A(I6132) );
  INV_X1 NOT_1337( .ZN(g6235), .A(g6062) );
  INV_X1 NOT_1338( .ZN(g2598), .A(I3726) );
  INV_X1 NOT_1339( .ZN(g3052), .A(I4273) );
  INV_X1 NOT_1340( .ZN(g1327), .A(I2334) );
  INV_X1 NOT_1341( .ZN(I2521), .A(g1063) );
  INV_X1 NOT_1342( .ZN(I3301), .A(g1730) );
  INV_X1 NOT_1343( .ZN(g5415), .A(I7081) );
  INV_X1 NOT_1344( .ZN(g3452), .A(g2625) );
  INV_X1 NOT_1345( .ZN(g6282), .A(I7996) );
  INV_X1 NOT_1346( .ZN(I2050), .A(g683) );
  INV_X1 NOT_1347( .ZN(I5400), .A(g3963) );
  INV_X1 NOT_1348( .ZN(g6566), .A(I8582) );
  INV_X1 NOT_1349( .ZN(I8494), .A(g6428) );
  INV_X1 NOT_1350( .ZN(I4501), .A(g2705) );
  INV_X1 NOT_1351( .ZN(I6534), .A(g4706) );
  INV_X1 NOT_1352( .ZN(I8518), .A(g6494) );
  INV_X1 NOT_1353( .ZN(I3605), .A(g1681) );
  INV_X1 NOT_1354( .ZN(g4723), .A(I6349) );
  INV_X1 NOT_1355( .ZN(I8567), .A(g6432) );
  INV_X1 NOT_1356( .ZN(g4101), .A(I5385) );
  INV_X1 NOT_1357( .ZN(g6134), .A(I7852) );
  INV_X1 NOT_1358( .ZN(g5664), .A(g5521) );
  INV_X1 NOT_1359( .ZN(g2625), .A(I3767) );
  INV_X1 NOT_1360( .ZN(I7270), .A(g5352) );
  INV_X1 NOT_1361( .ZN(g2232), .A(I3361) );
  INV_X1 NOT_1362( .ZN(g6548), .A(I8548) );
  INV_X1 NOT_1363( .ZN(I6927), .A(g5124) );
  INV_X1 NOT_1364( .ZN(g3086), .A(I4327) );
  INV_X1 NOT_1365( .ZN(I2724), .A(g1220) );
  INV_X1 NOT_1366( .ZN(g2253), .A(I3388) );
  INV_X1 NOT_1367( .ZN(I2179), .A(g293) );
  INV_X1 NOT_1368( .ZN(g3486), .A(g2869) );
  INV_X1 NOT_1369( .ZN(g2813), .A(g2457) );
  INV_X1 NOT_1370( .ZN(I2379), .A(g1123) );
  INV_X1 NOT_1371( .ZN(g1696), .A(I2700) );
  INV_X1 NOT_1372( .ZN(I7073), .A(g5281) );
  INV_X1 NOT_1373( .ZN(I7796), .A(g5917) );
  INV_X1 NOT_1374( .ZN(I6885), .A(g4872) );
  INV_X1 NOT_1375( .ZN(I6414), .A(g4497) );
  INV_X1 NOT_1376( .ZN(g3504), .A(g2675) );
  INV_X1 NOT_1377( .ZN(I6946), .A(g5124) );
  INV_X1 NOT_1378( .ZN(g1732), .A(I2738) );
  INV_X1 NOT_1379( .ZN(g3881), .A(I5116) );
  INV_X1 NOT_1380( .ZN(g2740), .A(I3909) );
  INV_X1 NOT_1381( .ZN(I2658), .A(g1001) );
  INV_X1 NOT_1382( .ZN(I3441), .A(g1502) );
  INV_X2 NOT_1383( .ZN(I7069), .A(g5281) );
  INV_X2 NOT_1384( .ZN(g3070), .A(I4297) );
  INV_X2 NOT_1385( .ZN(I8264), .A(g6296) );
  INV_X2 NOT_1386( .ZN(g6621), .A(I8721) );
  INV_X1 NOT_1387( .ZN(I2835), .A(g1209) );
  INV_X1 NOT_1388( .ZN(I7469), .A(g5625) );
  INV_X1 NOT_1389( .ZN(g3897), .A(g3251) );
  INV_X1 NOT_1390( .ZN(I5023), .A(g3263) );
  INV_X1 NOT_1391( .ZN(g1472), .A(g952) );
  INV_X1 NOT_1392( .ZN(g1043), .A(g486) );
  INV_X1 NOT_1393( .ZN(I5977), .A(g4319) );
  INV_X1 NOT_1394( .ZN(I8521), .A(g6495) );
  INV_X1 NOT_1395( .ZN(I6036), .A(g4370) );
  INV_X1 NOT_1396( .ZN(I8641), .A(g6524) );
  INV_X1 NOT_1397( .ZN(I2611), .A(g1209) );
  INV_X1 NOT_1398( .ZN(g893), .A(g23) );
  INV_X1 NOT_1399( .ZN(g2687), .A(I3833) );
  INV_X1 NOT_1400( .ZN(I8450), .A(g6412) );
  INV_X1 NOT_1401( .ZN(I3669), .A(g1739) );
  INV_X1 NOT_1402( .ZN(g1116), .A(I2154) );
  INV_X1 NOT_1403( .ZN(g2586), .A(I3711) );
  INV_X1 NOT_1404( .ZN(I3531), .A(g1593) );
  INV_X1 NOT_1405( .ZN(I5451), .A(g3967) );
  INV_X1 NOT_1406( .ZN(I6182), .A(g4249) );
  INV_X1 NOT_1407( .ZN(g6518), .A(I8470) );
  INV_X1 NOT_1408( .ZN(g6567), .A(I8585) );
  INV_X1 NOT_1409( .ZN(I8724), .A(g6533) );
  INV_X1 NOT_1410( .ZN(I6382), .A(g4460) );
  INV_X1 NOT_1411( .ZN(g996), .A(I2041) );
  INV_X1 NOT_1412( .ZN(g3331), .A(g3076) );
  INV_X1 NOT_1413( .ZN(I3890), .A(g2145) );
  INV_X1 NOT_1414( .ZN(g4772), .A(I6420) );
  INV_X1 NOT_1415( .ZN(g5247), .A(g4900) );
  INV_X1 NOT_1416( .ZN(g4531), .A(I6105) );
  INV_X1 NOT_1417( .ZN(I5633), .A(g3768) );
  INV_X1 NOT_1418( .ZN(I8878), .A(g6710) );
  INV_X1 NOT_1419( .ZN(g1681), .A(I2663) );
  INV_X1 NOT_1420( .ZN(I3505), .A(g1305) );
  INV_X1 NOT_1421( .ZN(g6593), .A(I8647) );
  INV_X1 NOT_1422( .ZN(g3766), .A(I4955) );
  INV_X1 NOT_1423( .ZN(g1533), .A(g878) );
  INV_X1 NOT_1424( .ZN(g5564), .A(g5382) );
  INV_X1 NOT_1425( .ZN(I5103), .A(g3440) );
  INV_X1 NOT_1426( .ZN(g2525), .A(I3650) );
  INV_X1 NOT_1427( .ZN(g3801), .A(g3388) );
  INV_X1 NOT_1428( .ZN(g3487), .A(g2622) );
  INV_X1 NOT_1429( .ZN(g1914), .A(I3013) );
  INV_X1 NOT_1430( .ZN(I5696), .A(g3942) );
  INV_X1 NOT_1431( .ZN(g2691), .A(g2317) );
  INV_X1 NOT_1432( .ZN(g4011), .A(g3486) );
  INV_X1 NOT_1433( .ZN(I6798), .A(g5042) );
  INV_X1 NOT_1434( .ZN(g4856), .A(I6576) );
  INV_X1 NOT_1435( .ZN(g5741), .A(g5602) );
  INV_X1 NOT_1436( .ZN(I2802), .A(g1204) );
  INV_X1 NOT_1437( .ZN(I3074), .A(g1426) );
  INV_X1 NOT_1438( .ZN(I3474), .A(g1450) );
  INV_X1 NOT_1439( .ZN(I5753), .A(g4022) );
  INV_X1 NOT_1440( .ZN(g5638), .A(I7397) );
  INV_X1 NOT_1441( .ZN(g6160), .A(g5926) );
  INV_X1 NOT_1442( .ZN(g3226), .A(I4477) );
  INV_X1 NOT_1443( .ZN(I5508), .A(g3867) );
  INV_X1 NOT_1444( .ZN(g6360), .A(I8144) );
  INV_X1 NOT_1445( .ZN(g6933), .A(I9220) );
  INV_X1 NOT_1446( .ZN(I5944), .A(g4356) );
  INV_X1 NOT_1447( .ZN(g2962), .A(g2008) );
  INV_X1 NOT_1448( .ZN(g6521), .A(I8479) );
  INV_X1 NOT_1449( .ZN(I9098), .A(g6864) );
  INV_X1 NOT_1450( .ZN(g2158), .A(I3281) );
  INV_X1 NOT_1451( .ZN(I5472), .A(g3846) );
  INV_X1 NOT_1452( .ZN(I8981), .A(g6793) );
  INV_X1 NOT_1453( .ZN(g2506), .A(I3632) );
  INV_X1 NOT_1454( .ZN(I3080), .A(g1519) );
  INV_X1 NOT_1455( .ZN(I8674), .A(g6521) );
  INV_X1 NOT_1456( .ZN(g1820), .A(I2880) );
  INV_X1 NOT_1457( .ZN(I5043), .A(g3247) );
  INV_X1 NOT_1458( .ZN(I6495), .A(g4607) );
  INV_X1 NOT_1459( .ZN(g1936), .A(g1756) );
  INV_X2 NOT_1460( .ZN(I6437), .A(g4501) );
  INV_X2 NOT_1461( .ZN(g3173), .A(I4410) );
  INV_X2 NOT_1462( .ZN(I6102), .A(g4399) );
  INV_X2 NOT_1463( .ZN(I6302), .A(g4440) );
  INV_X1 NOT_1464( .ZN(I8997), .A(g6790) );
  INV_X1 NOT_1465( .ZN(g1117), .A(g32) );
  INV_X1 NOT_1466( .ZN(I8541), .A(g6452) );
  INV_X1 NOT_1467( .ZN(g1317), .A(I2306) );
  INV_X1 NOT_1468( .ZN(g3491), .A(g2608) );
  INV_X1 NOT_1469( .ZN(g2587), .A(I3714) );
  INV_X1 NOT_1470( .ZN(I6579), .A(g4798) );
  INV_X1 NOT_1471( .ZN(I5116), .A(g3259) );
  INV_X1 NOT_1472( .ZN(I7852), .A(g5993) );
  INV_X1 NOT_1473( .ZN(I5316), .A(g3557) );
  INV_X1 NOT_1474( .ZN(g6724), .A(I8866) );
  INV_X1 NOT_1475( .ZN(I3569), .A(g1789) );
  INV_X1 NOT_1476( .ZN(g2111), .A(g1384) );
  INV_X1 NOT_1477( .ZN(g2275), .A(I3422) );
  INV_X1 NOT_1478( .ZN(g5466), .A(I7146) );
  INV_X1 NOT_1479( .ZN(I8332), .A(g6306) );
  INV_X1 NOT_1480( .ZN(g4713), .A(I6321) );
  INV_X1 NOT_1481( .ZN(I7701), .A(g5720) );
  INV_X1 NOT_1482( .ZN(g3369), .A(I4646) );
  INV_X1 NOT_1483( .ZN(I8153), .A(g6185) );
  INV_X1 NOT_1484( .ZN(g3007), .A(g2197) );
  INV_X1 NOT_1485( .ZN(g2615), .A(I3755) );
  INV_X1 NOT_1486( .ZN(g6878), .A(I9101) );
  INV_X1 NOT_1487( .ZN(I2864), .A(g1177) );
  INV_X1 NOT_1488( .ZN(g4569), .A(I6143) );
  INV_X1 NOT_1489( .ZN(g5571), .A(g5395) );
  INV_X1 NOT_1490( .ZN(g5861), .A(g5636) );
  INV_X1 NOT_1491( .ZN(g3868), .A(g3491) );
  INV_X1 NOT_1492( .ZN(g2174), .A(I3313) );
  INV_X1 NOT_1493( .ZN(g3459), .A(g2664) );
  INV_X1 NOT_1494( .ZN(g815), .A(I1877) );
  INV_X1 NOT_1495( .ZN(g1775), .A(g952) );
  INV_X1 NOT_1496( .ZN(g5448), .A(g5278) );
  INV_X1 NOT_1497( .ZN(g1922), .A(I3025) );
  INV_X1 NOT_1498( .ZN(g835), .A(g345) );
  INV_X1 NOT_1499( .ZN(g5711), .A(I7472) );
  INV_X1 NOT_1500( .ZN(g6835), .A(I9028) );
  INV_X1 NOT_1501( .ZN(g1581), .A(g910) );
  INV_X1 NOT_1502( .ZN(g6882), .A(I9113) );
  INV_X1 NOT_1503( .ZN(I6042), .A(g4374) );
  INV_X1 NOT_1504( .ZN(g1060), .A(g107) );
  INV_X1 NOT_1505( .ZN(g2284), .A(I3431) );
  INV_X1 NOT_1506( .ZN(I6786), .A(g4824) );
  INV_X1 NOT_1507( .ZN(g1460), .A(I2457) );
  INV_X1 NOT_1508( .ZN(g5774), .A(I7517) );
  INV_X1 NOT_1509( .ZN(g4857), .A(I6579) );
  INV_X1 NOT_1510( .ZN(g3793), .A(g3491) );
  INV_X1 NOT_1511( .ZN(g6611), .A(I8699) );
  INV_X1 NOT_1512( .ZN(g2591), .A(I3720) );
  INV_X1 NOT_1513( .ZN(g3015), .A(I4220) );
  INV_X1 NOT_1514( .ZN(g3227), .A(I4480) );
  INV_X1 NOT_1515( .ZN(g1739), .A(I2749) );
  INV_X1 NOT_1516( .ZN(I6054), .A(g4194) );
  INV_X1 NOT_1517( .ZN(g5538), .A(g5331) );
  INV_X1 NOT_1518( .ZN(I6296), .A(g4436) );
  INV_X1 NOT_1519( .ZN(I4646), .A(g2602) );
  INV_X1 NOT_1520( .ZN(I2623), .A(g1161) );
  INV_X1 NOT_1521( .ZN(g4126), .A(I5460) );
  INV_X1 NOT_1522( .ZN(g5509), .A(I7251) );
  INV_X1 NOT_1523( .ZN(g4400), .A(I5899) );
  INV_X2 NOT_1524( .ZN(g1937), .A(I3044) );
  INV_X2 NOT_1525( .ZN(g6541), .A(I8535) );
  INV_X2 NOT_1526( .ZN(I9185), .A(g6877) );
  INV_X2 NOT_1527( .ZN(I2476), .A(g971) );
  INV_X1 NOT_1528( .ZN(I7336), .A(g5534) );
  INV_X1 NOT_1529( .ZN(I8600), .A(g6451) );
  INV_X1 NOT_1530( .ZN(g2931), .A(g1988) );
  INV_X1 NOT_1531( .ZN(g4760), .A(I6386) );
  INV_X1 NOT_1532( .ZN(g1294), .A(I2287) );
  INV_X1 NOT_1533( .ZN(I1877), .A(g283) );
  INV_X1 NOT_1534( .ZN(g6332), .A(I8074) );
  INV_X1 NOT_1535( .ZN(g5067), .A(g4801) );
  INV_X1 NOT_1536( .ZN(g1190), .A(I2199) );
  INV_X1 NOT_1537( .ZN(I2175), .A(g25) );
  INV_X1 NOT_1538( .ZN(g6353), .A(I8113) );
  INV_X1 NOT_1539( .ZN(g5994), .A(g5873) );
  INV_X1 NOT_1540( .ZN(I3608), .A(g1461) );
  INV_X1 NOT_1541( .ZN(g2905), .A(g1994) );
  INV_X1 NOT_1542( .ZN(I6012), .A(g4167) );
  INV_X1 NOT_1543( .ZN(g6744), .A(I8910) );
  INV_X1 NOT_1544( .ZN(I3779), .A(g2125) );
  INV_X1 NOT_1545( .ZN(g6802), .A(I8972) );
  INV_X1 NOT_1546( .ZN(g2628), .A(I3770) );
  INV_X1 NOT_1547( .ZN(g1156), .A(I2175) );
  INV_X1 NOT_1548( .ZN(g2515), .A(I3641) );
  INV_X1 NOT_1549( .ZN(g5493), .A(I7197) );
  INV_X1 NOT_1550( .ZN(I7065), .A(g5281) );
  INV_X1 NOT_1551( .ZN(g5256), .A(g5077) );
  INV_X1 NOT_1552( .ZN(I6706), .A(g4731) );
  INV_X1 NOT_1553( .ZN(g4220), .A(I5644) );
  INV_X1 NOT_1554( .ZN(g3940), .A(I5177) );
  INV_X1 NOT_1555( .ZN(I6371), .A(g4569) );
  INV_X1 NOT_1556( .ZN(I4276), .A(g2170) );
  INV_X1 NOT_1557( .ZN(g4423), .A(I5920) );
  INV_X1 NOT_1558( .ZN(I3161), .A(g1270) );
  INV_X1 NOT_1559( .ZN(I3361), .A(g1331) );
  INV_X1 NOT_1560( .ZN(g5381), .A(I7039) );
  INV_X1 NOT_1561( .ZN(g3388), .A(I4667) );
  INV_X1 NOT_1562( .ZN(I9131), .A(g6855) );
  INV_X1 NOT_1563( .ZN(I6956), .A(g5124) );
  INV_X1 NOT_1564( .ZN(g6901), .A(I9170) );
  INV_X1 NOT_1565( .ZN(I5460), .A(g3771) );
  INV_X1 NOT_1566( .ZN(I5597), .A(g3821) );
  INV_X1 NOT_1567( .ZN(I8623), .A(g6542) );
  INV_X1 NOT_1568( .ZN(g3216), .A(I4459) );
  INV_X1 NOT_1569( .ZN(I3665), .A(g1824) );
  INV_X1 NOT_1570( .ZN(g5685), .A(g5552) );
  INV_X1 NOT_1571( .ZN(g6511), .A(I8453) );
  INV_X1 NOT_1572( .ZN(I8476), .A(g6457) );
  INV_X2 NOT_1573( .ZN(I2424), .A(g719) );
  INV_X2 NOT_1574( .ZN(g743), .A(I1844) );
  INV_X2 NOT_1575( .ZN(g862), .A(g319) );
  INV_X2 NOT_1576( .ZN(g2973), .A(I4170) );
  INV_X1 NOT_1577( .ZN(g1954), .A(I3065) );
  INV_X1 NOT_1578( .ZN(g3030), .A(I4243) );
  INV_X1 NOT_1579( .ZN(g1250), .A(g123) );
  INV_X1 NOT_1580( .ZN(I5739), .A(g3942) );
  INV_X1 NOT_1581( .ZN(g1363), .A(I2399) );
  INV_X1 NOT_1582( .ZN(I4986), .A(g3638) );
  INV_X1 NOT_1583( .ZN(I3999), .A(g1837) );
  INV_X1 NOT_1584( .ZN(g3247), .A(g2973) );
  INV_X1 NOT_1585( .ZN(g4127), .A(I5463) );
  INV_X1 NOT_1586( .ZN(I3346), .A(g1327) );
  INV_X1 NOT_1587( .ZN(g5950), .A(g5730) );
  INV_X1 NOT_1588( .ZN(g1053), .A(g197) );
  INV_X1 NOT_1589( .ZN(g2040), .A(g1738) );
  INV_X1 NOT_1590( .ZN(g6600), .A(I8668) );
  INV_X1 NOT_1591( .ZN(g6574), .A(g6484) );
  INV_X1 NOT_1592( .ZN(I2231), .A(g465) );
  INV_X1 NOT_1593( .ZN(I1844), .A(g208) );
  INV_X1 NOT_1594( .ZN(g2440), .A(I3575) );
  INV_X1 NOT_1595( .ZN(g3564), .A(g2618) );
  INV_X1 NOT_1596( .ZN(g6714), .A(g6670) );
  INV_X1 NOT_1597( .ZN(I2643), .A(g965) );
  INV_X1 NOT_1598( .ZN(g4146), .A(I5520) );
  INV_X1 NOT_1599( .ZN(I5668), .A(g3828) );
  INV_X1 NOT_1600( .ZN(g4633), .A(g4284) );
  INV_X1 NOT_1601( .ZN(I8285), .A(g6310) );
  INV_X1 NOT_1602( .ZN(I5840), .A(g3732) );
  INV_X1 NOT_1603( .ZN(I8500), .A(g6431) );
  INV_X1 NOT_1604( .ZN(g791), .A(I1865) );
  INV_X1 NOT_1605( .ZN(g4103), .A(I5391) );
  INV_X1 NOT_1606( .ZN(g6580), .A(g6491) );
  INV_X1 NOT_1607( .ZN(I7859), .A(g6032) );
  INV_X1 NOT_1608( .ZN(g5631), .A(g5536) );
  INV_X1 NOT_1609( .ZN(g3638), .A(g3108) );
  INV_X1 NOT_1610( .ZN(g5723), .A(I7484) );
  INV_X1 NOT_1611( .ZN(I9173), .A(g6876) );
  INV_X1 NOT_1612( .ZN(I3240), .A(g1460) );
  INV_X1 NOT_1613( .ZN(g4732), .A(I6362) );
  INV_X1 NOT_1614( .ZN(g3108), .A(I4354) );
  INV_X1 NOT_1615( .ZN(g3308), .A(g3060) );
  INV_X1 NOT_1616( .ZN(I6759), .A(g4778) );
  INV_X1 NOT_1617( .ZN(g2875), .A(g1940) );
  INV_X1 NOT_1618( .ZN(g4753), .A(I6377) );
  INV_X1 NOT_1619( .ZN(g4508), .A(I6036) );
  INV_X1 NOT_1620( .ZN(g917), .A(I1942) );
  INV_X1 NOT_1621( .ZN(I8809), .A(g6687) );
  INV_X1 NOT_1622( .ZN(I7342), .A(g5579) );
  INV_X1 NOT_1623( .ZN(g6623), .A(I8727) );
  INV_X1 NOT_1624( .ZN(g6076), .A(g5797) );
  INV_X1 NOT_1625( .ZN(I7081), .A(g5281) );
  INV_X1 NOT_1626( .ZN(g6889), .A(I9134) );
  INV_X1 NOT_1627( .ZN(g5751), .A(I7506) );
  INV_X1 NOT_1628( .ZN(I3316), .A(g1344) );
  INV_X1 NOT_1629( .ZN(g3589), .A(g3094) );
  INV_X1 NOT_1630( .ZN(I7481), .A(g5629) );
  INV_X1 NOT_1631( .ZN(I3034), .A(g1519) );
  INV_X1 NOT_1632( .ZN(g3466), .A(I4706) );
  INV_X1 NOT_1633( .ZN(g2410), .A(I3550) );
  INV_X1 NOT_1634( .ZN(I7692), .A(g5711) );
  INV_X1 NOT_1635( .ZN(I3434), .A(g1627) );
  INV_X1 NOT_1636( .ZN(I4516), .A(g2777) );
  INV_X1 NOT_1637( .ZN(I7497), .A(g5687) );
  INV_X1 NOT_1638( .ZN(g4116), .A(I5430) );
  INV_X1 NOT_1639( .ZN(g6375), .A(I8189) );
  INV_X1 NOT_1640( .ZN(g2884), .A(g1957) );
  INV_X1 NOT_1641( .ZN(I2044), .A(g681) );
  INV_X8 NOT_1642( .ZN(g3571), .A(g3084) );
  INV_X8 NOT_1643( .ZN(g2839), .A(g2535) );
  INV_X1 NOT_1644( .ZN(g3861), .A(I5084) );
  INV_X1 NOT_1645( .ZN(g6722), .A(I8860) );
  INV_X1 NOT_1646( .ZN(g4034), .A(I5333) );
  INV_X1 NOT_1647( .ZN(I7960), .A(g5925) );
  INV_X1 NOT_1648( .ZN(g852), .A(g634) );
  INV_X1 NOT_1649( .ZN(I2269), .A(g899) );
  INV_X1 NOT_1650( .ZN(g6651), .A(I8749) );
  INV_X1 NOT_1651( .ZN(g3448), .A(I4684) );
  INV_X1 NOT_1652( .ZN(g4565), .A(g4195) );
  INV_X1 NOT_1653( .ZN(I3681), .A(g1821) );
  INV_X1 NOT_1654( .ZN(I5053), .A(g3710) );
  INV_X1 NOT_1655( .ZN(g3455), .A(g2637) );
  INV_X1 NOT_1656( .ZN(g6285), .A(I8005) );
  INV_X1 NOT_1657( .ZN(g4147), .A(I5523) );
  INV_X1 NOT_1658( .ZN(g6500), .A(I8420) );
  INV_X1 NOT_1659( .ZN(g2172), .A(I3307) );
  INV_X1 NOT_1660( .ZN(I2712), .A(g1203) );
  INV_X1 NOT_1661( .ZN(I9227), .A(g6937) );
  INV_X1 NOT_1662( .ZN(I5568), .A(g3897) );
  INV_X1 NOT_1663( .ZN(g4533), .A(I6111) );
  INV_X1 NOT_1664( .ZN(g3846), .A(I5053) );
  INV_X1 NOT_1665( .ZN(g2618), .A(I3758) );
  INV_X1 NOT_1666( .ZN(I3596), .A(g1305) );
  INV_X1 NOT_1667( .ZN(g2667), .A(I3811) );
  INV_X1 NOT_1668( .ZN(g1683), .A(g1017) );
  INV_X1 NOT_1669( .ZN(g2343), .A(I3493) );
  INV_X1 NOT_1670( .ZN(g5168), .A(g5099) );
  INV_X1 NOT_1671( .ZN(I3013), .A(g1519) );
  INV_X1 NOT_1672( .ZN(g6339), .A(I8093) );
  INV_X1 NOT_1673( .ZN(g3196), .A(I4433) );
  INV_X1 NOT_1674( .ZN(g4914), .A(g4816) );
  INV_X1 NOT_1675( .ZN(g3803), .A(I5002) );
  INV_X1 NOT_1676( .ZN(g4210), .A(I5630) );
  INV_X1 NOT_1677( .ZN(I7267), .A(g5458) );
  INV_X1 NOT_1678( .ZN(g1894), .A(I2989) );
  INV_X1 NOT_1679( .ZN(I5157), .A(g3454) );
  INV_X1 NOT_1680( .ZN(g6838), .A(I9035) );
  INV_X1 NOT_1681( .ZN(I9203), .A(g6921) );
  INV_X1 NOT_1682( .ZN(I2961), .A(g1731) );
  INV_X1 NOT_1683( .ZN(g6424), .A(I8282) );
  INV_X1 NOT_1684( .ZN(g2134), .A(I3258) );
  INV_X1 NOT_1685( .ZN(I6362), .A(g4569) );
  INV_X1 NOT_1686( .ZN(g1735), .A(I2745) );
  INV_X1 NOT_1687( .ZN(I8273), .A(g6301) );
  INV_X1 NOT_1688( .ZN(g6809), .A(I8981) );
  INV_X1 NOT_1689( .ZN(g5890), .A(g5753) );
  INV_X1 NOT_1690( .ZN(g1782), .A(I2828) );
  INV_X1 NOT_1691( .ZN(I4340), .A(g1935) );
  INV_X1 NOT_1692( .ZN(I6452), .A(g4629) );
  INV_X1 NOT_1693( .ZN(I5929), .A(g4152) );
  INV_X1 NOT_1694( .ZN(g1661), .A(g1076) );
  INV_X1 NOT_1695( .ZN(I8044), .A(g6252) );
  INV_X1 NOT_1696( .ZN(g2555), .A(I3672) );
  INV_X1 NOT_1697( .ZN(g6231), .A(g6044) );
  INV_X8 NOT_1698( .ZN(g5011), .A(I6649) );
  INV_X8 NOT_1699( .ZN(I8444), .A(g6421) );
  INV_X1 NOT_1700( .ZN(g3067), .A(I4294) );
  INV_X1 NOT_1701( .ZN(I2414), .A(g784) );
  INV_X1 NOT_1702( .ZN(g729), .A(I1838) );
  INV_X1 NOT_1703( .ZN(g5411), .A(I7077) );
  INV_X1 NOT_1704( .ZN(g6523), .A(I8485) );
  INV_X1 NOT_1705( .ZN(g861), .A(g179) );
  INV_X1 NOT_1706( .ZN(I2946), .A(g1587) );
  INV_X1 NOT_1707( .ZN(g2792), .A(g2416) );
  INV_X1 NOT_1708( .ZN(g1627), .A(I2584) );
  INV_X1 NOT_1709( .ZN(g4117), .A(I5433) );
  INV_X1 NOT_1710( .ZN(g1292), .A(I2281) );
  INV_X1 NOT_1711( .ZN(I5626), .A(g3914) );
  INV_X1 NOT_1712( .ZN(g3093), .A(I4334) );
  INV_X1 NOT_1713( .ZN(g898), .A(g47) );
  INV_X1 NOT_1714( .ZN(g1998), .A(I3109) );
  INV_X1 NOT_1715( .ZN(g1646), .A(I2617) );
  INV_X1 NOT_1716( .ZN(g5992), .A(g5869) );
  INV_X1 NOT_1717( .ZN(g4601), .A(g4191) );
  INV_X1 NOT_1718( .ZN(g1084), .A(g98) );
  INV_X1 NOT_1719( .ZN(g6104), .A(I7808) );
  INV_X1 NOT_1720( .ZN(g854), .A(g646) );
  INV_X1 NOT_1721( .ZN(g1039), .A(g662) );
  INV_X1 NOT_1722( .ZN(g1484), .A(I2473) );
  INV_X1 NOT_1723( .ZN(I3581), .A(g1491) );
  INV_X1 NOT_1724( .ZN(g6499), .A(I8417) );
  INV_X1 NOT_1725( .ZN(g1439), .A(I2449) );
  INV_X1 NOT_1726( .ZN(I9028), .A(g6806) );
  INV_X1 NOT_1727( .ZN(I8961), .A(g6778) );
  INV_X1 NOT_1728( .ZN(g4775), .A(I6425) );
  INV_X1 NOT_1729( .ZN(I6470), .A(g4473) );
  INV_X1 NOT_1730( .ZN(g5573), .A(g5403) );
  INV_X1 NOT_1731( .ZN(g3847), .A(I5056) );
  INV_X1 NOT_1732( .ZN(g5480), .A(I7176) );
  INV_X1 NOT_1733( .ZN(I6425), .A(g4619) );
  INV_X1 NOT_1734( .ZN(I2831), .A(g1209) );
  INV_X1 NOT_1735( .ZN(g2494), .A(I3623) );
  INV_X1 NOT_1736( .ZN(I2182), .A(g692) );
  INV_X1 NOT_1737( .ZN(g2518), .A(I3644) );
  INV_X1 NOT_1738( .ZN(g1583), .A(g1001) );
  INV_X1 NOT_1739( .ZN(g1702), .A(g1107) );
  INV_X1 NOT_1740( .ZN(I2382), .A(g719) );
  INV_X1 NOT_1741( .ZN(I8414), .A(g6418) );
  INV_X1 NOT_1742( .ZN(g3263), .A(g3015) );
  INV_X1 NOT_1743( .ZN(I8946), .A(g6778) );
  INV_X1 NOT_1744( .ZN(g1919), .A(I3022) );
  INV_X1 NOT_1745( .ZN(I2805), .A(g1205) );
  INV_X1 NOT_1746( .ZN(I2916), .A(g1643) );
  INV_X1 NOT_1747( .ZN(g2776), .A(g2378) );
  INV_X1 NOT_1748( .ZN(I2749), .A(g1209) );
  INV_X1 NOT_1749( .ZN(g4784), .A(I6444) );
  INV_X1 NOT_1750( .ZN(g6044), .A(g5824) );
  INV_X1 NOT_1751( .ZN(g1276), .A(g847) );
  INV_X1 NOT_1752( .ZN(I4402), .A(g2283) );
  INV_X1 NOT_1753( .ZN(I3294), .A(g1720) );
  INV_X1 NOT_1754( .ZN(I3840), .A(g2125) );
  INV_X1 NOT_1755( .ZN(I6406), .A(g4473) );
  INV_X1 NOT_1756( .ZN(I5475), .A(g3852) );
  INV_X1 NOT_1757( .ZN(g6572), .A(I8600) );
  INV_X1 NOT_1758( .ZN(I4762), .A(g2862) );
  INV_X1 NOT_1759( .ZN(I7349), .A(g5532) );
  INV_X1 NOT_1760( .ZN(I6635), .A(g4745) );
  INV_X1 NOT_1761( .ZN(g2264), .A(I3405) );
  INV_X1 NOT_1762( .ZN(g6712), .A(g6676) );
  INV_X1 NOT_1763( .ZN(g851), .A(g606) );
  INV_X1 NOT_1764( .ZN(I6766), .A(g4783) );
  INV_X1 NOT_1765( .ZN(I6087), .A(g4392) );
  INV_X1 NOT_1766( .ZN(I6105), .A(g4400) );
  INV_X1 NOT_1767( .ZN(g6543), .A(I8541) );
  INV_X1 NOT_1768( .ZN(g4840), .A(I6528) );
  INV_X1 NOT_1769( .ZN(I6305), .A(g4441) );
  INV_X1 NOT_1770( .ZN(I6801), .A(g5045) );
  INV_X1 NOT_1771( .ZN(g2360), .A(g1793) );
  INV_X1 NOT_1772( .ZN(g2933), .A(I4123) );
  INV_X1 NOT_1773( .ZN(g3723), .A(I4903) );
  INV_X1 NOT_1774( .ZN(g1647), .A(I2620) );
  INV_X1 NOT_1775( .ZN(g4190), .A(I5600) );
  INV_X1 NOT_1776( .ZN(I5526), .A(g3848) );
  INV_X1 NOT_1777( .ZN(I5998), .A(g4157) );
  INV_X1 NOT_1778( .ZN(I8335), .A(g6308) );
  INV_X1 NOT_1779( .ZN(I8831), .A(g6665) );
  INV_X1 NOT_1780( .ZN(I9217), .A(g6931) );
  INV_X1 NOT_1781( .ZN(g1546), .A(g1101) );
  INV_X1 NOT_1782( .ZN(I2873), .A(g1161) );
  INV_X1 NOT_1783( .ZN(I2037), .A(g679) );
  INV_X1 NOT_1784( .ZN(g6534), .A(I8518) );
  INV_X1 NOT_1785( .ZN(g6729), .A(I8881) );
  INV_X8 NOT_1786( .ZN(g3605), .A(I4802) );
  INV_X8 NOT_1787( .ZN(I5084), .A(g3593) );
  INV_X8 NOT_1788( .ZN(I5603), .A(g3893) );
  INV_X1 NOT_1789( .ZN(g2996), .A(I4189) );
  INV_X1 NOT_1790( .ZN(I2653), .A(g996) );
  INV_X1 NOT_1791( .ZN(I5484), .A(g3875) );
  INV_X1 NOT_1792( .ZN(I3942), .A(g1833) );
  INV_X1 NOT_1793( .ZN(g1503), .A(g878) );
  INV_X1 NOT_1794( .ZN(I5439), .A(g3730) );
  INV_X1 NOT_1795( .ZN(I8916), .A(g6742) );
  INV_X1 NOT_1796( .ZN(g1925), .A(I3028) );
  INV_X1 NOT_1797( .ZN(I8749), .A(g6560) );
  INV_X1 NOT_1798( .ZN(g2179), .A(I3328) );
  INV_X1 NOT_1799( .ZN(g6014), .A(g5824) );
  INV_X1 NOT_1800( .ZN(g6885), .A(I9122) );
  INV_X1 NOT_1801( .ZN(I6045), .A(g4375) );
  INV_X1 NOT_1802( .ZN(g4704), .A(I6302) );
  INV_X1 NOT_1803( .ZN(g6414), .A(I8252) );
  INV_X1 NOT_1804( .ZN(I5702), .A(g3845) );
  INV_X1 NOT_1805( .ZN(g1320), .A(I2315) );
  INV_X1 NOT_1806( .ZN(g3041), .A(I4258) );
  INV_X1 NOT_1807( .ZN(g5383), .A(I7045) );
  INV_X1 NOT_1808( .ZN(g5924), .A(I7704) );
  INV_X1 NOT_1809( .ZN(g5220), .A(g4903) );
  INV_X1 NOT_1810( .ZN(I7119), .A(g5303) );
  INV_X1 NOT_1811( .ZN(g6903), .A(I9176) );
  INV_X1 NOT_1812( .ZN(g2777), .A(I3965) );
  INV_X1 NOT_1813( .ZN(g3441), .A(I4681) );
  INV_X1 NOT_1814( .ZN(g2835), .A(g2506) );
  INV_X1 NOT_1815( .ZN(I3053), .A(g1407) );
  INV_X1 NOT_1816( .ZN(I1958), .A(g702) );
  INV_X1 NOT_1817( .ZN(g4250), .A(I5702) );
  INV_X1 NOT_1818( .ZN(g6513), .A(I8459) );
  INV_X1 NOT_1819( .ZN(g913), .A(g658) );
  INV_X1 NOT_1820( .ZN(I6283), .A(g4613) );
  INV_X1 NOT_1821( .ZN(I7258), .A(g5458) );
  INV_X1 NOT_1822( .ZN(I5952), .A(g4367) );
  INV_X1 NOT_1823( .ZN(g4810), .A(I6488) );
  INV_X1 NOT_1824( .ZN(g2882), .A(g1854) );
  INV_X1 NOT_1825( .ZN(I7352), .A(g5533) );
  INV_X1 NOT_1826( .ZN(g3673), .A(g3075) );
  INV_X1 NOT_1827( .ZN(I2442), .A(g872) );
  INV_X1 NOT_1828( .ZN(g1789), .A(I2839) );
  INV_X1 NOT_1829( .ZN(g6036), .A(g5824) );
  INV_X1 NOT_1830( .ZN(I8632), .A(g6548) );
  INV_X1 NOT_1831( .ZN(I2364), .A(g1143) );
  INV_X1 NOT_1832( .ZN(g980), .A(I2037) );
  INV_X1 NOT_1833( .ZN(I8653), .A(g6531) );
  INV_X1 NOT_1834( .ZN(g1771), .A(I2808) );
  INV_X1 NOT_1835( .ZN(g3772), .A(g3466) );
  INV_X1 NOT_1836( .ZN(I6582), .A(g4765) );
  INV_X1 NOT_1837( .ZN(g5051), .A(I6689) );
  INV_X1 NOT_1838( .ZN(g2981), .A(g2179) );
  INV_X1 NOT_1839( .ZN(I8579), .A(g6438) );
  INV_X1 NOT_1840( .ZN(I8869), .A(g6694) );
  INV_X1 NOT_1841( .ZN(I4489), .A(g2975) );
  INV_X1 NOT_1842( .ZN(g3458), .A(g2656) );
  INV_X1 NOT_1843( .ZN(g865), .A(g188) );
  INV_X1 NOT_1844( .ZN(I2296), .A(g893) );
  INV_X1 NOT_1845( .ZN(g3890), .A(g3575) );
  INV_X1 NOT_1846( .ZN(g2997), .A(I4192) );
  INV_X1 NOT_1847( .ZN(I6015), .A(g4170) );
  INV_X2 NOT_1848( .ZN(g2541), .A(I3659) );
  INV_X2 NOT_1849( .ZN(I8752), .A(g6514) );
  INV_X2 NOT_1850( .ZN(I4471), .A(g3040) );
  INV_X1 NOT_1851( .ZN(I7170), .A(g5435) );
  INV_X1 NOT_1852( .ZN(g6422), .A(I8276) );
  INV_X1 NOT_1853( .ZN(g2353), .A(I3505) );
  INV_X1 NOT_1854( .ZN(g4929), .A(I6621) );
  INV_X1 NOT_1855( .ZN(I4955), .A(g3673) );
  INV_X1 NOT_1856( .ZN(I3626), .A(g1684) );
  INV_X1 NOT_1857( .ZN(g2744), .A(g2336) );
  INV_X1 NOT_1858( .ZN(g909), .A(I1935) );
  INV_X1 NOT_1859( .ZN(g1738), .A(g1108) );
  INV_X1 NOT_1860( .ZN(g2802), .A(g2437) );
  INV_X1 NOT_1861( .ZN(g3074), .A(I4303) );
  INV_X1 NOT_1862( .ZN(g949), .A(g79) );
  INV_X1 NOT_1863( .ZN(g1991), .A(I3102) );
  INV_X1 NOT_1864( .ZN(g6560), .A(I8564) );
  INV_X1 NOT_1865( .ZN(I5320), .A(g3559) );
  INV_X1 NOT_1866( .ZN(g4626), .A(g4270) );
  INV_X1 NOT_1867( .ZN(g1340), .A(I2373) );
  INV_X1 NOT_1868( .ZN(I2029), .A(g677) );
  INV_X1 NOT_1869( .ZN(I9021), .A(g6812) );
  INV_X1 NOT_1870( .ZN(g3480), .A(g2986) );
  INV_X1 NOT_1871( .ZN(g1690), .A(I2692) );
  INV_X1 NOT_1872( .ZN(g6653), .A(I8755) );
  INV_X1 NOT_1873( .ZN(g6102), .A(I7802) );
  INV_X1 NOT_1874( .ZN(I2281), .A(g900) );
  INV_X1 NOT_1875( .ZN(I7061), .A(g5281) );
  INV_X1 NOT_1876( .ZN(I7187), .A(g5387) );
  INV_X1 NOT_1877( .ZN(g6579), .A(g6490) );
  INV_X1 NOT_1878( .ZN(g5116), .A(g4810) );
  INV_X1 NOT_1879( .ZN(I5987), .A(g4224) );
  INV_X1 NOT_1880( .ZN(g5316), .A(I6976) );
  INV_X1 NOT_1881( .ZN(g1656), .A(I2635) );
  INV_X1 NOT_1882( .ZN(I6689), .A(g4758) );
  INV_X1 NOT_1883( .ZN(g5434), .A(I7110) );
  INV_X1 NOT_1884( .ZN(g2574), .A(I3681) );
  INV_X1 NOT_1885( .ZN(g2864), .A(g1887) );
  INV_X1 NOT_1886( .ZN(g4778), .A(I6430) );
  INV_X1 NOT_1887( .ZN(g855), .A(g650) );
  INV_X1 NOT_1888( .ZN(g5147), .A(I6809) );
  INV_X1 NOT_1889( .ZN(I3782), .A(g2145) );
  INV_X1 NOT_1890( .ZN(g4894), .A(g4813) );
  INV_X1 NOT_1891( .ZN(I2745), .A(g1249) );
  INV_X1 NOT_1892( .ZN(I8189), .A(g6179) );
  INV_X1 NOT_1893( .ZN(I4229), .A(g2284) );
  INV_X1 NOT_1894( .ZN(I6430), .A(g4620) );
  INV_X1 NOT_1895( .ZN(g3976), .A(I5252) );
  INV_X1 NOT_1896( .ZN(I2791), .A(g1236) );
  INV_X1 NOT_1897( .ZN(I6247), .A(g4609) );
  INV_X1 NOT_1898( .ZN(I7514), .A(g5590) );
  INV_X1 NOT_1899( .ZN(I2309), .A(g1236) );
  INV_X1 NOT_1900( .ZN(I9101), .A(g6855) );
  INV_X1 NOT_1901( .ZN(g1110), .A(I2140) );
  INV_X1 NOT_1902( .ZN(I8888), .A(g6708) );
  INV_X1 NOT_1903( .ZN(g2580), .A(I3691) );
  INV_X1 NOT_1904( .ZN(g5210), .A(I6874) );
  INV_X1 NOT_1905( .ZN(g6786), .A(I8946) );
  INV_X1 NOT_1906( .ZN(I6564), .A(g4712) );
  INV_X1 NOT_1907( .ZN(I8171), .A(g6170) );
  INV_X1 NOT_1908( .ZN(I2808), .A(g1161) );
  INV_X1 NOT_1909( .ZN(I8429), .A(g6425) );
  INV_X1 NOT_1910( .ZN(g5596), .A(I7358) );
  INV_X1 NOT_1911( .ZN(g6164), .A(g5926) );
  INV_X2 NOT_1912( .ZN(g6364), .A(I8156) );
  INV_X2 NOT_1913( .ZN(g6233), .A(g6052) );
  INV_X2 NOT_1914( .ZN(I5991), .A(g4226) );
  INV_X2 NOT_1915( .ZN(I2707), .A(g1190) );
  INV_X2 NOT_1916( .ZN(g4292), .A(g4059) );
  INV_X4 NOT_1917( .ZN(I7695), .A(g5714) );
  INV_X4 NOT_1918( .ZN(I7637), .A(g5751) );
  INV_X4 NOT_1919( .ZN(g2968), .A(g2179) );
  INV_X2 NOT_1920( .ZN(I5078), .A(g3719) );
  INV_X4 NOT_1921( .ZN(g1824), .A(I2890) );
  INV_X4 NOT_1922( .ZN(g4526), .A(I6090) );
  INV_X4 NOT_1923( .ZN(I5478), .A(g3859) );
  INV_X1 NOT_1924( .ZN(g1236), .A(I2234) );
  INV_X1 NOT_1925( .ZN(I7107), .A(g5277) );
  INV_X1 NOT_1926( .ZN(I5907), .A(g3883) );
  INV_X1 NOT_1927( .ZN(g6725), .A(I8869) );
  INV_X1 NOT_1928( .ZN(g1762), .A(I2791) );
  INV_X1 NOT_1929( .ZN(g2889), .A(g1975) );
  INV_X1 NOT_1930( .ZN(I6108), .A(g4403) );
  INV_X1 NOT_1931( .ZN(g4603), .A(I6170) );
  INV_X1 NOT_1932( .ZN(g6532), .A(I8512) );
  INV_X2 NOT_1933( .ZN(I6308), .A(g4443) );
  INV_X1 NOT_1934( .ZN(I5517), .A(g3885) );
  INV_X1 NOT_1935( .ZN(I9041), .A(g6835) );
  INV_X1 NOT_1936( .ZN(I2449), .A(g971) );
  INV_X1 NOT_1937( .ZN(g4439), .A(I5952) );
  INV_X1 NOT_1938( .ZN(g5117), .A(I6763) );
  INV_X1 NOT_1939( .ZN(g6553), .A(I8555) );
  INV_X1 NOT_1940( .ZN(g4850), .A(I6558) );
  INV_X1 NOT_1941( .ZN(I8684), .A(g6567) );
  INV_X1 NOT_1942( .ZN(I5876), .A(g3870) );
  INV_X1 NOT_1943( .ZN(I8745), .A(g6513) );
  INV_X1 NOT_1944( .ZN(g2175), .A(I3316) );
  INV_X1 NOT_1945( .ZN(g2871), .A(g1919) );
  INV_X2 NOT_1946( .ZN(I2604), .A(g1222) );
  INV_X1 NOT_1947( .ZN(g3183), .A(I4420) );
  INV_X1 NOT_1948( .ZN(g2722), .A(I3883) );
  INV_X1 NOT_1949( .ZN(I4462), .A(g2135) );
  INV_X1 NOT_1950( .ZN(I8309), .A(g6304) );
  INV_X1 NOT_1951( .ZN(g1556), .A(g878) );
  INV_X1 NOT_1952( .ZN(I6066), .A(g4382) );
  INV_X1 NOT_1953( .ZN(g3779), .A(g3466) );
  INV_X1 NOT_1954( .ZN(g1222), .A(I2225) );
  INV_X1 NOT_1955( .ZN(g4702), .A(I6296) );
  INV_X1 NOT_1956( .ZN(g6412), .A(I8246) );
  INV_X1 NOT_1957( .ZN(g896), .A(g22) );
  INV_X1 NOT_1958( .ZN(g3023), .A(g2215) );
  INV_X1 NOT_1959( .ZN(I7251), .A(g5458) );
  INV_X1 NOT_1960( .ZN(g1928), .A(I3031) );
  INV_X1 NOT_1961( .ZN(I7811), .A(g5921) );
  INV_X1 NOT_1962( .ZN(g6706), .A(I8828) );
  INV_X1 NOT_1963( .ZN(g5922), .A(I7698) );
  INV_X1 NOT_1964( .ZN(I8707), .A(g6520) );
  INV_X1 NOT_1965( .ZN(g1064), .A(g102) );
  INV_X1 NOT_1966( .ZN(I2584), .A(g839) );
  INV_X1 NOT_1967( .ZN(I5214), .A(g3567) );
  INV_X1 NOT_1968( .ZN(g6888), .A(I9131) );
  INV_X1 NOT_1969( .ZN(g1899), .A(I2998) );
  INV_X1 NOT_1970( .ZN(I6048), .A(g4376) );
  INV_X1 NOT_1971( .ZN(g5581), .A(I7339) );
  INV_X1 NOT_1972( .ZN(I6448), .A(g4626) );
  INV_X1 NOT_1973( .ZN(g6371), .A(I8177) );
  INV_X1 NOT_1974( .ZN(g4276), .A(I5731) );
  INV_X1 NOT_1975( .ZN(I4249), .A(g2525) );
  INV_X1 NOT_1976( .ZN(g5597), .A(I7361) );
  INV_X1 NOT_1977( .ZN(I3004), .A(g1426) );
  INV_X1 NOT_1978( .ZN(I1825), .A(g361) );
  INV_X1 NOT_1979( .ZN(g4561), .A(g4189) );
  INV_X1 NOT_1980( .ZN(g2838), .A(g2515) );
  INV_X1 NOT_1981( .ZN(I3647), .A(g1747) );
  INV_X1 NOT_1982( .ZN(g3451), .A(g2615) );
  INV_X1 NOT_1983( .ZN(I2162), .A(g197) );
  INV_X1 NOT_1984( .ZN(g1563), .A(g1006) );
  INV_X1 NOT_1985( .ZN(I9011), .A(g6819) );
  INV_X1 NOT_1986( .ZN(I4192), .A(g1847) );
  INV_X1 NOT_1987( .ZN(g2809), .A(I4019) );
  INV_X1 NOT_1988( .ZN(I3764), .A(g2044) );
  INV_X1 NOT_1989( .ZN(g5784), .A(I7583) );
  INV_X1 NOT_1990( .ZN(I3546), .A(g1586) );
  INV_X1 NOT_1991( .ZN(I5002), .A(g3612) );
  INV_X1 NOT_1992( .ZN(g4527), .A(I6093) );
  INV_X1 NOT_1993( .ZN(g4404), .A(I5907) );
  INV_X1 NOT_1994( .ZN(g1295), .A(I2290) );
  INV_X1 NOT_1995( .ZN(g4647), .A(g4296) );
  INV_X1 NOT_1996( .ZN(g3346), .A(I4623) );
  INV_X1 NOT_1997( .ZN(I5236), .A(g3545) );
  INV_X1 NOT_1998( .ZN(g2672), .A(I3816) );
  INV_X1 NOT_1999( .ZN(g2231), .A(I3358) );
  INV_X1 NOT_2000( .ZN(g4764), .A(I6400) );
  INV_X1 NOT_2001( .ZN(g5995), .A(g5824) );
  INV_X1 NOT_2002( .ZN(I9074), .A(g6844) );
  INV_X1 NOT_2003( .ZN(g5479), .A(I7173) );
  INV_X1 NOT_2004( .ZN(g2643), .A(I3785) );
  INV_X1 NOT_2005( .ZN(I6780), .A(g4825) );
  INV_X1 NOT_2006( .ZN(g6745), .A(I8913) );
  INV_X1 NOT_2007( .ZN(g1394), .A(g1206) );
  INV_X1 NOT_2008( .ZN(g4503), .A(I6023) );
  INV_X1 NOT_2009( .ZN(I7612), .A(g5605) );
  INV_X1 NOT_2010( .ZN(g1731), .A(I2735) );
  INV_X1 NOT_2011( .ZN(I2728), .A(g1232) );
  INV_X1 NOT_2012( .ZN(g1557), .A(g1017) );
  INV_X1 NOT_2013( .ZN(g2634), .A(I3776) );
  INV_X1 NOT_2014( .ZN(g1966), .A(I3077) );
  INV_X1 NOT_2015( .ZN(g4224), .A(g4046) );
  INV_X1 NOT_2016( .ZN(I5556), .A(g4059) );
  INV_X1 NOT_2017( .ZN(I2185), .A(g29) );
  INV_X1 NOT_2018( .ZN(g2104), .A(g1372) );
  INV_X1 NOT_2019( .ZN(g2099), .A(g1366) );
  INV_X1 NOT_2020( .ZN(g3240), .A(I4519) );
  INV_X1 NOT_2021( .ZN(I2385), .A(g784) );
  INV_X1 NOT_2022( .ZN(g6707), .A(I8831) );
  INV_X1 NOT_2023( .ZN(g1471), .A(I2464) );
  INV_X1 NOT_2024( .ZN(g4120), .A(I5442) );
  INV_X1 NOT_2025( .ZN(I4031), .A(g1846) );
  INV_X1 NOT_2026( .ZN(g4320), .A(g4011) );
  INV_X1 NOT_2027( .ZN(I4252), .A(g2555) );
  INV_X1 NOT_2028( .ZN(I3617), .A(g1305) );
  INV_X1 NOT_2029( .ZN(I3906), .A(g2234) );
  INV_X1 NOT_2030( .ZN(I6093), .A(g4394) );
  INV_X1 NOT_2031( .ZN(I8162), .A(g6189) );
  INV_X1 NOT_2032( .ZN(g3043), .A(I4264) );
  INV_X1 NOT_2033( .ZN(g971), .A(g658) );
  INV_X1 NOT_2034( .ZN(I5899), .A(g3748) );
  INV_X1 NOT_2035( .ZN(I4176), .A(g2268) );
  INV_X1 NOT_2036( .ZN(I6816), .A(g5111) );
  INV_X1 NOT_2037( .ZN(I3516), .A(g1295) );
  INV_X1 NOT_2038( .ZN(g2754), .A(g2347) );
  INV_X1 NOT_2039( .ZN(g4617), .A(g4242) );
  INV_X1 NOT_2040( .ZN(g3034), .A(I4249) );
  INV_X1 NOT_2041( .ZN(g1254), .A(g152) );
  INV_X1 NOT_2042( .ZN(g1814), .A(I2873) );
  INV_X4 NOT_2043( .ZN(g6575), .A(g6486) );
  INV_X4 NOT_2044( .ZN(g4516), .A(I6060) );
  INV_X1 NOT_2045( .ZN(g6715), .A(g6673) );
  INV_X1 NOT_2046( .ZN(g4771), .A(I6417) );
  INV_X1 NOT_2047( .ZN(g2044), .A(I3161) );
  INV_X1 NOT_2048( .ZN(I6685), .A(g4716) );
  INV_X1 NOT_2049( .ZN(g5250), .A(g4929) );
  INV_X1 NOT_2050( .ZN(g6604), .A(I8678) );
  INV_X1 NOT_2051( .ZN(g1038), .A(g127) );
  INV_X1 NOT_2052( .ZN(I6397), .A(g4473) );
  INV_X1 NOT_2053( .ZN(g6498), .A(I8414) );
  INV_X1 NOT_2054( .ZN(g1773), .A(I2814) );
  INV_X1 NOT_2055( .ZN(I2131), .A(g24) );
  INV_X1 NOT_2056( .ZN(g5432), .A(I7104) );
  INV_X1 NOT_2057( .ZN(g4299), .A(I5756) );
  INV_X1 NOT_2058( .ZN(g6833), .A(I9024) );
  INV_X1 NOT_2059( .ZN(I8730), .A(g6535) );
  INV_X1 NOT_2060( .ZN(g5453), .A(g5296) );
  INV_X1 NOT_2061( .ZN(I4270), .A(g2555) );
  INV_X1 NOT_2062( .ZN(g2862), .A(I4066) );
  INV_X1 NOT_2063( .ZN(I2635), .A(g1055) );
  INV_X1 NOT_2064( .ZN(g2712), .A(g2320) );
  INV_X1 NOT_2065( .ZN(I8881), .A(g6711) );
  INV_X1 NOT_2066( .ZN(I5394), .A(g4016) );
  INV_X1 NOT_2067( .ZN(g1769), .A(I2802) );
  INV_X1 NOT_2068( .ZN(g3914), .A(I5153) );
  INV_X1 NOT_2069( .ZN(g6584), .A(I8620) );
  INV_X1 NOT_2070( .ZN(I1859), .A(g277) );
  INV_X1 NOT_2071( .ZN(g6539), .A(I8531) );
  INV_X1 NOT_2072( .ZN(g6896), .A(I9155) );
  INV_X1 NOT_2073( .ZN(g1836), .A(I2922) );
  INV_X1 NOT_2074( .ZN(g5568), .A(g5423) );
  INV_X1 NOT_2075( .ZN(I8070), .A(g6116) );
  INV_X1 NOT_2076( .ZN(I5731), .A(g3942) );
  INV_X1 NOT_2077( .ZN(I8470), .A(g6461) );
  INV_X1 NOT_2078( .ZN(I8897), .A(g6707) );
  INV_X1 NOT_2079( .ZN(g1918), .A(I3019) );
  INV_X1 NOT_2080( .ZN(I3244), .A(g1772) );
  INV_X1 NOT_2081( .ZN(I7490), .A(g5583) );
  INV_X1 NOT_2082( .ZN(I4980), .A(g3546) );
  INV_X1 NOT_2083( .ZN(g5912), .A(g5853) );
  INV_X1 NOT_2084( .ZN(I4324), .A(g1918) );
  INV_X1 NOT_2085( .ZN(I3140), .A(g1317) );
  INV_X1 NOT_2086( .ZN(g2961), .A(g1861) );
  INV_X1 NOT_2087( .ZN(I5071), .A(g3263) );
  INV_X1 NOT_2088( .ZN(I3340), .A(g1282) );
  INV_X1 NOT_2089( .ZN(I5705), .A(g3942) );
  INV_X1 NOT_2090( .ZN(g6162), .A(g5926) );
  INV_X1 NOT_2091( .ZN(I3478), .A(g1450) );
  INV_X1 NOT_2092( .ZN(g6362), .A(I8150) );
  INV_X1 NOT_2093( .ZN(g6419), .A(I8267) );
  INV_X1 NOT_2094( .ZN(I6723), .A(g4761) );
  INV_X1 NOT_2095( .ZN(g4140), .A(I5502) );
  INV_X1 NOT_2096( .ZN(g6052), .A(g5824) );
  INV_X1 NOT_2097( .ZN(g2927), .A(g1979) );
  INV_X1 NOT_2098( .ZN(I5948), .A(g4360) );
  INV_X1 NOT_2099( .ZN(I9220), .A(g6930) );
  INV_X1 NOT_2100( .ZN(g2885), .A(g1963) );
  INV_X1 NOT_2101( .ZN(I7355), .A(g5535) );
  INV_X1 NOT_2102( .ZN(I8678), .A(g6565) );
  INV_X1 NOT_2103( .ZN(I2445), .A(g971) );
  INV_X1 NOT_2104( .ZN(g2660), .A(I3804) );
  INV_X1 NOT_2105( .ZN(g2946), .A(g2296) );
  INV_X2 NOT_2106( .ZN(g938), .A(g59) );
  INV_X2 NOT_2107( .ZN(g4435), .A(I5944) );
  INV_X1 NOT_2108( .ZN(I2373), .A(g1143) );
  INV_X1 NOT_2109( .ZN(g4517), .A(I6063) );
  INV_X1 NOT_2110( .ZN(I7698), .A(g5717) );
  INV_X1 NOT_2111( .ZN(I3656), .A(g1484) );
  INV_X1 NOT_2112( .ZN(g3601), .A(I4794) );
  INV_X1 NOT_2113( .ZN(I2491), .A(g821) );
  INV_X1 NOT_2114( .ZN(g2903), .A(g1902) );
  INV_X1 NOT_2115( .ZN(I8635), .A(g6552) );
  INV_X1 NOT_2116( .ZN(g6728), .A(I8878) );
  INV_X1 NOT_2117( .ZN(g6486), .A(g6363) );
  INV_X1 NOT_2118( .ZN(I2169), .A(g269) );
  INV_X1 NOT_2119( .ZN(g942), .A(g69) );
  INV_X1 NOT_2120( .ZN(g6730), .A(I8884) );
  INV_X1 NOT_2121( .ZN(I9161), .A(g6880) );
  INV_X1 NOT_2122( .ZN(g3775), .A(g3388) );
  INV_X1 NOT_2123( .ZN(g6504), .A(I8432) );
  INV_X1 NOT_2124( .ZN(g3922), .A(I5157) );
  INV_X1 NOT_2125( .ZN(I7463), .A(g5622) );
  INV_X1 NOT_2126( .ZN(I2578), .A(g1209) );
  INV_X1 NOT_2127( .ZN(g6385), .A(g6271) );
  INV_X1 NOT_2128( .ZN(g6881), .A(I9110) );
  INV_X1 NOT_2129( .ZN(I5409), .A(g3980) );
  INV_X1 NOT_2130( .ZN(g2036), .A(g1764) );
  INV_X1 NOT_2131( .ZN(g706), .A(I1825) );
  INV_X1 NOT_2132( .ZN(I6441), .A(g4624) );
  INV_X1 NOT_2133( .ZN(g4915), .A(g4669) );
  INV_X1 NOT_2134( .ZN(g2178), .A(I3325) );
  INV_X1 NOT_2135( .ZN(g2436), .A(I3569) );
  INV_X1 NOT_2136( .ZN(g2679), .A(I3823) );
  INV_X1 NOT_2137( .ZN(g6070), .A(g5824) );
  INV_X1 NOT_2138( .ZN(g2378), .A(I3525) );
  INV_X1 NOT_2139( .ZN(g3060), .A(I4285) );
  INV_X1 NOT_2140( .ZN(I3310), .A(g1640) );
  INV_X1 NOT_2141( .ZN(g6897), .A(I9158) );
  INV_X1 NOT_2142( .ZN(g1837), .A(I2925) );
  INV_X1 NOT_2143( .ZN(I8755), .A(g6561) );
  INV_X1 NOT_2144( .ZN(g3460), .A(g2667) );
  INV_X1 NOT_2145( .ZN(I8226), .A(g6328) );
  INV_X1 NOT_2146( .ZN(g6425), .A(I8285) );
  INV_X1 NOT_2147( .ZN(g2135), .A(I3261) );
  INV_X1 NOT_2148( .ZN(I4510), .A(g2753) );
  INV_X1 NOT_2149( .ZN(I9146), .A(g6890) );
  INV_X1 NOT_2150( .ZN(g4110), .A(I5412) );
  INV_X1 NOT_2151( .ZN(I7167), .A(g5434) );
  INV_X1 NOT_2152( .ZN(I7318), .A(g5452) );
  INV_X4 NOT_2153( .ZN(I4291), .A(g2241) );
  INV_X4 NOT_2154( .ZN(g5894), .A(g5731) );
  INV_X1 NOT_2155( .ZN(g2805), .A(g2443) );
  INV_X1 NOT_2156( .ZN(g910), .A(I1938) );
  INV_X1 NOT_2157( .ZN(g1788), .A(g985) );
  INV_X1 NOT_2158( .ZN(g2422), .A(I3560) );
  INV_X1 NOT_2159( .ZN(I6772), .A(g4788) );
  INV_X1 NOT_2160( .ZN(I7193), .A(g5466) );
  INV_X1 NOT_2161( .ZN(I8491), .A(g6480) );
  INV_X1 NOT_2162( .ZN(g3079), .A(I4312) );
  INV_X1 NOT_2163( .ZN(I6531), .A(g4704) );
  INV_X1 NOT_2164( .ZN(g4402), .A(g4017) );
  INV_X1 NOT_2165( .ZN(g784), .A(I1862) );
  INV_X1 NOT_2166( .ZN(g1249), .A(I2240) );
  INV_X1 NOT_2167( .ZN(g4824), .A(g4615) );
  INV_X1 NOT_2168( .ZN(g837), .A(g353) );
  INV_X1 NOT_2169( .ZN(g5661), .A(g5518) );
  INV_X1 NOT_2170( .ZN(g3840), .A(I5043) );
  INV_X1 NOT_2171( .ZN(g719), .A(I1835) );
  INV_X1 NOT_2172( .ZN(I3590), .A(g1781) );
  INV_X1 NOT_2173( .ZN(g6406), .A(I8232) );
  INV_X1 NOT_2174( .ZN(g5475), .A(I7161) );
  INV_X1 NOT_2175( .ZN(I7686), .A(g5705) );
  INV_X1 NOT_2176( .ZN(g1842), .A(g1612) );
  INV_X1 NOT_2177( .ZN(I2721), .A(g1219) );
  INV_X1 NOT_2178( .ZN(g1192), .A(g44) );
  INV_X1 NOT_2179( .ZN(I8459), .A(g6427) );
  INV_X1 NOT_2180( .ZN(g6105), .A(I7811) );
  INV_X1 NOT_2181( .ZN(g6087), .A(g5813) );
  INV_X1 NOT_2182( .ZN(g6801), .A(I8969) );
  INV_X1 NOT_2183( .ZN(g6305), .A(I8027) );
  INV_X1 NOT_2184( .ZN(g5292), .A(I6942) );
  INV_X1 NOT_2185( .ZN(I8767), .A(g6619) );
  INV_X1 NOT_2186( .ZN(g6487), .A(g6365) );
  INV_X1 NOT_2187( .ZN(I3556), .A(g1484) );
  INV_X1 NOT_2188( .ZN(g3501), .A(g2650) );
  INV_X1 NOT_2189( .ZN(I3222), .A(g1790) );
  INV_X1 NOT_2190( .ZN(I8535), .A(g6447) );
  INV_X1 NOT_2191( .ZN(g4657), .A(I6244) );
  INV_X1 NOT_2192( .ZN(I8582), .A(g6439) );
  INV_X1 NOT_2193( .ZN(g1854), .A(I2958) );
  INV_X1 NOT_2194( .ZN(I9116), .A(g6864) );
  INV_X1 NOT_2195( .ZN(I8261), .A(g6298) );
  INV_X1 NOT_2196( .ZN(g5084), .A(g4727) );
  INV_X1 NOT_2197( .ZN(g4222), .A(I5654) );
  INV_X1 NOT_2198( .ZN(g2437), .A(I3572) );
  INV_X1 NOT_2199( .ZN(g2653), .A(I3797) );
  INV_X1 NOT_2200( .ZN(I6992), .A(g5151) );
  INV_X1 NOT_2201( .ZN(I1932), .A(g667) );
  INV_X1 NOT_2202( .ZN(g2102), .A(I3222) );
  INV_X1 NOT_2203( .ZN(g5439), .A(g5261) );
  INV_X1 NOT_2204( .ZN(I3785), .A(g2346) );
  INV_X1 NOT_2205( .ZN(I2940), .A(g1653) );
  INV_X1 NOT_2206( .ZN(I5837), .A(g3850) );
  INV_X1 NOT_2207( .ZN(g2869), .A(g2433) );
  INV_X1 NOT_2208( .ZN(I2388), .A(g878) );
  INV_X1 NOT_2209( .ZN(I6573), .A(g4721) );
  INV_X1 NOT_2210( .ZN(I3563), .A(g1461) );
  INV_X1 NOT_2211( .ZN(g5702), .A(I7463) );
  INV_X1 NOT_2212( .ZN(I8246), .A(g6290) );
  INV_X1 NOT_2213( .ZN(g1219), .A(I2218) );
  INV_X1 NOT_2214( .ZN(g1640), .A(I2601) );
  INV_X1 NOT_2215( .ZN(g2752), .A(g2343) );
  INV_X1 NOT_2216( .ZN(g6373), .A(I8183) );
  INV_X1 NOT_2217( .ZN(g3363), .A(g3110) );
  INV_X1 NOT_2218( .ZN(g6491), .A(g6373) );
  INV_X1 NOT_2219( .ZN(g5919), .A(I7689) );
  INV_X1 NOT_2220( .ZN(I2671), .A(g1017) );
  INV_X1 NOT_2221( .ZN(g1812), .A(I2867) );
  INV_X1 NOT_2222( .ZN(I8721), .A(g6534) );
  INV_X1 NOT_2223( .ZN(I2428), .A(g774) );
  INV_X1 NOT_2224( .ZN(g4563), .A(g4190) );
  INV_X1 NOT_2225( .ZN(g3053), .A(I4276) );
  INV_X1 NOT_2226( .ZN(g1176), .A(I2190) );
  INV_X1 NOT_2227( .ZN(g2265), .A(I3408) );
  INV_X1 NOT_2228( .ZN(g3453), .A(g2628) );
  INV_X1 NOT_2229( .ZN(g6283), .A(I7999) );
  INV_X1 NOT_2230( .ZN(g6369), .A(I8171) );
  INV_X1 NOT_2231( .ZN(g2042), .A(I3155) );
  INV_X1 NOT_2232( .ZN(g6602), .A(I8674) );
  INV_X1 NOT_2233( .ZN(I5249), .A(g3589) );
  INV_X2 NOT_2234( .ZN(g6407), .A(I8235) );
  INV_X1 NOT_2235( .ZN(g6578), .A(g6489) );
  INV_X1 NOT_2236( .ZN(g4844), .A(I6540) );
  INV_X1 NOT_2237( .ZN(g2164), .A(I3291) );
  INV_X1 NOT_2238( .ZN(g1286), .A(g854) );
  INV_X1 NOT_2239( .ZN(g2364), .A(I3516) );
  INV_X1 NOT_2240( .ZN(g2233), .A(I3364) );
  INV_X1 NOT_2241( .ZN(g4194), .A(I5612) );
  INV_X1 NOT_2242( .ZN(g1911), .A(I3010) );
  INV_X1 NOT_2243( .ZN(g4394), .A(I5885) );
  INV_X1 NOT_2244( .ZN(g6535), .A(I8521) );
  INV_X1 NOT_2245( .ZN(I6976), .A(g5136) );
  INV_X1 NOT_2246( .ZN(g3912), .A(g3505) );
  INV_X1 NOT_2247( .ZN(I2741), .A(g1222) );
  INV_X1 NOT_2248( .ZN(g5527), .A(I7267) );
  INV_X1 NOT_2249( .ZN(g6582), .A(I8614) );
  INV_X1 NOT_2250( .ZN(I8940), .A(g6783) );
  INV_X1 NOT_2251( .ZN(g4731), .A(I6359) );
  INV_X1 NOT_2252( .ZN(I2910), .A(g1645) );
  INV_X1 NOT_2253( .ZN(I3071), .A(g1504) );
  INV_X1 NOT_2254( .ZN(g5647), .A(g5509) );
  INV_X1 NOT_2255( .ZN(I3705), .A(g2316) );
  INV_X1 NOT_2256( .ZN(I3471), .A(g1450) );
  INV_X1 NOT_2257( .ZN(g2296), .A(I3441) );
  INV_X1 NOT_2258( .ZN(g1733), .A(I2741) );
  INV_X1 NOT_2259( .ZN(I2638), .A(g1123) );
  INV_X1 NOT_2260( .ZN(g1270), .A(g844) );
  INV_X1 NOT_2261( .ZN(g5546), .A(g5388) );
  INV_X1 NOT_2262( .ZN(I5854), .A(g3857) );
  INV_X1 NOT_2263( .ZN(I4465), .A(g2945) );
  INV_X1 NOT_2264( .ZN(g6015), .A(g5857) );
  INV_X1 NOT_2265( .ZN(g4705), .A(I6305) );
  INV_X1 NOT_2266( .ZN(g6415), .A(I8255) );
  INV_X1 NOT_2267( .ZN(I6126), .A(g4240) );
  INV_X1 NOT_2268( .ZN(I6400), .A(g4473) );
  INV_X1 NOT_2269( .ZN(g4242), .A(I5686) );
  INV_X1 NOT_2270( .ZN(I2883), .A(g1143) );
  INV_X1 NOT_2271( .ZN(I8671), .A(g6519) );
  INV_X1 NOT_2272( .ZN(g5925), .A(I7707) );
  INV_X1 NOT_2273( .ZN(I8030), .A(g6239) );
  INV_X1 NOT_2274( .ZN(I4433), .A(g2103) );
  INV_X1 NOT_2275( .ZN(g1324), .A(I2327) );
  INV_X1 NOT_2276( .ZN(I5708), .A(g3942) );
  INV_X1 NOT_2277( .ZN(I5520), .A(g3835) );
  INV_X1 NOT_2278( .ZN(g6721), .A(I8857) );
  INV_X1 NOT_2279( .ZN(I5640), .A(g3770) );
  INV_X1 NOT_2280( .ZN(g5120), .A(I6772) );
  INV_X1 NOT_2281( .ZN(I8564), .A(g6429) );
  INV_X1 NOT_2282( .ZN(g2706), .A(I3861) );
  INV_X1 NOT_2283( .ZN(I5252), .A(g3546) );
  INV_X1 NOT_2284( .ZN(I3773), .A(g2524) );
  INV_X1 NOT_2285( .ZN(g1177), .A(I2193) );
  INV_X1 NOT_2286( .ZN(g4150), .A(I5532) );
  INV_X1 NOT_2287( .ZN(I2165), .A(g690) );
  INV_X1 NOT_2288( .ZN(g1206), .A(I2212) );
  INV_X1 NOT_2289( .ZN(g4350), .A(g4010) );
  INV_X2 NOT_2290( .ZN(g2888), .A(g1972) );
  INV_X2 NOT_2291( .ZN(I7358), .A(g5565) );
  INV_X1 NOT_2292( .ZN(I4195), .A(g2173) );
  INV_X1 NOT_2293( .ZN(g2029), .A(I3134) );
  INV_X1 NOT_2294( .ZN(I7506), .A(g5584) );
  INV_X1 NOT_2295( .ZN(I5376), .A(g4014) );
  INV_X1 NOT_2296( .ZN(g2171), .A(I3304) );
  INV_X1 NOT_2297( .ZN(I4337), .A(g1934) );
  INV_X1 NOT_2298( .ZN(I8910), .A(g6730) );
  INV_X1 NOT_2299( .ZN(g2787), .A(g2405) );
  INV_X1 NOT_2300( .ZN(g6502), .A(I8426) );
  INV_X1 NOT_2301( .ZN(g2956), .A(g1861) );
  INV_X1 NOT_2302( .ZN(I6023), .A(g4151) );
  INV_X1 NOT_2303( .ZN(I8638), .A(g6553) );
  INV_X1 NOT_2304( .ZN(g1287), .A(g855) );
  INV_X1 NOT_2305( .ZN(g2675), .A(I3819) );
  INV_X1 NOT_2306( .ZN(I3836), .A(g1832) );
  INV_X4 NOT_2307( .ZN(I3212), .A(g1806) );
  INV_X1 NOT_2308( .ZN(I7587), .A(g5605) );
  INV_X1 NOT_2309( .ZN(g6940), .A(I9233) );
  INV_X1 NOT_2310( .ZN(g4769), .A(g4606) );
  INV_X1 NOT_2311( .ZN(g1849), .A(I2949) );
  INV_X1 NOT_2312( .ZN(g3778), .A(g3388) );
  INV_X1 NOT_2313( .ZN(g6188), .A(g5950) );
  INV_X1 NOT_2314( .ZN(I2196), .A(g3) );
  INV_X1 NOT_2315( .ZN(g5299), .A(I6949) );
  INV_X1 NOT_2316( .ZN(g1781), .A(I2825) );
  INV_X1 NOT_2317( .ZN(I6051), .A(g4185) );
  INV_X1 NOT_2318( .ZN(g1898), .A(I2995) );
  INV_X1 NOT_2319( .ZN(g3782), .A(g3388) );
  INV_X1 NOT_2320( .ZN(I8217), .A(g6319) );
  INV_X1 NOT_2321( .ZN(I8758), .A(g6562) );
  INV_X1 NOT_2322( .ZN(I8066), .A(g6114) );
  INV_X1 NOT_2323( .ZN(g5892), .A(g5742) );
  INV_X1 NOT_2324( .ZN(I6327), .A(g4451) );
  INV_X1 NOT_2325( .ZN(g6428), .A(I8290) );
  INV_X1 NOT_2326( .ZN(g3075), .A(I4306) );
  INV_X1 NOT_2327( .ZN(g4229), .A(g4059) );
  INV_X1 NOT_2328( .ZN(g2109), .A(I3235) );
  INV_X1 NOT_2329( .ZN(I7284), .A(g5383) );
  INV_X1 NOT_2330( .ZN(I4255), .A(g2179) );
  INV_X1 NOT_2331( .ZN(I6346), .A(g4563) );
  INV_X1 NOT_2332( .ZN(I8165), .A(g6189) );
  INV_X1 NOT_2333( .ZN(g4822), .A(g4614) );
  INV_X1 NOT_2334( .ZN(g1291), .A(I2278) );
  INV_X1 NOT_2335( .ZN(I5124), .A(g3719) );
  INV_X2 NOT_2336( .ZN(I2067), .A(g686) );
  INV_X2 NOT_2337( .ZN(g6564), .A(I8576) );
  INV_X1 NOT_2338( .ZN(I5324), .A(g3466) );
  INV_X1 NOT_2339( .ZN(I7832), .A(g5943) );
  INV_X1 NOT_2340( .ZN(g6826), .A(I9011) );
  INV_X1 NOT_2341( .ZN(I5469), .A(g3838) );
  INV_X1 NOT_2342( .ZN(I2290), .A(g971) );
  INV_X1 NOT_2343( .ZN(g1344), .A(I2379) );
  INV_X1 NOT_2344( .ZN(I4354), .A(g1953) );
  INV_X1 NOT_2345( .ZN(g5140), .A(I6798) );
  INV_X1 NOT_2346( .ZN(I5177), .A(g3267) );
  INV_X1 NOT_2347( .ZN(g3084), .A(I4321) );
  INV_X1 NOT_2348( .ZN(g5478), .A(I7170) );
  INV_X1 NOT_2349( .ZN(g1819), .A(I2877) );
  INV_X1 NOT_2350( .ZN(I6753), .A(g4772) );
  INV_X1 NOT_2351( .ZN(g2957), .A(g1861) );
  INV_X1 NOT_2352( .ZN(I8803), .A(g6685) );
  INV_X1 NOT_2353( .ZN(g1088), .A(I2119) );
  INV_X1 NOT_2354( .ZN(g1852), .A(I2952) );
  INV_X4 NOT_2355( .ZN(I6072), .A(g4385) );
  INV_X4 NOT_2356( .ZN(g6609), .A(I8693) );
  INV_X1 NOT_2357( .ZN(g5435), .A(I7113) );
  INV_X1 NOT_2358( .ZN(g6308), .A(I8034) );
  INV_X1 NOT_2359( .ZN(I3062), .A(g1776) );
  INV_X1 NOT_2360( .ZN(g5082), .A(g4723) );
  INV_X1 NOT_2361( .ZN(g2449), .A(I3584) );
  INV_X1 NOT_2362( .ZN(I3620), .A(g1484) );
  INV_X1 NOT_2363( .ZN(I3462), .A(g1450) );
  INV_X1 NOT_2364( .ZN(I8538), .A(g6450) );
  INV_X1 NOT_2365( .ZN(g2575), .A(I3684) );
  INV_X1 NOT_2366( .ZN(g2865), .A(g2296) );
  INV_X1 NOT_2367( .ZN(g6883), .A(I9116) );
  INV_X1 NOT_2368( .ZN(g5876), .A(I7640) );
  INV_X1 NOT_2369( .ZN(g4837), .A(g4473) );
  INV_X1 NOT_2370( .ZN(I8509), .A(g6437) );
  INV_X1 NOT_2371( .ZN(I2700), .A(g1173) );
  INV_X1 NOT_2372( .ZN(g2604), .A(I3736) );
  INV_X1 NOT_2373( .ZN(I4267), .A(g2525) );
  INV_X1 NOT_2374( .ZN(g2098), .A(g1363) );
  INV_X1 NOT_2375( .ZN(I4312), .A(g2555) );
  INV_X1 NOT_2376( .ZN(g4620), .A(g4251) );
  INV_X1 NOT_2377( .ZN(g4462), .A(I5977) );
  INV_X1 NOT_2378( .ZN(g6589), .A(I8635) );
  INV_X1 NOT_2379( .ZN(g945), .A(g536) );
  INV_X1 NOT_2380( .ZN(I8662), .A(g6525) );
  INV_X1 NOT_2381( .ZN(I3788), .A(g2554) );
  INV_X1 NOT_2382( .ZN(g6466), .A(I8332) );
  INV_X1 NOT_2383( .ZN(g5915), .A(I7679) );
  INV_X1 NOT_2384( .ZN(g3952), .A(I5182) );
  INV_X2 NOT_2385( .ZN(I6434), .A(g4622) );
  INV_X2 NOT_2386( .ZN(I8467), .A(g6457) );
  INV_X1 NOT_2387( .ZN(I8994), .A(g6789) );
  INV_X1 NOT_2388( .ZN(I8290), .A(g6291) );
  INV_X1 NOT_2389( .ZN(g1114), .A(I2150) );
  INV_X1 NOT_2390( .ZN(g6165), .A(g5926) );
  INV_X1 NOT_2391( .ZN(g6571), .A(I8597) );
  INV_X1 NOT_2392( .ZN(g6365), .A(I8159) );
  INV_X1 NOT_2393( .ZN(g2584), .A(I3705) );
  INV_X1 NOT_2394( .ZN(g4788), .A(I6452) );
  INV_X1 NOT_2395( .ZN(g6048), .A(g5824) );
  INV_X1 NOT_2396( .ZN(I1841), .A(g207) );
  INV_X1 NOT_2397( .ZN(g6711), .A(I8843) );
  INV_X1 NOT_2398( .ZN(I8093), .A(g6122) );
  INV_X1 NOT_2399( .ZN(g5110), .A(I6740) );
  INV_X1 NOT_2400( .ZN(g4249), .A(I5699) );
  INV_X1 NOT_2401( .ZN(g5310), .A(g5067) );
  INV_X1 NOT_2402( .ZN(I3298), .A(g1725) );
  INV_X1 NOT_2403( .ZN(g1825), .A(I2893) );
  INV_X1 NOT_2404( .ZN(g6827), .A(I9014) );
  INV_X1 NOT_2405( .ZN(g1650), .A(I2627) );
  INV_X1 NOT_2406( .ZN(I3485), .A(g1450) );
  INV_X2 NOT_2407( .ZN(g3527), .A(I4743) );
  INV_X1 NOT_2408( .ZN(g809), .A(I1874) );
  INV_X1 NOT_2409( .ZN(I6697), .A(g4722) );
  INV_X1 NOT_2410( .ZN(g4842), .A(I6534) );
  INV_X1 NOT_2411( .ZN(g849), .A(g598) );
  INV_X1 NOT_2412( .ZN(g2268), .A(I3419) );
  INV_X1 NOT_2413( .ZN(g4192), .A(I5606) );
  INV_X1 NOT_2414( .ZN(g4392), .A(I5879) );
  INV_X1 NOT_2415( .ZN(g3546), .A(g3095) );
  INV_X1 NOT_2416( .ZN(g4485), .A(I5987) );
  INV_X1 NOT_2417( .ZN(I2817), .A(g1222) );
  INV_X1 NOT_2418( .ZN(g5824), .A(g5631) );
  INV_X1 NOT_2419( .ZN(g1336), .A(I2361) );
  INV_X1 NOT_2420( .ZN(g6803), .A(I8975) );
  INV_X1 NOT_2421( .ZN(g3970), .A(I5236) );
  INV_X1 NOT_2422( .ZN(g1594), .A(g1143) );
  INV_X1 NOT_2423( .ZN(g4854), .A(I6570) );
  INV_X2 NOT_2424( .ZN(g6538), .A(g6469) );
  INV_X1 NOT_2425( .ZN(g1972), .A(I3083) );
  INV_X1 NOT_2426( .ZN(I5923), .A(g4299) );
  INV_X1 NOT_2427( .ZN(g6509), .A(I8447) );
  INV_X1 NOT_2428( .ZN(g1806), .A(I2857) );
  INV_X1 NOT_2429( .ZN(g5877), .A(I7643) );
  INV_X1 NOT_2430( .ZN(g5590), .A(I7352) );
  INV_X1 NOT_2431( .ZN(g1943), .A(I3050) );
  INV_X1 NOT_2432( .ZN(I3708), .A(g1946) );
  INV_X1 NOT_2433( .ZN(g3224), .A(I4471) );
  INV_X1 NOT_2434( .ZN(g2086), .A(I3198) );
  INV_X1 NOT_2435( .ZN(g2728), .A(I3890) );
  INV_X1 NOT_2436( .ZN(I3031), .A(g1504) );
  INV_X1 NOT_2437( .ZN(I4468), .A(g2583) );
  INV_X1 NOT_2438( .ZN(g3320), .A(g3067) );
  INV_X1 NOT_2439( .ZN(g6067), .A(g5788) );
  INV_X4 NOT_2440( .ZN(g1887), .A(I2982) );
  INV_X4 NOT_2441( .ZN(I3431), .A(g1275) );
  INV_X1 NOT_2442( .ZN(g1122), .A(I2162) );
  INV_X1 NOT_2443( .ZN(g6418), .A(I8264) );
  INV_X1 NOT_2444( .ZN(g6467), .A(I8335) );
  INV_X1 NOT_2445( .ZN(g1322), .A(I2321) );
  INV_X1 NOT_2446( .ZN(g4520), .A(I6072) );
  INV_X1 NOT_2447( .ZN(g1934), .A(I3037) );
  INV_X1 NOT_2448( .ZN(I2041), .A(g680) );
  INV_X1 NOT_2449( .ZN(I3376), .A(g1328) );
  INV_X1 NOT_2450( .ZN(g4431), .A(I5938) );
  INV_X1 NOT_2451( .ZN(g4252), .A(I5708) );
  INV_X1 NOT_2452( .ZN(I1874), .A(g282) );
  INV_X1 NOT_2453( .ZN(I3405), .A(g1321) );
  INV_X1 NOT_2454( .ZN(g3906), .A(g3575) );
  INV_X1 NOT_2455( .ZN(g2470), .A(I3602) );
  INV_X1 NOT_2456( .ZN(g3789), .A(g3388) );
  INV_X1 NOT_2457( .ZN(g5064), .A(I6706) );
  INV_X1 NOT_2458( .ZN(g2025), .A(g1276) );
  INV_X1 NOT_2459( .ZN(g6493), .A(g6375) );
  INV_X1 NOT_2460( .ZN(g5899), .A(g5753) );
  INV_X1 NOT_2461( .ZN(I6775), .A(g4790) );
  INV_X1 NOT_2462( .ZN(g4376), .A(I5843) );
  INV_X1 NOT_2463( .ZN(g4405), .A(I5910) );
  INV_X1 NOT_2464( .ZN(g3771), .A(I4964) );
  INV_X1 NOT_2465( .ZN(I5825), .A(g3914) );
  INV_X1 NOT_2466( .ZN(g872), .A(g143) );
  INV_X1 NOT_2467( .ZN(g1550), .A(g996) );
  INV_X1 NOT_2468( .ZN(I6060), .A(g4380) );
  INV_X1 NOT_2469( .ZN(g4286), .A(I5743) );
  INV_X1 NOT_2470( .ZN(g4765), .A(I6403) );
  INV_X1 NOT_2471( .ZN(I1880), .A(g276) );
  INV_X1 NOT_2472( .ZN(I4198), .A(g2276) );
  INV_X4 NOT_2473( .ZN(g3299), .A(g3049) );
  INV_X1 NOT_2474( .ZN(g5563), .A(g5381) );
  INV_X1 NOT_2475( .ZN(I4398), .A(g2086) );
  INV_X1 NOT_2476( .ZN(g4911), .A(I6615) );
  INV_X1 NOT_2477( .ZN(I3733), .A(g2031) );
  INV_X1 NOT_2478( .ZN(g6700), .A(I8818) );
  INV_X1 NOT_2479( .ZN(g1395), .A(I2428) );
  INV_X1 NOT_2480( .ZN(g1891), .A(I2986) );
  INV_X1 NOT_2481( .ZN(g1337), .A(I2364) );
  INV_X1 NOT_2482( .ZN(g5237), .A(g5083) );
  INV_X1 NOT_2483( .ZN(g3892), .A(g3575) );
  INV_X1 NOT_2484( .ZN(g2678), .A(g2312) );
  INV_X1 NOT_2485( .ZN(I3225), .A(g1813) );
  INV_X1 NOT_2486( .ZN(g6421), .A(I8273) );
  INV_X1 NOT_2487( .ZN(I2890), .A(g1123) );
  INV_X1 NOT_2488( .ZN(I8585), .A(g6442) );
  INV_X1 NOT_2489( .ZN(I5594), .A(g3821) );
  INV_X1 NOT_2490( .ZN(g4270), .A(I5723) );
  INV_X1 NOT_2491( .ZN(I7372), .A(g5493) );
  INV_X1 NOT_2492( .ZN(g1807), .A(I2860) );
  INV_X1 NOT_2493( .ZN(g4225), .A(g4059) );
  INV_X1 NOT_2494( .ZN(g2682), .A(I3826) );
  INV_X1 NOT_2495( .ZN(g2766), .A(g2361) );
  INV_X1 NOT_2496( .ZN(I6995), .A(g5220) );
  INV_X1 NOT_2497( .ZN(I1935), .A(g666) );
  INV_X1 NOT_2498( .ZN(g2087), .A(g1352) );
  INV_X1 NOT_2499( .ZN(g2105), .A(g1375) );
  INV_X1 NOT_2500( .ZN(I6937), .A(g5124) );
  INV_X4 NOT_2501( .ZN(I7143), .A(g5323) );
  INV_X4 NOT_2502( .ZN(I8441), .A(g6419) );
  INV_X1 NOT_2503( .ZN(g2801), .A(I4003) );
  INV_X1 NOT_2504( .ZN(I2411), .A(g736) );
  INV_X1 NOT_2505( .ZN(g5089), .A(I6723) );
  INV_X1 NOT_2506( .ZN(g5489), .A(I7187) );
  INV_X1 NOT_2507( .ZN(I5065), .A(g3714) );
  INV_X1 NOT_2508( .ZN(g4124), .A(I5454) );
  INV_X1 NOT_2509( .ZN(g714), .A(g131) );
  INV_X1 NOT_2510( .ZN(I3540), .A(g1670) );
  INV_X1 NOT_2511( .ZN(g4980), .A(g4678) );
  INV_X1 NOT_2512( .ZN(g2748), .A(I3923) );
  INV_X1 NOT_2513( .ZN(g6562), .A(I8570) );
  INV_X1 NOT_2514( .ZN(I3206), .A(g1823) );
  INV_X1 NOT_2515( .ZN(g5705), .A(I7466) );
  INV_X1 NOT_2516( .ZN(I2992), .A(g1741) );
  INV_X1 NOT_2517( .ZN(g3478), .A(g2695) );
  INV_X1 NOT_2518( .ZN(g1142), .A(I2169) );
  INV_X1 NOT_2519( .ZN(g2755), .A(g2350) );
  INV_X1 NOT_2520( .ZN(I4258), .A(g2169) );
  INV_X1 NOT_2521( .ZN(g5242), .A(g5085) );
  INV_X1 NOT_2522( .ZN(I8168), .A(g6170) );
  INV_X4 NOT_2523( .ZN(g6723), .A(I8863) );
  INV_X4 NOT_2524( .ZN(g1255), .A(g161) );
  INV_X1 NOT_2525( .ZN(I5033), .A(g3527) );
  INV_X1 NOT_2526( .ZN(g6101), .A(I7799) );
  INV_X1 NOT_2527( .ZN(g6817), .A(I8988) );
  INV_X1 NOT_2528( .ZN(I5433), .A(g3728) );
  INV_X1 NOT_2529( .ZN(g4206), .A(I5626) );
  INV_X1 NOT_2530( .ZN(g3082), .A(I4315) );
  INV_X1 NOT_2531( .ZN(g3482), .A(g2713) );
  INV_X1 NOT_2532( .ZN(I8531), .A(g6444) );
  INV_X1 NOT_2533( .ZN(g1692), .A(I2696) );
  INV_X1 NOT_2534( .ZN(g6605), .A(I8681) );
  INV_X1 NOT_2535( .ZN(g1726), .A(I2728) );
  INV_X1 NOT_2536( .ZN(g3876), .A(I5109) );
  INV_X1 NOT_2537( .ZN(g2173), .A(I3310) );
  INV_X1 NOT_2538( .ZN(I6942), .A(g5124) );
  INV_X1 NOT_2539( .ZN(g2091), .A(g1355) );
  INV_X1 NOT_2540( .ZN(I5496), .A(g3839) );
  INV_X1 NOT_2541( .ZN(g1960), .A(I3071) );
  INV_X1 NOT_2542( .ZN(g2491), .A(I3620) );
  INV_X1 NOT_2543( .ZN(g5150), .A(I6816) );
  INV_X1 NOT_2544( .ZN(g4849), .A(I6555) );
  INV_X1 NOT_2545( .ZN(g2169), .A(I3298) );
  INV_X1 NOT_2546( .ZN(g2283), .A(I3428) );
  INV_X1 NOT_2547( .ZN(I7113), .A(g5295) );
  INV_X1 NOT_2548( .ZN(I8411), .A(g6415) );
  INV_X1 NOT_2549( .ZN(I5337), .A(g3564) );
  INV_X1 NOT_2550( .ZN(I5913), .A(g3751) );
  INV_X1 NOT_2551( .ZN(g2602), .A(g2061) );
  INV_X1 NOT_2552( .ZN(g6585), .A(I8623) );
  INV_X1 NOT_2553( .ZN(g2007), .A(g1411) );
  INV_X1 NOT_2554( .ZN(g5773), .A(I7514) );
  INV_X4 NOT_2555( .ZN(g4399), .A(I5896) );
  INV_X4 NOT_2556( .ZN(I3797), .A(g2125) );
  INV_X1 NOT_2557( .ZN(I6250), .A(g4514) );
  INV_X1 NOT_2558( .ZN(g2059), .A(g1402) );
  INV_X1 NOT_2559( .ZN(g2920), .A(g1947) );
  INV_X1 NOT_2560( .ZN(I4170), .A(g2157) );
  INV_X1 NOT_2561( .ZN(g4781), .A(I6437) );
  INV_X1 NOT_2562( .ZN(g6441), .A(I8309) );
  INV_X1 NOT_2563( .ZN(I8074), .A(g6118) );
  INV_X1 NOT_2564( .ZN(g2767), .A(g2364) );
  INV_X1 NOT_2565( .ZN(g4900), .A(I6607) );
  INV_X1 NOT_2566( .ZN(g1783), .A(I2831) );
  INV_X1 NOT_2567( .ZN(g3110), .A(I4358) );
  INV_X1 NOT_2568( .ZN(I4821), .A(g2877) );
  INV_X1 NOT_2569( .ZN(I2688), .A(g1030) );
  INV_X1 NOT_2570( .ZN(I2857), .A(g1161) );
  INV_X1 NOT_2571( .ZN(g2535), .A(I3653) );
  INV_X1 NOT_2572( .ZN(I3291), .A(g1714) );
  INV_X1 NOT_2573( .ZN(g1979), .A(I3090) );
  INV_X1 NOT_2574( .ZN(g1112), .A(g336) );
  INV_X1 NOT_2575( .ZN(g1267), .A(g843) );
  INV_X1 NOT_2576( .ZN(I7494), .A(g5691) );
  INV_X1 NOT_2577( .ZN(g4510), .A(I6042) );
  INV_X1 NOT_2578( .ZN(I3144), .A(g1319) );
  INV_X1 NOT_2579( .ZN(g5918), .A(I7686) );
  INV_X1 NOT_2580( .ZN(g1001), .A(I2044) );
  INV_X1 NOT_2581( .ZN(g3002), .A(g2215) );
  INV_X1 NOT_2582( .ZN(I8573), .A(g6435) );
  INV_X1 NOT_2583( .ZN(I8863), .A(g6700) );
  INV_X1 NOT_2584( .ZN(I4483), .A(g3082) );
  INV_X1 NOT_2585( .ZN(g1293), .A(I2284) );
  INV_X1 NOT_2586( .ZN(g6368), .A(I8168) );
  INV_X1 NOT_2587( .ZN(g4144), .A(I5514) );
  INV_X1 NOT_2588( .ZN(I8713), .A(g6522) );
  INV_X1 NOT_2589( .ZN(I7593), .A(g5605) );
  INV_X1 NOT_2590( .ZN(I3819), .A(g2044) );
  INV_X1 NOT_2591( .ZN(g3236), .A(I4507) );
  INV_X1 NOT_2592( .ZN(g1329), .A(I2340) );
  INV_X1 NOT_2593( .ZN(I3694), .A(g1811) );
  INV_X1 NOT_2594( .ZN(g1761), .A(I2788) );
  INV_X1 NOT_2595( .ZN(g857), .A(g170) );
  INV_X4 NOT_2596( .ZN(g5993), .A(g5872) );
  INV_X4 NOT_2597( .ZN(g6531), .A(I8509) );
  INV_X1 NOT_2598( .ZN(I5081), .A(g3589) );
  INV_X1 NOT_2599( .ZN(I3923), .A(g2581) );
  INV_X1 NOT_2600( .ZN(I4306), .A(g1898) );
  INV_X1 NOT_2601( .ZN(I2760), .A(g1193) );
  INV_X1 NOT_2602( .ZN(g2664), .A(I3808) );
  INV_X1 NOT_2603( .ZN(I5481), .A(g3866) );
  INV_X1 NOT_2604( .ZN(I3488), .A(g1295) );
  INV_X1 NOT_2605( .ZN(g6743), .A(I8907) );
  INV_X1 NOT_2606( .ZN(g6890), .A(I9137) );
  INV_X1 NOT_2607( .ZN(g1830), .A(I2904) );
  INV_X1 NOT_2608( .ZN(I5692), .A(g3942) );
  INV_X1 NOT_2609( .ZN(I7264), .A(g5458) );
  INV_X1 NOT_2610( .ZN(g4852), .A(I6564) );
  INV_X1 NOT_2611( .ZN(g6505), .A(I8435) );
  INV_X1 NOT_2612( .ZN(I3215), .A(g1820) );
  INV_X1 NOT_2613( .ZN(g1221), .A(g46) );
  INV_X1 NOT_2614( .ZN(g6411), .A(I8243) );
  INV_X1 NOT_2615( .ZN(g6734), .A(I8894) );
  INV_X1 NOT_2616( .ZN(g3222), .A(I4465) );
  INV_X1 NOT_2617( .ZN(I3886), .A(g2215) );
  INV_X1 NOT_2618( .ZN(I8857), .A(g6698) );
  INV_X1 NOT_2619( .ZN(g1703), .A(I2707) );
  INV_X1 NOT_2620( .ZN(I2608), .A(g1143) );
  INV_X1 NOT_2621( .ZN(g5921), .A(I7695) );
  INV_X1 NOT_2622( .ZN(g4215), .A(I5637) );
  INV_X1 NOT_2623( .ZN(I2779), .A(g1038) );
  INV_X1 NOT_2624( .ZN(I7996), .A(g6137) );
  INV_X4 NOT_2625( .ZN(g6074), .A(g5794) );
  INV_X4 NOT_2626( .ZN(g3064), .A(I4291) );
  INV_X4 NOT_2627( .ZN(g3785), .A(g3466) );
  INV_X1 NOT_2628( .ZN(g1624), .A(I2581) );
  INV_X1 NOT_2629( .ZN(g1953), .A(I3062) );
  INV_X1 NOT_2630( .ZN(I4003), .A(g2284) );
  INV_X1 NOT_2631( .ZN(g5895), .A(g5742) );
  INV_X1 NOT_2632( .ZN(g4114), .A(I5424) );
  INV_X1 NOT_2633( .ZN(g4314), .A(g4080) );
  INV_X1 NOT_2634( .ZN(I2588), .A(g1193) );
  INV_X1 NOT_2635( .ZN(I3650), .A(g1650) );
  INV_X1 NOT_2636( .ZN(g6080), .A(g5805) );
  INV_X1 NOT_2637( .ZN(I2361), .A(g1075) );
  INV_X1 NOT_2638( .ZN(g6573), .A(I8603) );
  INV_X1 NOT_2639( .ZN(I4391), .A(g2275) );
  INV_X1 NOT_2640( .ZN(g6713), .A(g6679) );
  INV_X1 NOT_2641( .ZN(I3408), .A(g1644) );
  INV_X1 NOT_2642( .ZN(g3237), .A(I4510) );
  INV_X1 NOT_2643( .ZN(I7835), .A(g5926) );
  INV_X1 NOT_2644( .ZN(I2327), .A(g1222) );
  INV_X1 NOT_2645( .ZN(g6569), .A(I8591) );
  INV_X1 NOT_2646( .ZN(g2030), .A(I3137) );
  INV_X1 NOT_2647( .ZN(g5788), .A(I7587) );
  INV_X1 NOT_2648( .ZN(g2430), .A(I3563) );
  INV_X1 NOT_2649( .ZN(I2346), .A(g1193) );
  INV_X1 NOT_2650( .ZN(g4136), .A(I5490) );
  INV_X1 NOT_2651( .ZN(I8183), .A(g6176) );
  INV_X1 NOT_2652( .ZN(I4223), .A(g2176) );
  INV_X1 NOT_2653( .ZN(I8220), .A(g6322) );
  INV_X1 NOT_2654( .ZN(g4768), .A(I6410) );
  INV_X1 NOT_2655( .ZN(g1848), .A(I2946) );
  INV_X1 NOT_2656( .ZN(I9140), .A(g6888) );
  INV_X1 NOT_2657( .ZN(g2826), .A(g2481) );
  INV_X1 NOT_2658( .ZN(g1699), .A(I2703) );
  INV_X1 NOT_2659( .ZN(g1747), .A(I2760) );
  INV_X1 NOT_2660( .ZN(g838), .A(g564) );
  INV_X1 NOT_2661( .ZN(I6075), .A(g4386) );
  INV_X1 NOT_2662( .ZN(I2696), .A(g1156) );
  INV_X1 NOT_2663( .ZN(I4757), .A(g2861) );
  INV_X1 NOT_2664( .ZN(I7799), .A(g5918) );
  INV_X1 NOT_2665( .ZN(I3065), .A(g1426) );
  INV_X1 NOT_2666( .ZN(g3557), .A(g2598) );
  INV_X1 NOT_2667( .ZN(I5746), .A(g4022) );
  INV_X1 NOT_2668( .ZN(g4806), .A(g4473) );
  INV_X1 NOT_2669( .ZN(g5392), .A(I7058) );
  INV_X1 NOT_2670( .ZN(I8423), .A(g6423) );
  INV_X1 NOT_2671( .ZN(I9035), .A(g6812) );
  INV_X1 NOT_2672( .ZN(I6949), .A(g5050) );
  INV_X1 NOT_2673( .ZN(g4943), .A(I6635) );
  INV_X1 NOT_2674( .ZN(I3465), .A(g1724) );
  INV_X1 NOT_2675( .ZN(I3322), .A(g1333) );
  INV_X1 NOT_2676( .ZN(I9082), .A(g6849) );
  INV_X1 NOT_2677( .ZN(g3705), .A(g3014) );
  INV_X1 NOT_2678( .ZN(I8588), .A(g6443) );
  INV_X1 NOT_2679( .ZN(I4522), .A(g2801) );
  INV_X1 NOT_2680( .ZN(I2753), .A(g1174) );
  INV_X1 NOT_2681( .ZN(g842), .A(g571) );
  INV_X1 NOT_2682( .ZN(I6292), .A(g4434) );
  INV_X1 NOT_2683( .ZN(I4315), .A(g2245) );
  INV_X1 NOT_2684( .ZN(g3242), .A(g3083) );
  INV_X1 NOT_2685( .ZN(g4122), .A(I5448) );
  INV_X1 NOT_2686( .ZN(g4228), .A(I5668) );
  INV_X1 NOT_2687( .ZN(g4322), .A(I5793) );
  INV_X4 NOT_2688( .ZN(I2240), .A(g19) );
  INV_X4 NOT_2689( .ZN(I1938), .A(g332) );
  INV_X4 NOT_2690( .ZN(g2108), .A(I3232) );
  INV_X1 NOT_2691( .ZN(g2609), .A(I3749) );
  INV_X1 NOT_2692( .ZN(I6646), .A(g4687) );
  INV_X1 NOT_2693( .ZN(g2308), .A(I3452) );
  INV_X1 NOT_2694( .ZN(I8665), .A(g6527) );
  INV_X1 NOT_2695( .ZN(I8051), .A(g6108) );
  INV_X1 NOT_2696( .ZN(I7153), .A(g5358) );
  INV_X1 NOT_2697( .ZN(g2883), .A(g1954) );
  INV_X1 NOT_2698( .ZN(I6084), .A(g4391) );
  INV_X1 NOT_2699( .ZN(I6039), .A(g4182) );
  INV_X1 NOT_2700( .ZN(I5068), .A(g3571) );
  INV_X1 NOT_2701( .ZN(I3096), .A(g1439) );
  INV_X1 NOT_2702( .ZN(g1644), .A(I2611) );
  INV_X1 NOT_2703( .ZN(I3496), .A(g1326) );
  INV_X1 NOT_2704( .ZN(g715), .A(g135) );
  INV_X1 NOT_2705( .ZN(I3550), .A(g1295) );
  INV_X1 NOT_2706( .ZN(I7802), .A(g5920) );
  INV_X1 NOT_2707( .ZN(g5708), .A(I7469) );
  INV_X1 NOT_2708( .ZN(g1119), .A(I2159) );
  INV_X1 NOT_2709( .ZN(g1319), .A(I2312) );
  INV_X1 NOT_2710( .ZN(g2066), .A(g1341) );
  INV_X1 NOT_2711( .ZN(g3150), .A(I4391) );
  INV_X1 NOT_2712( .ZN(g5219), .A(I6885) );
  INV_X1 NOT_2713( .ZN(I3137), .A(g1315) );
  INV_X1 NOT_2714( .ZN(I8103), .A(g6134) );
  INV_X1 NOT_2715( .ZN(I3395), .A(g1286) );
  INV_X1 NOT_2716( .ZN(I3337), .A(g1338) );
  INV_X1 NOT_2717( .ZN(g4496), .A(I6008) );
  INV_X1 NOT_2718( .ZN(g1352), .A(I2391) );
  INV_X1 NOT_2719( .ZN(I9110), .A(g6864) );
  INV_X1 NOT_2720( .ZN(g1577), .A(g1001) );
  INV_X1 NOT_2721( .ZN(g4550), .A(I6126) );
  INV_X1 NOT_2722( .ZN(g3773), .A(g3466) );
  INV_X1 NOT_2723( .ZN(g4845), .A(I6543) );
  INV_X1 NOT_2724( .ZN(I4537), .A(g2877) );
  INV_X1 NOT_2725( .ZN(I8696), .A(g6569) );
  INV_X1 NOT_2726( .ZN(g2165), .A(I3294) );
  INV_X1 NOT_2727( .ZN(g5958), .A(g5818) );
  INV_X1 NOT_2728( .ZN(I2147), .A(g6) );
  INV_X1 NOT_2729( .ZN(g6608), .A(I8690) );
  INV_X1 NOT_2730( .ZN(g4195), .A(I5615) );
  INV_X1 NOT_2731( .ZN(g4137), .A(I5493) );
  INV_X1 NOT_2732( .ZN(g830), .A(g338) );
  INV_X1 NOT_2733( .ZN(I5716), .A(g3942) );
  INV_X1 NOT_2734( .ZN(g3769), .A(g3622) );
  INV_X1 NOT_2735( .ZN(I9002), .A(g6802) );
  INV_X1 NOT_2736( .ZN(g2827), .A(g2485) );
  INV_X1 NOT_2737( .ZN(I6952), .A(g5124) );
  INV_X1 NOT_2738( .ZN(I5848), .A(g3856) );
  INV_X1 NOT_2739( .ZN(g3836), .A(I5033) );
  INV_X1 NOT_2740( .ZN(g3212), .A(I4455) );
  INV_X1 NOT_2741( .ZN(g6423), .A(I8279) );
  INV_X4 NOT_2742( .ZN(I4243), .A(g1853) );
  INV_X4 NOT_2743( .ZN(g2333), .A(I3485) );
  INV_X4 NOT_2744( .ZN(I8240), .A(g6287) );
  INV_X1 NOT_2745( .ZN(g1975), .A(I3086) );
  INV_X1 NOT_2746( .ZN(I5699), .A(g3844) );
  INV_X1 NOT_2747( .ZN(g4807), .A(g4473) );
  INV_X1 NOT_2748( .ZN(I9236), .A(g6939) );
  INV_X1 NOT_2749( .ZN(g3967), .A(I5223) );
  INV_X1 NOT_2750( .ZN(I6561), .A(g4707) );
  INV_X1 NOT_2751( .ZN(g6588), .A(I8632) );
  INV_X1 NOT_2752( .ZN(I4935), .A(g3369) );
  INV_X1 NOT_2753( .ZN(I2596), .A(g985) );
  INV_X1 NOT_2754( .ZN(g6161), .A(g5926) );
  INV_X1 NOT_2755( .ZN(g1274), .A(g856) );
  INV_X1 NOT_2756( .ZN(g6361), .A(I8147) );
  INV_X1 NOT_2757( .ZN(g1426), .A(I2445) );
  INV_X1 NOT_2758( .ZN(g2196), .A(I3337) );
  INV_X1 NOT_2759( .ZN(I7600), .A(g5605) );
  INV_X1 NOT_2760( .ZN(g2803), .A(g2440) );
  INV_X1 NOT_2761( .ZN(I6004), .A(g4159) );
  INV_X1 NOT_2762( .ZN(g3229), .A(I4486) );
  INV_X1 NOT_2763( .ZN(I6986), .A(g5230) );
  INV_X1 NOT_2764( .ZN(g6051), .A(g5824) );
  INV_X1 NOT_2765( .ZN(g5270), .A(I6927) );
  INV_X1 NOT_2766( .ZN(g804), .A(I1871) );
  INV_X1 NOT_2767( .ZN(I3255), .A(g1650) );
  INV_X1 NOT_2768( .ZN(g2538), .A(I3656) );
  INV_X1 NOT_2769( .ZN(g1325), .A(I2330) );
  INV_X1 NOT_2770( .ZN(g1821), .A(I2883) );
  INV_X4 NOT_2771( .ZN(g844), .A(g578) );
  INV_X1 NOT_2772( .ZN(I3481), .A(g1461) );
  INV_X1 NOT_2773( .ZN(I8034), .A(g6242) );
  INV_X1 NOT_2774( .ZN(g4142), .A(I5508) );
  INV_X1 NOT_2775( .ZN(g4248), .A(I5696) );
  INV_X1 NOT_2776( .ZN(g2509), .A(I3635) );
  INV_X1 NOT_2777( .ZN(I6546), .A(g4692) );
  INV_X1 NOT_2778( .ZN(I3726), .A(g2030) );
  INV_X1 NOT_2779( .ZN(g4815), .A(I6495) );
  INV_X1 NOT_2780( .ZN(I5644), .A(g4059) );
  INV_X1 NOT_2781( .ZN(I8147), .A(g6182) );
  INV_X1 NOT_2782( .ZN(g5124), .A(I6780) );
  INV_X1 NOT_2783( .ZN(g6103), .A(I7805) );
  INV_X1 NOT_2784( .ZN(I5119), .A(g3714) );
  INV_X1 NOT_2785( .ZN(g4692), .A(I6280) );
  INV_X1 NOT_2786( .ZN(g2467), .A(I3599) );
  INV_X1 NOT_2787( .ZN(I8681), .A(g6566) );
  INV_X1 NOT_2788( .ZN(g4726), .A(I6352) );
  INV_X1 NOT_2789( .ZN(g5469), .A(I7153) );
  INV_X1 NOT_2790( .ZN(g4154), .A(I5548) );
  INV_X4 NOT_2791( .ZN(I2601), .A(g1161) );
  INV_X4 NOT_2792( .ZN(g6696), .A(I8806) );
  INV_X1 NOT_2793( .ZN(g1636), .A(I2593) );
  INV_X1 NOT_2794( .ZN(g3921), .A(g3512) );
  INV_X1 NOT_2795( .ZN(g5540), .A(I7284) );
  INV_X1 NOT_2796( .ZN(I5577), .A(g4022) );
  INV_X1 NOT_2797( .ZN(g1106), .A(I2128) );
  INV_X1 NOT_2798( .ZN(g6732), .A(I8888) );
  INV_X1 NOT_2799( .ZN(g853), .A(g642) );
  INV_X1 NOT_2800( .ZN(g2256), .A(I3395) );
  INV_X1 NOT_2801( .ZN(g1790), .A(I2842) );
  INV_X1 NOT_2802( .ZN(I2922), .A(g1774) );
  INV_X1 NOT_2803( .ZN(g6508), .A(I8444) );
  INV_X1 NOT_2804( .ZN(I5893), .A(g3747) );
  INV_X1 NOT_2805( .ZN(I3979), .A(g1836) );
  INV_X1 NOT_2806( .ZN(I2581), .A(g946) );
  INV_X1 NOT_2807( .ZN(I3112), .A(g1439) );
  INV_X1 NOT_2808( .ZN(g1461), .A(I2460) );
  INV_X1 NOT_2809( .ZN(g3462), .A(g2679) );
  INV_X1 NOT_2810( .ZN(g1756), .A(I2779) );
  INV_X1 NOT_2811( .ZN(g2381), .A(I3528) );
  INV_X1 NOT_2812( .ZN(I6789), .A(g4871) );
  INV_X1 NOT_2813( .ZN(g4783), .A(I6441) );
  INV_X1 NOT_2814( .ZN(g6043), .A(g5824) );
  INV_X1 NOT_2815( .ZN(I7871), .A(g6097) );
  INV_X1 NOT_2816( .ZN(I2460), .A(g952) );
  INV_X1 NOT_2817( .ZN(I3001), .A(g1267) );
  INV_X1 NOT_2818( .ZN(g4112), .A(I5418) );
  INV_X1 NOT_2819( .ZN(g4218), .A(I5640) );
  INV_X1 NOT_2820( .ZN(g2197), .A(I3340) );
  INV_X2 NOT_2821( .ZN(g4267), .A(I5720) );
  INV_X1 NOT_2822( .ZN(I4166), .A(g2390) );
  INV_X1 NOT_2823( .ZN(g2397), .A(I3540) );
  INV_X1 NOT_2824( .ZN(I4366), .A(g2244) );
  INV_X1 NOT_2825( .ZN(g5199), .A(I6867) );
  INV_X1 NOT_2826( .ZN(g5399), .A(I7065) );
  INV_X1 NOT_2827( .ZN(g1046), .A(g489) );
  INV_X1 NOT_2828( .ZN(I3761), .A(g2505) );
  INV_X1 NOT_2829( .ZN(g3788), .A(g3466) );
  INV_X2 NOT_2830( .ZN(g6034), .A(g5824) );
  INV_X1 NOT_2831( .ZN(g6434), .A(I8300) );
  INV_X1 NOT_2832( .ZN(g6565), .A(I8579) );
  INV_X1 NOT_2833( .ZN(I6299), .A(g4438) );
  INV_X1 NOT_2834( .ZN(g4293), .A(I5750) );
  INV_X1 NOT_2835( .ZN(g4129), .A(I5469) );
  INV_X1 NOT_2836( .ZN(g5797), .A(I7596) );
  INV_X1 NOT_2837( .ZN(I3830), .A(g2179) );
  INV_X1 NOT_2838( .ZN(I2995), .A(g1742) );
  INV_X1 NOT_2839( .ZN(g6147), .A(I7871) );
  INV_X1 NOT_2840( .ZN(g1345), .A(I2382) );
  INV_X1 NOT_2841( .ZN(g1841), .A(I2929) );
  INV_X1 NOT_2842( .ZN(g6347), .A(I8103) );
  INV_X1 NOT_2843( .ZN(I1832), .A(g143) );
  INV_X1 NOT_2844( .ZN(I2479), .A(g1049) );
  INV_X1 NOT_2845( .ZN(I7339), .A(g5540) );
  INV_X1 NOT_2846( .ZN(g1191), .A(g38) );
  INV_X1 NOT_2847( .ZN(I2668), .A(g1011) );
  INV_X1 NOT_2848( .ZN(g1391), .A(I2424) );
  INV_X1 NOT_2849( .ZN(I1853), .A(g211) );
  INV_X1 NOT_2850( .ZN(g3192), .A(I4429) );
  INV_X1 NOT_2851( .ZN(g6533), .A(I8515) );
  INV_X1 NOT_2852( .ZN(g3085), .A(I4324) );
  INV_X1 NOT_2853( .ZN(I3746), .A(g2035) );
  INV_X1 NOT_2854( .ZN(I7838), .A(g5947) );
  INV_X4 NOT_2855( .ZN(g4727), .A(I6355) );
  INV_X4 NOT_2856( .ZN(I4964), .A(g3673) );
  INV_X1 NOT_2857( .ZN(g3485), .A(g2986) );
  INV_X1 NOT_2858( .ZN(I2190), .A(g297) );
  INV_X1 NOT_2859( .ZN(g1695), .A(g1106) );
  INV_X1 NOT_2860( .ZN(g6697), .A(I8809) );
  INV_X1 NOT_2861( .ZN(g1637), .A(I2596) );
  INV_X1 NOT_2862( .ZN(g1107), .A(I2131) );
  INV_X1 NOT_2863( .ZN(g2631), .A(I3773) );
  INV_X1 NOT_2864( .ZN(g6596), .A(I8656) );
  INV_X1 NOT_2865( .ZN(g3854), .A(I5071) );
  INV_X1 NOT_2866( .ZN(I5106), .A(g3247) );
  INV_X1 NOT_2867( .ZN(I8597), .A(g6445) );
  INV_X1 NOT_2868( .ZN(g2817), .A(g2461) );
  INV_X1 NOT_2869( .ZN(I6244), .A(g4519) );
  INV_X1 NOT_2870( .ZN(I7077), .A(g5281) );
  INV_X1 NOT_2871( .ZN(g4703), .A(I6299) );
  INV_X1 NOT_2872( .ZN(g6413), .A(I8249) );
  INV_X1 NOT_2873( .ZN(I5790), .A(g3803) );
  INV_X1 NOT_2874( .ZN(g1858), .A(I2964) );
  INV_X1 NOT_2875( .ZN(I6078), .A(g4387) );
  INV_X1 NOT_2876( .ZN(I6340), .A(g4561) );
  INV_X1 NOT_2877( .ZN(I7643), .A(g5752) );
  INV_X1 NOT_2878( .ZN(I3068), .A(g1439) );
  INV_X1 NOT_2879( .ZN(g5923), .A(I7701) );
  INV_X1 NOT_2880( .ZN(I9038), .A(g6833) );
  INV_X1 NOT_2881( .ZN(I3468), .A(g1802) );
  INV_X4 NOT_2882( .ZN(I4279), .A(g2230) );
  INV_X4 NOT_2883( .ZN(I5756), .A(g3922) );
  INV_X1 NOT_2884( .ZN(g6820), .A(I8997) );
  INV_X1 NOT_2885( .ZN(g4624), .A(g4265) );
  INV_X1 NOT_2886( .ZN(I6959), .A(g5089) );
  INV_X1 NOT_2887( .ZN(I5622), .A(g3914) );
  INV_X1 NOT_2888( .ZN(g3219), .A(I4462) );
  INV_X1 NOT_2889( .ZN(I5027), .A(g3267) );
  INV_X1 NOT_2890( .ZN(I4318), .A(g2171) );
  INV_X1 NOT_2891( .ZN(I7634), .A(g5727) );
  INV_X1 NOT_2892( .ZN(I5427), .A(g3726) );
  INV_X4 NOT_2893( .ZN(g3031), .A(I4246) );
  INV_X4 NOT_2894( .ZN(g1115), .A(g40) );
  INV_X1 NOT_2895( .ZN(g6117), .A(g5880) );
  INV_X1 NOT_2896( .ZN(g1315), .A(I2296) );
  INV_X1 NOT_2897( .ZN(g1811), .A(I2864) );
  INV_X1 NOT_2898( .ZN(g1642), .A(g809) );
  INV_X1 NOT_2899( .ZN(I8479), .A(g6482) );
  INV_X1 NOT_2900( .ZN(g2585), .A(I3708) );
  INV_X1 NOT_2901( .ZN(I7104), .A(g5273) );
  INV_X1 NOT_2902( .ZN(I5904), .A(g3749) );
  INV_X1 NOT_2903( .ZN(I8668), .A(g6530) );
  INV_X1 NOT_2904( .ZN(g5886), .A(g5753) );
  INV_X1 NOT_2905( .ZN(I8840), .A(g6657) );
  INV_X1 NOT_2906( .ZN(g2041), .A(I3152) );
  INV_X1 NOT_2907( .ZN(g6601), .A(I8671) );
  INV_X1 NOT_2908( .ZN(I5514), .A(g3882) );
  INV_X1 NOT_2909( .ZN(I3349), .A(g1334) );
  INV_X1 NOT_2910( .ZN(I2053), .A(g684) );
  INV_X1 NOT_2911( .ZN(g5114), .A(I6756) );
  INV_X1 NOT_2912( .ZN(I5403), .A(g3970) );
  INV_X1 NOT_2913( .ZN(g5314), .A(I6972) );
  INV_X1 NOT_2914( .ZN(I2453), .A(g952) );
  INV_X1 NOT_2915( .ZN(g1654), .A(g878) );
  INV_X1 NOT_2916( .ZN(g4716), .A(I6330) );
  INV_X1 NOT_2917( .ZN(g4149), .A(I5529) );
  INV_X1 NOT_2918( .ZN(g6922), .A(I9203) );
  INV_X8 NOT_2919( .ZN(I8156), .A(g6167) );
  INV_X1 NOT_2920( .ZN(I3198), .A(g1819) );
  INV_X1 NOT_2921( .ZN(I3855), .A(g2550) );
  INV_X1 NOT_2922( .ZN(I5391), .A(g3975) );
  INV_X1 NOT_2923( .ZN(g3911), .A(I5148) );
  INV_X1 NOT_2924( .ZN(g6581), .A(g6493) );
  INV_X1 NOT_2925( .ZN(g4848), .A(I6552) );
  INV_X1 NOT_2926( .ZN(I5637), .A(g3914) );
  INV_X1 NOT_2927( .ZN(g1880), .A(g1603) );
  INV_X1 NOT_2928( .ZN(g4198), .A(I5618) );
  INV_X1 NOT_2929( .ZN(g4699), .A(I6289) );
  INV_X1 NOT_2930( .ZN(g6597), .A(I8659) );
  INV_X1 NOT_2931( .ZN(g4855), .A(I6573) );
  INV_X1 NOT_2932( .ZN(g4398), .A(I5893) );
  INV_X1 NOT_2933( .ZN(g2772), .A(I3961) );
  INV_X1 NOT_2934( .ZN(I4321), .A(g1917) );
  INV_X1 NOT_2935( .ZN(g5136), .A(I6786) );
  INV_X1 NOT_2936( .ZN(g3225), .A(I4474) );
  INV_X1 NOT_2937( .ZN(I5223), .A(g3537) );
  INV_X1 NOT_2938( .ZN(g2743), .A(g2333) );
  INV_X1 NOT_2939( .ZN(g6784), .A(I8940) );
  INV_X1 NOT_2940( .ZN(g2890), .A(g1875) );
  INV_X1 NOT_2941( .ZN(g3073), .A(I4300) );
  INV_X1 NOT_2942( .ZN(g1978), .A(g1387) );
  INV_X1 NOT_2943( .ZN(g3796), .A(g3388) );
  INV_X1 NOT_2944( .ZN(g1017), .A(I2053) );
  INV_X1 NOT_2945( .ZN(I2929), .A(g1659) );
  INV_X2 NOT_2946( .ZN(g798), .A(I1868) );
  INV_X1 NOT_2947( .ZN(g2505), .A(I3629) );
  INV_X1 NOT_2948( .ZN(I3644), .A(g1685) );
  INV_X1 NOT_2949( .ZN(g3124), .A(I4371) );
  INV_X1 NOT_2950( .ZN(g1935), .A(I3040) );
  INV_X1 NOT_2951( .ZN(g3980), .A(I5264) );
  INV_X1 NOT_2952( .ZN(g2856), .A(g2010) );
  INV_X1 NOT_2953( .ZN(g2734), .A(I3902) );
  INV_X1 NOT_2954( .ZN(I8432), .A(g6411) );
  INV_X1 NOT_2955( .ZN(I3319), .A(g1636) );
  INV_X1 NOT_2956( .ZN(g1982), .A(I3093) );
  INV_X1 NOT_2957( .ZN(g754), .A(I1850) );
  INV_X1 NOT_2958( .ZN(g4524), .A(I6084) );
  INV_X1 NOT_2959( .ZN(g836), .A(g349) );
  INV_X1 NOT_2960( .ZN(I8453), .A(g6414) );
  INV_X1 NOT_2961( .ZN(g6840), .A(I9041) );
  INV_X1 NOT_2962( .ZN(I4519), .A(g2788) );
  INV_X1 NOT_2963( .ZN(g4644), .A(I6231) );
  INV_X1 NOT_2964( .ZN(I3152), .A(g1322) );
  INV_X1 NOT_2965( .ZN(I3258), .A(g1760) );
  INV_X1 NOT_2966( .ZN(g3540), .A(I4762) );
  INV_X1 NOT_2967( .ZN(I3352), .A(g1285) );
  INV_X1 NOT_2968( .ZN(g1328), .A(I2337) );
  INV_X1 NOT_2969( .ZN(g5887), .A(g5742) );
  INV_X1 NOT_2970( .ZN(g4119), .A(I5439) );
  INV_X1 NOT_2971( .ZN(g5465), .A(I7143) );
  INV_X4 NOT_2972( .ZN(g1542), .A(g878) );
  INV_X4 NOT_2973( .ZN(g1330), .A(I2343) );
  INV_X1 NOT_2974( .ZN(g3177), .A(I4414) );
  INV_X1 NOT_2975( .ZN(I3717), .A(g2154) );
  INV_X1 NOT_2976( .ZN(g5230), .A(I6895) );
  INV_X1 NOT_2977( .ZN(g845), .A(g582) );
  INV_X1 NOT_2978( .ZN(g4152), .A(I5542) );
  INV_X1 NOT_2979( .ZN(g6501), .A(I8423) );
  INV_X1 NOT_2980( .ZN(g4577), .A(g4202) );
  INV_X1 NOT_2981( .ZN(g4717), .A(g4465) );
  INV_X1 NOT_2982( .ZN(g5433), .A(I7107) );
  INV_X1 NOT_2983( .ZN(I5654), .A(g3742) );
  INV_X1 NOT_2984( .ZN(I6930), .A(g5017) );
  INV_X1 NOT_2985( .ZN(g2863), .A(g2296) );
  INV_X1 NOT_2986( .ZN(I6464), .A(g4562) );
  INV_X1 NOT_2987( .ZN(I3599), .A(g1484) );
  INV_X1 NOT_2988( .ZN(g2713), .A(I3868) );
  INV_X1 NOT_2989( .ZN(I3274), .A(g1773) );
  INV_X1 NOT_2990( .ZN(g4386), .A(I5865) );
  INV_X1 NOT_2991( .ZN(g3199), .A(g1861) );
  INV_X1 NOT_2992( .ZN(g5550), .A(g5331) );
  INV_X1 NOT_2993( .ZN(I3614), .A(g1295) );
  INV_X1 NOT_2994( .ZN(g3781), .A(I4976) );
  INV_X1 NOT_2995( .ZN(I3370), .A(g1805) );
  INV_X1 NOT_2996( .ZN(g5137), .A(I6789) );
  INV_X1 NOT_2997( .ZN(g5395), .A(I7061) );
  INV_X1 NOT_2998( .ZN(g5891), .A(g5731) );
  INV_X4 NOT_2999( .ZN(g3898), .A(g3575) );
  INV_X4 NOT_3000( .ZN(g3900), .A(g3575) );
  INV_X8 NOT_3001( .ZN(I3325), .A(g1340) );
  INV_X1 NOT_3002( .ZN(g4426), .A(I5929) );
  INV_X1 NOT_3003( .ZN(I2735), .A(g1118) );
  INV_X1 NOT_3004( .ZN(g3797), .A(g3388) );
  INV_X1 NOT_3005( .ZN(I9085), .A(g6850) );
  INV_X1 NOT_3006( .ZN(g1902), .A(I3001) );
  INV_X1 NOT_3007( .ZN(g6163), .A(g5926) );
  INV_X1 NOT_3008( .ZN(g4614), .A(g4308) );
  INV_X1 NOT_3009( .ZN(I2782), .A(g1177) );
  INV_X1 NOT_3010( .ZN(I7679), .A(g5726) );
  INV_X1 NOT_3011( .ZN(g6363), .A(I8153) );
  INV_X1 NOT_3012( .ZN(g4370), .A(I5831) );
  INV_X1 NOT_3013( .ZN(I8626), .A(g6543) );
  INV_X1 NOT_3014( .ZN(g3510), .A(g2709) );
  INV_X1 NOT_3015( .ZN(I5612), .A(g3910) );
  INV_X1 NOT_3016( .ZN(g6032), .A(g5770) );
  INV_X1 NOT_3017( .ZN(g4125), .A(I5457) );
  INV_X1 NOT_3018( .ZN(g2688), .A(I3836) );
  INV_X4 NOT_3019( .ZN(g2857), .A(I4059) );
  INV_X4 NOT_3020( .ZN(g3291), .A(g3037) );
  INV_X1 NOT_3021( .ZN(I3083), .A(g1426) );
  INV_X1 NOT_3022( .ZN(g2976), .A(g2197) );
  INV_X1 NOT_3023( .ZN(g1823), .A(I2887) );
  INV_X1 NOT_3024( .ZN(I2949), .A(g1263) );
  INV_X1 NOT_3025( .ZN(g1366), .A(I2402) );
  INV_X1 NOT_3026( .ZN(g5266), .A(I6923) );
  INV_X1 NOT_3027( .ZN(I2627), .A(g1053) );
  INV_X1 NOT_3028( .ZN(g1056), .A(g89) );
  INV_X1 NOT_3029( .ZN(g6568), .A(I8588) );
  INV_X1 NOT_3030( .ZN(I5328), .A(g3502) );
  INV_X1 NOT_3031( .ZN(g1529), .A(g1076) );
  INV_X1 NOT_3032( .ZN(I7805), .A(g5923) );
  INV_X1 NOT_3033( .ZN(I5542), .A(g3984) );
  INV_X1 NOT_3034( .ZN(I2998), .A(g1257) );
  INV_X1 NOT_3035( .ZN(g1649), .A(g985) );
  INV_X1 NOT_3036( .ZN(g1348), .A(I2385) );
  INV_X1 NOT_3037( .ZN(g3259), .A(g2996) );
  INV_X1 NOT_3038( .ZN(I4358), .A(g2525) );
  INV_X1 NOT_3039( .ZN(g5248), .A(g4911) );
  INV_X1 NOT_3040( .ZN(g4636), .A(g4286) );
  INV_X1 NOT_3041( .ZN(g1355), .A(I2394) );
  INV_X1 NOT_3042( .ZN(g4106), .A(I5400) );
  INV_X1 NOT_3043( .ZN(g5255), .A(g4933) );
  INV_X1 NOT_3044( .ZN(g3852), .A(I5065) );
  INV_X1 NOT_3045( .ZN(I9031), .A(g6809) );
  INV_X1 NOT_3046( .ZN(g2760), .A(I3942) );
  INV_X1 NOT_3047( .ZN(g3488), .A(g2728) );
  INV_X1 NOT_3048( .ZN(I8894), .A(g6709) );
  INV_X1 NOT_3049( .ZN(g4790), .A(I6456) );
  INV_X1 NOT_3050( .ZN(g5692), .A(I7451) );
  INV_X8 NOT_3051( .ZN(I4587), .A(g2962) );
  INV_X8 NOT_3052( .ZN(g5097), .A(I6733) );
  INV_X1 NOT_3053( .ZN(g5726), .A(I7487) );
  INV_X1 NOT_3054( .ZN(g4187), .A(I5591) );
  INV_X1 NOT_3055( .ZN(I9176), .A(g6881) );
  INV_X1 NOT_3056( .ZN(g4387), .A(I5868) );
  INV_X1 NOT_3057( .ZN(I9005), .A(g6817) );
  INV_X1 NOT_3058( .ZN(g1063), .A(g675) );
  INV_X1 NOT_3059( .ZN(g3886), .A(g3346) );
  INV_X1 NOT_3060( .ZN(g4622), .A(g4252) );
  INV_X1 NOT_3061( .ZN(g2608), .A(I3746) );
  INV_X2 NOT_3062( .ZN(I2919), .A(g1787) );
  INV_X1 NOT_3063( .ZN(g2779), .A(g2394) );
  INV_X1 NOT_3064( .ZN(g4904), .A(g4812) );
  INV_X1 NOT_3065( .ZN(g3114), .A(I4362) );
  INV_X1 NOT_3066( .ZN(I2952), .A(g1594) );
  INV_X1 NOT_3067( .ZN(g1279), .A(g848) );
  INV_X1 NOT_3068( .ZN(g4514), .A(I6054) );
  INV_X1 NOT_3069( .ZN(g1720), .A(g1111) );
  INV_X1 NOT_3070( .ZN(g4003), .A(g3441) );
  INV_X1 NOT_3071( .ZN(g1118), .A(g36) );
  INV_X1 NOT_3072( .ZN(I3391), .A(g1646) );
  INV_X1 NOT_3073( .ZN(g1318), .A(I2309) );
  INV_X1 NOT_3074( .ZN(g4403), .A(I5904) );
  INV_X1 NOT_3075( .ZN(I5490), .A(g3832) );
  INV_X1 NOT_3076( .ZN(g5112), .A(I6750) );
  INV_X1 NOT_3077( .ZN(g2588), .A(I3717) );
  INV_X1 NOT_3078( .ZN(g4145), .A(I5517) );
  INV_X1 NOT_3079( .ZN(g4841), .A(I6531) );
  INV_X4 NOT_3080( .ZN(I8603), .A(g6449) );
  INV_X4 NOT_3081( .ZN(g2361), .A(I3513) );
  INV_X4 NOT_3082( .ZN(I6769), .A(g4786) );
  INV_X1 NOT_3083( .ZN(g4763), .A(I6397) );
  INV_X1 NOT_3084( .ZN(g4191), .A(I5603) );
  INV_X1 NOT_3085( .ZN(g4391), .A(I5876) );
  INV_X1 NOT_3086( .ZN(I5056), .A(g3567) );
  INV_X1 NOT_3087( .ZN(I2986), .A(g1504) );
  INV_X1 NOT_3088( .ZN(I3307), .A(g1339) );
  INV_X1 NOT_3089( .ZN(g1193), .A(I2204) );
  INV_X1 NOT_3090( .ZN(I5529), .A(g3854) );
  INV_X1 NOT_3091( .ZN(I4420), .A(g2096) );
  INV_X1 NOT_3092( .ZN(I5148), .A(g3450) );
  INV_X1 NOT_3093( .ZN(g3136), .A(I4382) );
  INV_X1 NOT_3094( .ZN(g2327), .A(I3481) );
  INV_X1 NOT_3095( .ZN(I6918), .A(g5124) );
  INV_X1 NOT_3096( .ZN(I4507), .A(g2739) );
  INV_X1 NOT_3097( .ZN(g5329), .A(I6989) );
  INV_X2 NOT_3098( .ZN(g1549), .A(g878) );
  INV_X1 NOT_3099( .ZN(g4107), .A(I5403) );
  INV_X1 NOT_3100( .ZN(I7042), .A(g5310) );
  INV_X1 NOT_3101( .ZN(g947), .A(g74) );
  INV_X1 NOT_3102( .ZN(g6894), .A(I9149) );
  INV_X1 NOT_3103( .ZN(g1834), .A(I2916) );
  INV_X1 NOT_3104( .ZN(I4794), .A(g2814) );
  INV_X1 NOT_3105( .ZN(g4307), .A(I5774) );
  INV_X1 NOT_3106( .ZN(I5851), .A(g3739) );
  INV_X1 NOT_3107( .ZN(g4536), .A(I6118) );
  INV_X1 NOT_3108( .ZN(I3858), .A(g2197) );
  INV_X1 NOT_3109( .ZN(I8702), .A(g6572) );
  INV_X1 NOT_3110( .ZN(g2346), .A(I3496) );
  INV_X1 NOT_3111( .ZN(g6735), .A(I8897) );
  INV_X1 NOT_3112( .ZN(I3016), .A(g1754) );
  INV_X1 NOT_3113( .ZN(I2970), .A(g1504) );
  INV_X1 NOT_3114( .ZN(g5727), .A(I7490) );
  INV_X1 NOT_3115( .ZN(I7164), .A(g5433) );
  INV_X1 NOT_3116( .ZN(g2103), .A(I3225) );
  INV_X1 NOT_3117( .ZN(g858), .A(g301) );
  INV_X16 NOT_3118( .ZN(I2925), .A(g1762) );
  INV_X1 NOT_3119( .ZN(g4858), .A(I6582) );
  INV_X1 NOT_3120( .ZN(I3522), .A(g1664) );
  INV_X1 NOT_3121( .ZN(g4016), .A(I5320) );
  INV_X1 NOT_3122( .ZN(I3115), .A(g1519) );
  INV_X1 NOT_3123( .ZN(I3251), .A(g1471) );
  INV_X1 NOT_3124( .ZN(I3811), .A(g2145) );
  INV_X1 NOT_3125( .ZN(I8276), .A(g6303) );
  INV_X1 NOT_3126( .ZN(g1321), .A(I2318) );
  INV_X1 NOT_3127( .ZN(I3047), .A(g1426) );
  INV_X1 NOT_3128( .ZN(g1670), .A(I2648) );
  INV_X1 NOT_3129( .ZN(g3228), .A(I4483) );
  INV_X1 NOT_3130( .ZN(g3465), .A(g2986) );
  INV_X1 NOT_3131( .ZN(g3322), .A(g3070) );
  INV_X1 NOT_3132( .ZN(I5463), .A(g3783) );
  INV_X1 NOT_3133( .ZN(g3230), .A(I4489) );
  INV_X1 NOT_3134( .ZN(g4522), .A(I6078) );
  INV_X1 NOT_3135( .ZN(g4115), .A(I5427) );
  INV_X1 NOT_3136( .ZN(g2753), .A(I3927) );
  INV_X1 NOT_3137( .ZN(g4251), .A(I5705) );
  INV_X1 NOT_3138( .ZN(g1232), .A(I2228) );
  INV_X4 NOT_3139( .ZN(I4300), .A(g2234) );
  INV_X4 NOT_3140( .ZN(g6526), .A(I8494) );
  INV_X1 NOT_3141( .ZN(g1813), .A(I2870) );
  INV_X1 NOT_3142( .ZN(I8527), .A(g6440) );
  INV_X1 NOT_3143( .ZN(I8647), .A(g6528) );
  INV_X1 NOT_3144( .ZN(I2617), .A(g1193) );
  INV_X1 NOT_3145( .ZN(I5720), .A(g4022) );
  INV_X1 NOT_3146( .ZN(g2043), .A(I3158) );
  INV_X1 NOT_3147( .ZN(g6039), .A(g5824) );
  INV_X1 NOT_3148( .ZN(I8764), .A(g6564) );
  INV_X1 NOT_3149( .ZN(g2443), .A(I3578) );
  INV_X1 NOT_3150( .ZN(g6484), .A(g6361) );
  INV_X1 NOT_3151( .ZN(g3096), .A(I4343) );
  INV_X1 NOT_3152( .ZN(g5468), .A(I7150) );
  INV_X1 NOT_3153( .ZN(g1519), .A(I2491) );
  INV_X1 NOT_3154( .ZN(g1740), .A(g1116) );
  INV_X1 NOT_3155( .ZN(I7012), .A(g5316) );
  INV_X1 NOT_3156( .ZN(g6850), .A(I9077) );
  INV_X1 NOT_3157( .ZN(I6895), .A(g5010) );
  INV_X1 NOT_3158( .ZN(I1835), .A(g205) );
  INV_X1 NOT_3159( .ZN(g3845), .A(I5050) );
  INV_X1 NOT_3160( .ZN(I5843), .A(g3851) );
  INV_X1 NOT_3161( .ZN(g2316), .A(I3468) );
  INV_X1 NOT_3162( .ZN(I3537), .A(g1305) );
  INV_X1 NOT_3163( .ZN(I8503), .A(g6434) );
  INV_X1 NOT_3164( .ZN(g1552), .A(g1030) );
  INV_X1 NOT_3165( .ZN(I5457), .A(g3766) );
  INV_X1 NOT_3166( .ZN(g2565), .A(I3675) );
  INV_X1 NOT_3167( .ZN(g6583), .A(I8617) );
  INV_X1 NOT_3168( .ZN(g850), .A(g602) );
  INV_X1 NOT_3169( .ZN(g5576), .A(g5415) );
  INV_X1 NOT_3170( .ZN(g4537), .A(g4410) );
  INV_X1 NOT_3171( .ZN(I7029), .A(g5149) );
  INV_X32 NOT_3172( .ZN(g2347), .A(I3499) );
  INV_X1 NOT_3173( .ZN(I5686), .A(g3942) );
  INV_X1 NOT_3174( .ZN(I4123), .A(g2043) );
  INV_X1 NOT_3175( .ZN(g3807), .A(I5006) );
  INV_X1 NOT_3176( .ZN(g1586), .A(g1052) );
  INV_X1 NOT_3177( .ZN(g3859), .A(I5078) );
  INV_X1 NOT_3178( .ZN(g6276), .A(I7960) );
  INV_X1 NOT_3179( .ZN(g4612), .A(g4320) );
  INV_X1 NOT_3180( .ZN(g2914), .A(g1928) );
  INV_X1 NOT_3181( .ZN(g6616), .A(I8710) );
  INV_X1 NOT_3182( .ZN(I3629), .A(g1759) );
  INV_X1 NOT_3183( .ZN(g6561), .A(I8567) );
  INV_X1 NOT_3184( .ZN(I3328), .A(g1273) );
  INV_X1 NOT_3185( .ZN(I2738), .A(g1236) );
  INV_X1 NOT_3186( .ZN(I8617), .A(g6539) );
  INV_X1 NOT_3187( .ZN(g1341), .A(I2376) );
  INV_X1 NOT_3188( .ZN(g2413), .A(I3553) );
  INV_X1 NOT_3189( .ZN(I4351), .A(g2233) );
  INV_X1 NOT_3190( .ZN(g3342), .A(g3086) );
  INV_X1 NOT_3191( .ZN(g4128), .A(I5466) );
  INV_X1 NOT_3192( .ZN(g1710), .A(g1109) );
  INV_X1 NOT_3193( .ZN(g4629), .A(g4276) );
  INV_X1 NOT_3194( .ZN(I6485), .A(g4603) );
  INV_X1 NOT_3195( .ZN(g6527), .A(I8497) );
  INV_X1 NOT_3196( .ZN(g6404), .A(I8226) );
  INV_X1 NOT_3197( .ZN(g4328), .A(g4092) );
  INV_X1 NOT_3198( .ZN(I2140), .A(g28) );
  INV_X1 NOT_3199( .ZN(g1645), .A(I2614) );
  INV_X1 NOT_3200( .ZN(I2340), .A(g1142) );
  INV_X1 NOT_3201( .ZN(g4130), .A(I5472) );
  INV_X1 NOT_3202( .ZN(I5938), .A(g4351) );
  INV_X1 NOT_3203( .ZN(I7963), .A(g6276) );
  INV_X1 NOT_3204( .ZN(I3800), .A(g2145) );
  INV_X1 NOT_3205( .ZN(g3481), .A(g2612) );
  INV_X1 NOT_3206( .ZN(I2907), .A(g1498) );
  INV_X4 NOT_3207( .ZN(g2820), .A(g2470) );
  INV_X4 NOT_3208( .ZN(g2936), .A(g2026) );
  INV_X1 NOT_3209( .ZN(g5524), .A(I7264) );
  INV_X1 NOT_3210( .ZN(g6503), .A(I8429) );
  INV_X1 NOT_3211( .ZN(g3354), .A(g3096) );
  INV_X1 NOT_3212( .ZN(I4410), .A(g2088) );
  INV_X1 NOT_3213( .ZN(I7808), .A(g5919) );
  INV_X1 NOT_3214( .ZN(g2117), .A(I3244) );
  INV_X1 NOT_3215( .ZN(g3960), .A(I5204) );
  INV_X1 NOT_3216( .ZN(g2317), .A(I3471) );
  INV_X1 NOT_3217( .ZN(g5119), .A(I6769) );
  INV_X1 NOT_3218( .ZN(g6925), .A(I9208) );
  INV_X1 NOT_3219( .ZN(I7707), .A(g5701) );
  INV_X1 NOT_3220( .ZN(I5606), .A(g3821) );
  INV_X1 NOT_3221( .ZN(g1659), .A(I2638) );
  INV_X1 NOT_3222( .ZN(g1358), .A(g1119) );
  INV_X1 NOT_3223( .ZN(g5352), .A(I7002) );
  INV_X1 NOT_3224( .ZN(g5577), .A(g5420) );
  INV_X1 NOT_3225( .ZN(g4213), .A(I5633) );
  INV_X1 NOT_3226( .ZN(g5717), .A(I7478) );
  INV_X1 NOT_3227( .ZN(I3902), .A(g2576) );
  INV_X1 NOT_3228( .ZN(g6120), .A(I7832) );
  INV_X1 NOT_3229( .ZN(g2922), .A(g1960) );
  INV_X1 NOT_3230( .ZN(g1587), .A(g1123) );
  INV_X1 NOT_3231( .ZN(I6812), .A(g5110) );
  INV_X1 NOT_3232( .ZN(I8991), .A(g6788) );
  INV_X16 NOT_3233( .ZN(g3783), .A(I4980) );
  INV_X1 NOT_3234( .ZN(g1111), .A(I2143) );
  INV_X1 NOT_3235( .ZN(I3090), .A(g1504) );
  INV_X1 NOT_3236( .ZN(I9008), .A(g6818) );
  INV_X1 NOT_3237( .ZN(g5893), .A(g5753) );
  INV_X1 NOT_3238( .ZN(g1275), .A(g842) );
  INV_X1 NOT_3239( .ZN(g6277), .A(I7963) );
  INV_X1 NOT_3240( .ZN(g2581), .A(I3694) );
  INV_X1 NOT_3241( .ZN(I3823), .A(g2125) );
  INV_X1 NOT_3242( .ZN(g3267), .A(g3030) );
  INV_X1 NOT_3243( .ZN(I4667), .A(g2908) );
  INV_X1 NOT_3244( .ZN(g3312), .A(I4587) );
  INV_X1 NOT_3245( .ZN(I7865), .A(g6095) );
  INV_X1 NOT_3246( .ZN(I4343), .A(g2525) );
  INV_X1 NOT_3247( .ZN(g2060), .A(g1369) );
  INV_X1 NOT_3248( .ZN(g6617), .A(I8713) );
  INV_X1 NOT_3249( .ZN(g6906), .A(I9185) );
  INV_X1 NOT_3250( .ZN(g5975), .A(g5821) );
  INV_X1 NOT_3251( .ZN(g4512), .A(I6048) );
  INV_X1 NOT_3252( .ZN(I4282), .A(g2525) );
  INV_X1 NOT_3253( .ZN(g2460), .A(I3590) );
  INV_X1 NOT_3254( .ZN(I7604), .A(g5605) );
  INV_X1 NOT_3255( .ZN(I8907), .A(g6702) );
  INV_X1 NOT_3256( .ZN(I3056), .A(g1519) );
  INV_X1 NOT_3257( .ZN(g3001), .A(I4198) );
  INV_X1 NOT_3258( .ZN(g1174), .A(g37) );
  INV_X1 NOT_3259( .ZN(g4823), .A(I6507) );
  INV_X1 NOT_3260( .ZN(I2663), .A(g1006) );
  INV_X1 NOT_3261( .ZN(g4166), .A(I5568) );
  INV_X1 NOT_3262( .ZN(g6516), .A(g6409) );
  INV_X4 NOT_3263( .ZN(g5274), .A(I6933) );
  INV_X4 NOT_3264( .ZN(I8435), .A(g6413) );
  INV_X1 NOT_3265( .ZN(I3148), .A(g1595) );
  INV_X1 NOT_3266( .ZN(I8690), .A(g6571) );
  INV_X1 NOT_3267( .ZN(g1985), .A(I3096) );
  INV_X1 NOT_3268( .ZN(I4334), .A(g2256) );
  INV_X1 NOT_3269( .ZN(I8482), .A(g6461) );
  INV_X1 NOT_3270( .ZN(g2739), .A(I3906) );
  INV_X1 NOT_3271( .ZN(g3761), .A(g3605) );
  INV_X1 NOT_3272( .ZN(I3155), .A(g1612) );
  INV_X1 NOT_3273( .ZN(I3355), .A(g1608) );
  INV_X1 NOT_3274( .ZN(I2402), .A(g774) );
  INV_X1 NOT_3275( .ZN(g4529), .A(I6099) );
  INV_X1 NOT_3276( .ZN(g1284), .A(g851) );
  INV_X1 NOT_3277( .ZN(g4148), .A(I5526) );
  INV_X1 NOT_3278( .ZN(I6733), .A(g4773) );
  INV_X1 NOT_3279( .ZN(I8656), .A(g6532) );
  INV_X1 NOT_3280( .ZN(g3830), .A(I5019) );
  INV_X1 NOT_3281( .ZN(I9122), .A(g6864) );
  INV_X1 NOT_3282( .ZN(g2079), .A(g1348) );
  INV_X1 NOT_3283( .ZN(g4155), .A(I5551) );
  INV_X1 NOT_3284( .ZN(g4851), .A(I6561) );
  INV_X1 NOT_3285( .ZN(g6892), .A(I9143) );
  INV_X1 NOT_3286( .ZN(g1832), .A(I2910) );
  INV_X1 NOT_3287( .ZN(I9230), .A(g6936) );
  INV_X1 NOT_3288( .ZN(g1853), .A(I2955) );
  INV_X1 NOT_3289( .ZN(g2840), .A(g2538) );
  INV_X1 NOT_3290( .ZN(I2877), .A(g1123) );
  INV_X16 NOT_3291( .ZN(I5879), .A(g3745) );
  INV_X1 NOT_3292( .ZN(g5544), .A(g5331) );
  INV_X1 NOT_3293( .ZN(g2390), .A(I3531) );
  INV_X1 NOT_3294( .ZN(I6324), .A(g4450) );
  INV_X1 NOT_3295( .ZN(g1559), .A(g965) );
  INV_X1 NOT_3296( .ZN(I6069), .A(g4213) );
  INV_X1 NOT_3297( .ZN(I8110), .A(g6143) );
  INV_X1 NOT_3298( .ZN(g4463), .A(g4364) );
  INV_X1 NOT_3299( .ZN(g943), .A(g496) );
  INV_X1 NOT_3300( .ZN(g1931), .A(I3034) );
  INV_X1 NOT_3301( .ZN(g6709), .A(I8837) );
  INV_X1 NOT_3302( .ZN(g3932), .A(I5169) );
  INV_X1 NOT_3303( .ZN(I6540), .A(g4714) );
  INV_X1 NOT_3304( .ZN(I3720), .A(g2155) );
  INV_X1 NOT_3305( .ZN(g6078), .A(g5801) );
  INV_X1 NOT_3306( .ZN(I1871), .A(g281) );
  INV_X1 NOT_3307( .ZN(I6377), .A(g4569) );
  INV_X1 NOT_3308( .ZN(g5061), .A(I6701) );
  INV_X1 NOT_3309( .ZN(g6478), .A(I8342) );
  INV_X1 NOT_3310( .ZN(I2464), .A(g850) );
  INV_X1 NOT_3311( .ZN(I3367), .A(g1283) );
  INV_X1 NOT_3312( .ZN(g5387), .A(I7051) );
  INV_X1 NOT_3313( .ZN(I9137), .A(g6864) );
  INV_X1 NOT_3314( .ZN(g1905), .A(I3004) );
  INV_X1 NOT_3315( .ZN(I8002), .A(g6110) );
  INV_X4 NOT_3316( .ZN(g866), .A(g314) );
  INV_X4 NOT_3317( .ZN(I2785), .A(g1222) );
  INV_X1 NOT_3318( .ZN(I7086), .A(g5281) );
  INV_X1 NOT_3319( .ZN(I5615), .A(g3914) );
  INV_X1 NOT_3320( .ZN(g6035), .A(g5824) );
  INV_X1 NOT_3321( .ZN(g4720), .A(I6340) );
  INV_X1 NOT_3322( .ZN(I3843), .A(g2145) );
  INV_X1 NOT_3323( .ZN(g4118), .A(I5436) );
  INV_X1 NOT_3324( .ZN(g4619), .A(g4248) );
  INV_X1 NOT_3325( .ZN(g6517), .A(I8467) );
  INV_X1 NOT_3326( .ZN(g1204), .A(g39) );
  INV_X1 NOT_3327( .ZN(g3677), .A(g3140) );
  INV_X1 NOT_3328( .ZN(g6876), .A(I9095) );
  INV_X1 NOT_3329( .ZN(g4843), .A(I6537) );
  INV_X1 NOT_3330( .ZN(g3866), .A(I5091) );
  INV_X1 NOT_3331( .ZN(g2954), .A(g2381) );
  INV_X1 NOT_3332( .ZN(I4593), .A(g2966) );
  INV_X1 NOT_3333( .ZN(g5046), .A(I6680) );
  INV_X1 NOT_3334( .ZN(g2163), .A(I3288) );
  INV_X1 NOT_3335( .ZN(g6656), .A(I8764) );
  INV_X1 NOT_3336( .ZN(g4193), .A(I5609) );
  INV_X1 NOT_3337( .ZN(I2237), .A(g465) );
  INV_X1 NOT_3338( .ZN(g2032), .A(g1749) );
  INV_X1 NOT_3339( .ZN(g4393), .A(I5882) );
  INV_X1 NOT_3340( .ZN(I5545), .A(g3814) );
  INV_X1 NOT_3341( .ZN(g5403), .A(I7069) );
  INV_X1 NOT_3342( .ZN(I1838), .A(g206) );
  INV_X1 NOT_3343( .ZN(g3848), .A(I5059) );
  INV_X1 NOT_3344( .ZN(I5591), .A(g3821) );
  INV_X1 NOT_3345( .ZN(I4264), .A(g2212) );
  INV_X32 NOT_3346( .ZN(I2394), .A(g719) );
  INV_X1 NOT_3347( .ZN(g5391), .A(I7055) );
  INV_X1 NOT_3348( .ZN(g2568), .A(I3678) );
  INV_X1 NOT_3349( .ZN(I2731), .A(g1117) );
  INV_X1 NOT_3350( .ZN(I4050), .A(g2059) );
  INV_X1 NOT_3351( .ZN(g3241), .A(I4522) );
  INV_X1 NOT_3352( .ZN(g2912), .A(g2001) );
  INV_X1 NOT_3353( .ZN(g4121), .A(I5445) );
  INV_X1 NOT_3354( .ZN(g1969), .A(I3080) );
  INV_X1 NOT_3355( .ZN(I3232), .A(g1782) );
  INV_X1 NOT_3356( .ZN(g4321), .A(I5790) );
  INV_X1 NOT_3357( .ZN(g5307), .A(I6959) );
  INV_X1 NOT_3358( .ZN(g2157), .A(I3278) );
  INV_X1 NOT_3359( .ZN(g5536), .A(g5467) );
  INV_X1 NOT_3360( .ZN(g2357), .A(I3509) );
  INV_X1 NOT_3361( .ZN(g1123), .A(I2165) );
  INV_X1 NOT_3362( .ZN(g1323), .A(I2324) );
  INV_X1 NOT_3363( .ZN(g4625), .A(g4267) );
  INV_X1 NOT_3364( .ZN(I3909), .A(g2044) );
  INV_X1 NOT_3365( .ZN(g4232), .A(I5674) );
  INV_X1 NOT_3366( .ZN(g6402), .A(I8220) );
  INV_X1 NOT_3367( .ZN(g6824), .A(I9005) );
  INV_X1 NOT_3368( .ZN(g1666), .A(g1088) );
  INV_X1 NOT_3369( .ZN(g4938), .A(I6630) );
  INV_X1 NOT_3370( .ZN(I6819), .A(g5019) );
  INV_X1 NOT_3371( .ZN(g6236), .A(g6070) );
  INV_X1 NOT_3372( .ZN(I3519), .A(g1305) );
  INV_X1 NOT_3373( .ZN(I8295), .A(g6295) );
  INV_X1 NOT_3374( .ZN(I2955), .A(g1729) );
  INV_X1 NOT_3375( .ZN(I7487), .A(g5684) );
  INV_X32 NOT_3376( .ZN(g856), .A(g654) );
  INV_X1 NOT_3377( .ZN(I6923), .A(g5124) );
  INV_X1 NOT_3378( .ZN(g1528), .A(g878) );
  INV_X1 NOT_3379( .ZN(I5204), .A(g3534) );
  INV_X1 NOT_3380( .ZN(I5630), .A(g3914) );
  INV_X1 NOT_3381( .ZN(I6488), .A(g4603) );
  INV_X1 NOT_3382( .ZN(g1351), .A(I2388) );
  INV_X1 NOT_3383( .ZN(g1648), .A(I2623) );
  INV_X1 NOT_3384( .ZN(I2814), .A(g1222) );
  INV_X1 NOT_3385( .ZN(g1875), .A(I2970) );
  INV_X1 NOT_3386( .ZN(g4519), .A(I6069) );
  INV_X1 NOT_3387( .ZN(g5115), .A(I6759) );
  INV_X1 NOT_3388( .ZN(g6590), .A(I8638) );
  INV_X1 NOT_3389( .ZN(g5251), .A(g5069) );
  INV_X1 NOT_3390( .ZN(g6877), .A(I9098) );
  INV_X1 NOT_3391( .ZN(g3258), .A(I4537) );
  INV_X1 NOT_3392( .ZN(I4777), .A(g2962) );
  INV_X1 NOT_3393( .ZN(I6701), .A(g4726) );
  INV_X1 NOT_3394( .ZN(g5315), .A(g5116) );
  INV_X1 NOT_3395( .ZN(g3867), .A(I5094) );
  INV_X1 NOT_3396( .ZN(I2150), .A(g10) );
  INV_X1 NOT_3397( .ZN(g1655), .A(g985) );
  INV_X1 NOT_3398( .ZN(g6657), .A(I8767) );
  INV_X1 NOT_3399( .ZN(g4606), .A(g4193) );
  INV_X1 NOT_3400( .ZN(I3687), .A(g1814) );
  INV_X1 NOT_3401( .ZN(I8089), .A(g6120) );
  INV_X1 NOT_3402( .ZN(I2773), .A(g1191) );
  INV_X1 NOT_3403( .ZN(g5874), .A(I7634) );
  INV_X1 NOT_3404( .ZN(g1410), .A(g1233) );
  INV_X1 NOT_3405( .ZN(I8966), .A(g6796) );
  INV_X1 NOT_3406( .ZN(I5750), .A(g4022) );
  INV_X1 NOT_3407( .ZN(I7045), .A(g5167) );
  INV_X1 NOT_3408( .ZN(I6114), .A(g4405) );
  INV_X1 NOT_3409( .ZN(g3975), .A(I5249) );
  INV_X1 NOT_3410( .ZN(I7173), .A(g5436) );
  INV_X32 NOT_3411( .ZN(g1884), .A(I2979) );
  INV_X1 NOT_3412( .ZN(I7091), .A(g5281) );
  INV_X1 NOT_3413( .ZN(g6899), .A(I9164) );
  INV_X1 NOT_3414( .ZN(I4799), .A(g2967) );
  INV_X1 NOT_3415( .ZN(I2212), .A(g123) );
  INV_X1 NOT_3416( .ZN(g929), .A(g49) );
  INV_X1 NOT_3417( .ZN(g6785), .A(I8943) );
  INV_X1 NOT_3418( .ZN(g5880), .A(g5824) );
  INV_X1 NOT_3419( .ZN(I5040), .A(g3271) );
  INV_X1 NOT_3420( .ZN(I2967), .A(g1682) );
  INV_X1 NOT_3421( .ZN(g5537), .A(g5385) );
  INV_X1 NOT_3422( .ZN(g2778), .A(g2391) );
  INV_X1 NOT_3423( .ZN(I1862), .A(g278) );
  INV_X1 NOT_3424( .ZN(I3525), .A(g1461) );
  INV_X1 NOT_3425( .ZN(g3370), .A(g3124) );
  INV_X1 NOT_3426( .ZN(g2894), .A(g1891) );
  INV_X1 NOT_3427( .ZN(I7007), .A(g5314) );
  INV_X1 NOT_3428( .ZN(g1372), .A(I2408) );
  INV_X1 NOT_3429( .ZN(g4141), .A(I5505) );
  INV_X1 NOT_3430( .ZN(g6563), .A(I8573) );
  INV_X1 NOT_3431( .ZN(I6008), .A(g4163) );
  INV_X1 NOT_3432( .ZN(I3691), .A(g1732) );
  INV_X1 NOT_3433( .ZN(g4525), .A(I6087) );
  INV_X1 NOT_3434( .ZN(g1143), .A(I2172) );
  INV_X4 NOT_3435( .ZN(g3984), .A(g3564) );
  INV_X4 NOT_3436( .ZN(I8150), .A(g6185) );
  INV_X1 NOT_3437( .ZN(g1282), .A(g849) );
  INV_X1 NOT_3438( .ZN(I8438), .A(g6416) );
  INV_X1 NOT_3439( .ZN(g3083), .A(I4318) );
  INV_X1 NOT_3440( .ZN(g1988), .A(I3099) );
  INV_X1 NOT_3441( .ZN(I4802), .A(g2877) );
  INV_X1 NOT_3442( .ZN(I6972), .A(g5135) );
  INV_X1 NOT_3443( .ZN(g3483), .A(g2716) );
  INV_X1 NOT_3444( .ZN(I7261), .A(g5458) );
  INV_X1 NOT_3445( .ZN(g6194), .A(I7906) );
  INV_X1 NOT_3446( .ZN(g1334), .A(I2355) );
  INV_X1 NOT_3447( .ZN(I3158), .A(g1829) );
  INV_X1 NOT_3448( .ZN(I3659), .A(g1491) );
  INV_X1 NOT_3449( .ZN(I3358), .A(g1323) );
  INV_X1 NOT_3450( .ZN(g5328), .A(I6986) );
  INV_X1 NOT_3451( .ZN(I1927), .A(g665) );
  INV_X1 NOT_3452( .ZN(g6489), .A(g6369) );
  INV_X1 NOT_3453( .ZN(g5542), .A(g5331) );
  INV_X1 NOT_3454( .ZN(g5330), .A(I6992) );
  INV_X1 NOT_3455( .ZN(g3306), .A(g3057) );
  INV_X1 NOT_3456( .ZN(g2998), .A(I4195) );
  INV_X1 NOT_3457( .ZN(g4158), .A(I5556) );
  INV_X1 NOT_3458( .ZN(g4659), .A(I6250) );
  INV_X1 NOT_3459( .ZN(g1555), .A(I2521) );
  INV_X1 NOT_3460( .ZN(g3790), .A(g3388) );
  INV_X1 NOT_3461( .ZN(I3587), .A(g1461) );
  INV_X1 NOT_3462( .ZN(g1792), .A(I2848) );
  INV_X1 NOT_3463( .ZN(g2603), .A(I3733) );
  INV_X1 NOT_3464( .ZN(g2039), .A(I3148) );
  INV_X4 NOT_3465( .ZN(g3187), .A(I4424) );
  INV_X1 NOT_3466( .ZN(g2484), .A(I3611) );
  INV_X1 NOT_3467( .ZN(g3387), .A(I4664) );
  INV_X1 NOT_3468( .ZN(g3461), .A(g2986) );
  INV_X1 NOT_3469( .ZN(g4587), .A(g4215) );
  INV_X1 NOT_3470( .ZN(I6033), .A(g4179) );
  INV_X1 NOT_3471( .ZN(g5554), .A(g5455) );
  INV_X1 NOT_3472( .ZN(g3622), .A(I4821) );
  INV_X1 NOT_3473( .ZN(g4111), .A(I5415) );
  INV_X1 NOT_3474( .ZN(I8229), .A(g6330) );
  INV_X1 NOT_3475( .ZN(I9149), .A(g6884) );
  INV_X1 NOT_3476( .ZN(I2620), .A(g1177) );
  INV_X1 NOT_3477( .ZN(g1113), .A(I2147) );
  INV_X1 NOT_3478( .ZN(I4492), .A(g3001) );
  INV_X1 NOT_3479( .ZN(g4615), .A(g4322) );
  INV_X1 NOT_3480( .ZN(g2583), .A(g1830) );
  INV_X1 NOT_3481( .ZN(g3904), .A(g3575) );
  INV_X1 NOT_3482( .ZN(g3200), .A(I4437) );
  INV_X1 NOT_3483( .ZN(I6096), .A(g4397) );
  INV_X1 NOT_3484( .ZN(g3046), .A(I4267) );
  INV_X1 NOT_3485( .ZN(g899), .A(I1924) );
  INV_X1 NOT_3486( .ZN(g4374), .A(I5837) );
  INV_X1 NOT_3487( .ZN(I3284), .A(g1702) );
  INV_X1 NOT_3488( .ZN(g2919), .A(g1937) );
  INV_X1 NOT_3489( .ZN(g1908), .A(I3007) );
  INV_X1 NOT_3490( .ZN(I2788), .A(g1236) );
  INV_X1 NOT_3491( .ZN(g1094), .A(I2122) );
  INV_X1 NOT_3492( .ZN(I5618), .A(g3821) );
  INV_X1 NOT_3493( .ZN(g2952), .A(g2381) );
  INV_X1 NOT_3494( .ZN(I6337), .A(g4455) );
  INV_X16 NOT_3495( .ZN(I5343), .A(g3599) );
  INV_X1 NOT_3496( .ZN(g2276), .A(I3425) );
  INV_X1 NOT_3497( .ZN(g1567), .A(I2537) );
  INV_X1 NOT_3498( .ZN(g4284), .A(I5739) );
  INV_X1 NOT_3499( .ZN(g5512), .A(I7254) );
  INV_X1 NOT_3500( .ZN(g4545), .A(g4416) );
  INV_X1 NOT_3501( .ZN(g5090), .A(g4741) );
  INV_X1 NOT_3502( .ZN(g6409), .A(g6285) );
  INV_X1 NOT_3503( .ZN(g5490), .A(I7190) );
  INV_X1 NOT_3504( .ZN(I7689), .A(g5708) );
  INV_X1 NOT_3505( .ZN(g4380), .A(I5851) );
  INV_X1 NOT_3506( .ZN(I2842), .A(g1177) );
  INV_X1 NOT_3507( .ZN(g1776), .A(I2821) );
  INV_X1 NOT_3508( .ZN(g1593), .A(g1054) );
  INV_X1 NOT_3509( .ZN(g2004), .A(I3115) );
  INV_X1 NOT_3510( .ZN(g4853), .A(I6567) );
  INV_X1 NOT_3511( .ZN(g6836), .A(I9031) );
  INV_X1 NOT_3512( .ZN(I2485), .A(g766) );
  INV_X1 NOT_3513( .ZN(I3794), .A(g2044) );
  INV_X1 NOT_3514( .ZN(g2986), .A(g2010) );
  INV_X1 NOT_3515( .ZN(g4020), .A(I5324) );
  INV_X1 NOT_3516( .ZN(g6212), .A(I7910) );
  INV_X1 NOT_3517( .ZN(I5548), .A(g4059) );
  INV_X1 NOT_3518( .ZN(g5456), .A(g5300) );
  INV_X1 NOT_3519( .ZN(g2647), .A(I3791) );
  INV_X1 NOT_3520( .ZN(I8837), .A(g6665) );
  INV_X1 NOT_3521( .ZN(g5148), .A(I6812) );
  INV_X1 NOT_3522( .ZN(g5649), .A(I7404) );
  INV_X16 NOT_3523( .ZN(g4507), .A(I6033) );
  INV_X1 NOT_3524( .ZN(g3223), .A(I4468) );
  INV_X1 NOT_3525( .ZN(I4623), .A(g2962) );
  INV_X1 NOT_3526( .ZN(I1947), .A(g699) );
  INV_X1 NOT_3527( .ZN(g2764), .A(g2357) );
  INV_X1 NOT_3528( .ZN(I8620), .A(g6541) );
  INV_X1 NOT_3529( .ZN(I8462), .A(g6430) );
  INV_X1 NOT_3530( .ZN(I9119), .A(g6855) );
  INV_X1 NOT_3531( .ZN(I2854), .A(g1236) );
  INV_X1 NOT_3532( .ZN(g4559), .A(g4187) );
  INV_X1 NOT_3533( .ZN(g5155), .A(g5099) );
  INV_X1 NOT_3534( .ZN(g5355), .A(I7007) );
  INV_X1 NOT_3535( .ZN(I9152), .A(g6889) );
  INV_X1 NOT_3536( .ZN(g3016), .A(I4223) );
  INV_X1 NOT_3537( .ZN(g6229), .A(g6036) );
  INV_X1 NOT_3538( .ZN(g1160), .A(I2179) );
  INV_X16 NOT_3539( .ZN(g5260), .A(g4938) );
  INV_X1 NOT_3540( .ZN(I6081), .A(g4388) );
  INV_X1 NOT_3541( .ZN(I4375), .A(g2254) );
  INV_X1 NOT_3542( .ZN(g6822), .A(g6786) );
  INV_X1 NOT_3543( .ZN(g1641), .A(I2604) );
  INV_X1 NOT_3544( .ZN(g3251), .A(I4534) );
  INV_X1 NOT_3545( .ZN(I6692), .A(g4720) );
  INV_X1 NOT_3546( .ZN(g1450), .A(I2453) );
  INV_X1 NOT_3547( .ZN(g5063), .A(g4799) );
  INV_X1 NOT_3548( .ZN(I7910), .A(g5905) );
  INV_X1 NOT_3549( .ZN(I8249), .A(g6289) );
  INV_X1 NOT_3550( .ZN(g4628), .A(g4273) );
  INV_X1 NOT_3551( .ZN(g4515), .A(I6057) );
  INV_X1 NOT_3552( .ZN(g2120), .A(I3251) );
  INV_X1 NOT_3553( .ZN(I4285), .A(g2555) );
  INV_X1 NOT_3554( .ZN(g2320), .A(I3474) );
  INV_X1 NOT_3555( .ZN(g4100), .A(I5382) );
  INV_X1 NOT_3556( .ZN(g1724), .A(I2724) );
  INV_X1 NOT_3557( .ZN(g3874), .A(I5103) );
  INV_X1 NOT_3558( .ZN(I2958), .A(g1257) );
  INV_X1 NOT_3559( .ZN(I5094), .A(g3705) );
  INV_X1 NOT_3560( .ZN(I2376), .A(g729) );
  INV_X1 NOT_3561( .ZN(I8485), .A(g6479) );
  INV_X1 NOT_3562( .ZN(g5720), .A(I7481) );
  INV_X1 NOT_3563( .ZN(I2405), .A(g1112) );
  INV_X1 NOT_3564( .ZN(g2906), .A(g1911) );
  INV_X1 NOT_3565( .ZN(g2789), .A(g2410) );
  INV_X1 NOT_3566( .ZN(g1878), .A(I2973) );
  INV_X1 NOT_3567( .ZN(g5118), .A(I6766) );
  INV_X1 NOT_3568( .ZN(I9170), .A(g6883) );
  INV_X16 NOT_3569( .ZN(I1917), .A(g48) );
  AND2_X1 AND2_0( .ZN(g2771), .A1(g2497), .A2(g1975) );
  AND2_X1 AND2_1( .ZN(g6620), .A1(g6516), .A2(g6117) );
  AND2_X1 AND2_2( .ZN(g5193), .A1(g532), .A2(g4967) );
  AND4_X1 AND4_0( .ZN(I5360), .A1(g3532), .A2(g3536), .A3(g3539), .A4(g3544) );
  AND2_X1 AND2_3( .ZN(g5598), .A1(g5046), .A2(g5509) );
  AND2_X1 AND2_4( .ZN(g6249), .A1(g1332), .A2(g5892) );
  AND2_X1 AND2_5( .ZN(g4666), .A1(g4630), .A2(g4627) );
  AND2_X1 AND2_6( .ZN(g3629), .A1(g2809), .A2(g2738) );
  AND2_X2 AND2_7( .ZN(g3328), .A1(g2701), .A2(g1894) );
  AND2_X2 AND2_8( .ZN(g6085), .A1(g1161), .A2(g5731) );
  AND2_X2 AND2_9( .ZN(g4351), .A1(g166), .A2(g3776) );
  AND2_X1 AND2_10( .ZN(g4648), .A1(g4407), .A2(g79) );
  AND2_X1 AND2_11( .ZN(g5232), .A1(g548), .A2(g4980) );
  AND2_X1 AND2_12( .ZN(g2340), .A1(g1398), .A2(g1387) );
  AND2_X1 AND2_13( .ZN(g5938), .A1(g5114), .A2(g5791) );
  AND2_X1 AND2_14( .ZN(g5909), .A1(g5787), .A2(g3384) );
  AND2_X1 AND2_15( .ZN(g1802), .A1(g89), .A2(g1064) );
  AND2_X1 AND2_16( .ZN(g3554), .A1(g2941), .A2(g179) );
  AND2_X1 AND2_17( .ZN(g4410), .A1(g3903), .A2(g1474) );
  AND2_X1 AND2_18( .ZN(g6640), .A1(g1612), .A2(g6549) );
  AND2_X1 AND2_19( .ZN(g4172), .A1(g3930), .A2(g1366) );
  AND2_X1 AND2_20( .ZN(g4372), .A1(g406), .A2(g3790) );
  AND2_X1 AND2_21( .ZN(g3512), .A1(g2928), .A2(g1764) );
  AND2_X1 AND2_22( .ZN(g3490), .A1(g353), .A2(g2959) );
  AND2_X1 AND2_23( .ZN(g4667), .A1(g4653), .A2(g4651) );
  AND2_X1 AND2_24( .ZN(g3166), .A1(g2042), .A2(g1233) );
  AND2_X1 AND2_25( .ZN(g3366), .A1(g248), .A2(g2893) );
  AND2_X1 AND2_26( .ZN(g6829), .A1(g6806), .A2(g5958) );
  AND2_X1 AND2_27( .ZN(g3649), .A1(g3104), .A2(g2764) );
  AND2_X1 AND2_28( .ZN(g6911), .A1(g6904), .A2(g6902) );
  AND2_X1 AND2_29( .ZN(g3155), .A1(g248), .A2(g2461) );
  AND2_X1 AND2_30( .ZN(g3698), .A1(g2284), .A2(g2835) );
  AND2_X1 AND2_31( .ZN(g6270), .A1(g1726), .A2(g6062) );
  AND2_X1 AND2_32( .ZN(g4792), .A1(g1417), .A2(g4471) );
  AND3_X1 AND3_0( .ZN(g6473), .A1(g2036), .A2(g6397), .A3(g1628) );
  AND2_X1 AND2_33( .ZN(g4621), .A1(g3953), .A2(g4364) );
  AND2_X1 AND2_34( .ZN(g5158), .A1(g504), .A2(g4993) );
  AND2_X1 AND2_35( .ZN(g6124), .A1(g5705), .A2(g5958) );
  AND2_X1 AND2_36( .ZN(g6324), .A1(g3880), .A2(g6212) );
  AND3_X1 AND3_1( .ZN(g6469), .A1(g2121), .A2(g2032), .A3(g6394) );
  AND2_X1 AND2_37( .ZN(g3279), .A1(g2599), .A2(g2612) );
  AND2_X1 AND2_38( .ZN(g3619), .A1(g2449), .A2(g3057) );
  AND2_X1 AND2_39( .ZN(g3167), .A1(g1883), .A2(g921) );
  AND2_X1 AND2_40( .ZN(g5311), .A1(g5013), .A2(g4468) );
  AND2_X1 AND2_41( .ZN(g3367), .A1(g2809), .A2(g1960) );
  AND2_X1 AND2_42( .ZN(g3652), .A1(g2544), .A2(g3096) );
  AND3_X1 AND3_2( .ZN(g3843), .A1(g2856), .A2(g945), .A3(g3533) );
  AND2_X1 AND2_43( .ZN(g4593), .A1(g4277), .A2(g947) );
  AND2_X1 AND2_44( .ZN(g3686), .A1(g2256), .A2(g2819) );
  AND2_X1 AND2_45( .ZN(g5180), .A1(g414), .A2(g4950) );
  AND2_X1 AND2_46( .ZN(g5380), .A1(g188), .A2(g5264) );
  AND2_X1 AND2_47( .ZN(g4160), .A1(g3923), .A2(g1345) );
  AND2_X1 AND2_48( .ZN(g3321), .A1(g2252), .A2(g2713) );
  AND2_X2 AND2_49( .ZN(g2089), .A1(g1123), .A2(g1578) );
  AND2_X2 AND2_50( .ZN(g6245), .A1(g1329), .A2(g5889) );
  AND2_X2 AND2_51( .ZN(g4360), .A1(g184), .A2(g3785) );
  AND2_X2 AND2_52( .ZN(g3670), .A1(g2234), .A2(g2792) );
  AND2_X1 AND2_53( .ZN(g3625), .A1(g2619), .A2(g2320) );
  AND2_X1 AND2_54( .ZN(g6291), .A1(g5210), .A2(g6161) );
  AND2_X1 AND2_55( .ZN(g4050), .A1(I5359), .A2(I5360) );
  AND2_X1 AND2_56( .ZN(g5559), .A1(g5024), .A2(g5453) );
  AND2_X1 AND2_57( .ZN(g6144), .A1(g3183), .A2(g5997) );
  AND2_X1 AND2_58( .ZN(g6344), .A1(g6272), .A2(g6080) );
  AND2_X1 AND2_59( .ZN(g2948), .A1(g2137), .A2(g1595) );
  AND2_X1 AND2_60( .ZN(g6259), .A1(g1699), .A2(g6044) );
  AND2_X1 AND2_61( .ZN(g4179), .A1(g390), .A2(g3902) );
  AND2_X1 AND2_62( .ZN(g2955), .A1(g2381), .A2(g297) );
  AND2_X1 AND2_63( .ZN(g6088), .A1(g1143), .A2(g5753) );
  AND2_X1 AND2_64( .ZN(g6852), .A1(g6847), .A2(g2295) );
  AND2_X1 AND2_65( .ZN(g6923), .A1(g6918), .A2(g6917) );
  AND2_X1 AND2_66( .ZN(g5515), .A1(g590), .A2(g5364) );
  AND2_X1 AND2_67( .ZN(g1499), .A1(g1101), .A2(g1094) );
  AND2_X1 AND2_68( .ZN(g4835), .A1(g4533), .A2(g4530) );
  AND2_X1 AND2_69( .ZN(g3687), .A1(g2245), .A2(g2820) );
  AND3_X1 AND3_3( .ZN(g4271), .A1(g2121), .A2(g1749), .A3(g4004) );
  AND3_X1 AND3_4( .ZN(g4611), .A1(g3985), .A2(g119), .A3(g4300) );
  AND2_X1 AND2_70( .ZN(g3341), .A1(g2998), .A2(g2709) );
  AND2_X1 AND2_71( .ZN(g6650), .A1(g6580), .A2(g6235) );
  AND2_X1 AND2_72( .ZN(g4541), .A1(g631), .A2(g4199) );
  AND2_X1 AND2_73( .ZN(g3645), .A1(g2497), .A2(g3090) );
  AND2_X1 AND2_74( .ZN(g5123), .A1(g4670), .A2(g1936) );
  AND2_X1 AND2_75( .ZN(g3691), .A1(g2268), .A2(g2828) );
  AND2_X1 AND2_76( .ZN(g4209), .A1(g3816), .A2(g865) );
  AND2_X1 AND2_77( .ZN(g4353), .A1(g3989), .A2(g3332) );
  AND2_X1 AND2_78( .ZN(g6336), .A1(g6246), .A2(g6065) );
  AND2_X1 AND2_79( .ZN(g6768), .A1(g6750), .A2(g3477) );
  AND2_X1 AND2_80( .ZN(g4744), .A1(g3434), .A2(g4582) );
  AND2_X1 AND2_81( .ZN(g3659), .A1(g2672), .A2(g2361) );
  AND2_X1 AND2_82( .ZN(g5351), .A1(g5326), .A2(g3459) );
  AND2_X1 AND2_83( .ZN(g3358), .A1(g2842), .A2(g1369) );
  AND2_X1 AND2_84( .ZN(g5648), .A1(g4507), .A2(g5545) );
  AND2_X1 AND2_85( .ZN(g6934), .A1(g6932), .A2(g3605) );
  AND2_X1 AND2_86( .ZN(g3275), .A1(g2172), .A2(g2615) );
  AND2_X1 AND2_87( .ZN(g3311), .A1(g218), .A2(g2872) );
  AND2_X1 AND2_88( .ZN(g5410), .A1(g378), .A2(g5274) );
  AND2_X1 AND2_89( .ZN(g3615), .A1(g2422), .A2(g3046) );
  AND2_X1 AND2_90( .ZN(g2062), .A1(g1499), .A2(g1666) );
  AND2_X1 AND2_91( .ZN(g3374), .A1(g2809), .A2(g1969) );
  AND2_X1 AND2_92( .ZN(g4600), .A1(g4054), .A2(g4289) );
  AND2_X1 AND2_93( .ZN(g6096), .A1(g1193), .A2(g5753) );
  AND2_X1 AND2_94( .ZN(g1436), .A1(g834), .A2(g830) );
  AND2_X1 AND2_95( .ZN(g5172), .A1(g441), .A2(g4877) );
  AND2_X1 AND2_96( .ZN(g3180), .A1(g260), .A2(g2506) );
  AND2_X1 AND2_97( .ZN(g5618), .A1(g5506), .A2(g4933) );
  AND2_X1 AND2_98( .ZN(g5143), .A1(g157), .A2(g5099) );
  AND2_X2 AND2_99( .ZN(g6913), .A1(g6900), .A2(g6898) );
  AND2_X2 AND2_100( .ZN(g5235), .A1(g554), .A2(g4980) );
  AND2_X1 AND2_101( .ZN(g4580), .A1(g706), .A2(g4262) );
  AND2_X1 AND2_102( .ZN(g2085), .A1(g1123), .A2(g1567) );
  AND2_X1 AND2_103( .ZN(g6266), .A1(g1721), .A2(g6057) );
  AND2_X1 AND2_104( .ZN(g5555), .A1(g5014), .A2(g5442) );
  AND2_X1 AND2_105( .ZN(g2941), .A1(g2166), .A2(g170) );
  AND2_X1 AND2_106( .ZN(g6248), .A1(g465), .A2(g5894) );
  AND2_X1 AND2_107( .ZN(g6342), .A1(g6264), .A2(g6076) );
  AND2_X1 AND2_108( .ZN(g5621), .A1(g5508), .A2(g4943) );
  AND2_X1 AND2_109( .ZN(g3628), .A1(g2449), .A2(g3070) );
  AND2_X1 AND2_110( .ZN(g6255), .A1(g1335), .A2(g5895) );
  AND2_X1 AND2_111( .ZN(g6081), .A1(g1177), .A2(g5731) );
  AND2_X1 AND2_112( .ZN(g3630), .A1(g3167), .A2(g1756) );
  AND2_X1 AND2_113( .ZN(g6692), .A1(g6616), .A2(g6615) );
  AND2_X1 AND2_114( .ZN(g3300), .A1(g2232), .A2(g2682) );
  AND2_X1 AND2_115( .ZN(g6154), .A1(g3219), .A2(g6015) );
  AND2_X1 AND2_116( .ZN(g6354), .A1(g5866), .A2(g6193) );
  AND2_X1 AND2_117( .ZN(g4184), .A1(g3934), .A2(g2136) );
  AND2_X1 AND2_118( .ZN(g5494), .A1(g5443), .A2(g3455) );
  AND2_X1 AND2_119( .ZN(g4384), .A1(g414), .A2(g3797) );
  AND2_X1 AND2_120( .ZN(g4339), .A1(g3971), .A2(g3289) );
  AND2_X1 AND2_121( .ZN(g4838), .A1(g4648), .A2(g84) );
  AND2_X1 AND2_122( .ZN(g3123), .A1(g230), .A2(g2391) );
  AND2_X1 AND2_123( .ZN(g3323), .A1(g2253), .A2(g2716) );
  AND2_X2 AND2_124( .ZN(g4672), .A1(g4635), .A2(g4631) );
  AND2_X2 AND2_125( .ZN(g2733), .A1(g2422), .A2(g1943) );
  AND2_X1 AND2_126( .ZN(g3666), .A1(g3128), .A2(g2787) );
  AND2_X1 AND2_127( .ZN(g6129), .A1(g5717), .A2(g5975) );
  AND2_X1 AND2_128( .ZN(g6329), .A1(g3888), .A2(g6212) );
  AND2_X1 AND2_129( .ZN(g2073), .A1(g1088), .A2(g1499) );
  AND2_X1 AND2_130( .ZN(g5360), .A1(g4431), .A2(g5160) );
  AND2_X1 AND2_131( .ZN(g6828), .A1(g6803), .A2(g5958) );
  AND2_X1 AND2_132( .ZN(g5050), .A1(g4285), .A2(g4807) );
  AND2_X1 AND2_133( .ZN(g3351), .A1(g2760), .A2(g1931) );
  AND2_X1 AND2_134( .ZN(g6830), .A1(g6809), .A2(g5975) );
  AND2_X1 AND2_135( .ZN(g3648), .A1(g2722), .A2(g2343) );
  AND2_X1 AND2_136( .ZN(g3655), .A1(g2197), .A2(g2768) );
  AND3_X1 AND3_5( .ZN(g1706), .A1(g766), .A2(g719), .A3(g729) );
  AND2_X1 AND2_137( .ZN(g6068), .A1(g5824), .A2(g1726) );
  AND2_X1 AND2_138( .ZN(g4044), .A1(g410), .A2(g3388) );
  AND3_X1 AND3_6( .ZN(g6468), .A1(g2032), .A2(g6394), .A3(g1609) );
  AND2_X1 AND2_139( .ZN(g3172), .A1(g2449), .A2(g2491) );
  AND2_X1 AND2_140( .ZN(g3278), .A1(g2175), .A2(g2628) );
  AND2_X1 AND2_141( .ZN(g3372), .A1(g254), .A2(g2905) );
  AND2_X1 AND2_142( .ZN(g2781), .A1(g2544), .A2(g1982) );
  AND2_X1 AND2_143( .ZN(g3618), .A1(g3016), .A2(g2712) );
  AND2_X2 AND2_144( .ZN(g3667), .A1(g2245), .A2(g2789) );
  AND2_X2 AND2_145( .ZN(g3143), .A1(g242), .A2(g2437) );
  AND2_X1 AND2_146( .ZN(g3282), .A1(g131), .A2(g2863) );
  AND2_X1 AND2_147( .ZN(g6716), .A1(g6682), .A2(g932) );
  AND2_X1 AND2_148( .ZN(g6149), .A1(g3200), .A2(g5997) );
  AND2_X1 AND2_149( .ZN(g3693), .A1(g2256), .A2(g2830) );
  AND2_X1 AND2_150( .ZN(g3134), .A1(g230), .A2(g2413) );
  AND2_X1 AND2_151( .ZN(g3334), .A1(g236), .A2(g2883) );
  AND3_X1 AND3_7( .ZN(g6848), .A1(g3741), .A2(g328), .A3(g6843) );
  AND2_X1 AND2_152( .ZN(g5153), .A1(g492), .A2(g4904) );
  AND2_X1 AND2_153( .ZN(g5209), .A1(g560), .A2(g5025) );
  AND2_X1 AND2_154( .ZN(g5353), .A1(g5327), .A2(g3463) );
  AND2_X1 AND2_155( .ZN(g6241), .A1(g1325), .A2(g5887) );
  AND2_X1 AND2_156( .ZN(g1808), .A1(g706), .A2(g49) );
  AND2_X1 AND2_157( .ZN(g3113), .A1(g224), .A2(g2364) );
  AND2_X1 AND2_158( .ZN(g5558), .A1(g5018), .A2(g5450) );
  AND2_X1 AND2_159( .ZN(g6644), .A1(g6575), .A2(g6230) );
  AND2_X1 AND2_160( .ZN(g6152), .A1(g3212), .A2(g6015) );
  AND2_X1 AND2_161( .ZN(g6258), .A1(g512), .A2(g5899) );
  AND2_X1 AND2_162( .ZN(g4178), .A1(g3959), .A2(g2110) );
  AND2_X1 AND2_163( .ZN(g1575), .A1(g980), .A2(g965) );
  AND2_X1 AND2_164( .ZN(g4378), .A1(g410), .A2(g3792) );
  AND2_X1 AND2_165( .ZN(g4831), .A1(g4528), .A2(g4524) );
  AND2_X1 AND2_166( .ZN(g4182), .A1(g394), .A2(g3904) );
  AND2_X1 AND2_167( .ZN(g5492), .A1(g5441), .A2(g3452) );
  AND2_X1 AND2_168( .ZN(g5600), .A1(g5502), .A2(g4900) );
  AND2_X1 AND2_169( .ZN(g6614), .A1(g932), .A2(g6556) );
  AND2_X1 AND2_170( .ZN(g4947), .A1(g184), .A2(g4741) );
  AND2_X1 AND2_171( .ZN(g3360), .A1(g2783), .A2(g1947) );
  AND2_X2 AND2_172( .ZN(g6125), .A1(g5708), .A2(g5975) );
  AND2_X1 AND2_173( .ZN(g1419), .A1(g613), .A2(g918) );
  AND2_X1 AND2_174( .ZN(g3641), .A1(g2644), .A2(g2333) );
  AND2_X1 AND2_175( .ZN(g4873), .A1(g4838), .A2(g4173) );
  AND2_X1 AND2_176( .ZN(g4037), .A1(g2896), .A2(g3388) );
  AND2_X1 AND2_177( .ZN(g3724), .A1(g117), .A2(g3251) );
  AND2_X1 AND2_178( .ZN(g4495), .A1(g3913), .A2(g4292) );
  AND2_X1 AND2_179( .ZN(g3379), .A1(g3104), .A2(g1988) );
  AND2_X1 AND2_180( .ZN(g5175), .A1(g5094), .A2(g1384) );
  AND2_X1 AND2_181( .ZN(g3658), .A1(g3118), .A2(g2776) );
  AND2_X1 AND2_182( .ZN(g6061), .A1(g5824), .A2(g1711) );
  AND2_X1 AND2_183( .ZN(g5500), .A1(g5430), .A2(g5074) );
  AND2_X1 AND2_184( .ZN(g3611), .A1(g2370), .A2(g3037) );
  AND2_X1 AND2_185( .ZN(g2137), .A1(g760), .A2(g1638) );
  AND2_X1 AND2_186( .ZN(g4042), .A1(g406), .A2(g3388) );
  AND2_X1 AND2_187( .ZN(g5184), .A1(g453), .A2(g4877) );
  AND2_X1 AND2_188( .ZN(g4442), .A1(g4239), .A2(g2882) );
  AND2_X1 AND2_189( .ZN(g4164), .A1(g3958), .A2(g2091) );
  AND2_X1 AND2_190( .ZN(g2807), .A1(g2568), .A2(g2001) );
  AND2_X1 AND2_191( .ZN(g5424), .A1(g390), .A2(g5296) );
  AND2_X1 AND2_192( .ZN(g6145), .A1(g3187), .A2(g6015) );
  AND2_X1 AND2_193( .ZN(g2859), .A1(g2112), .A2(g1649) );
  AND3_X1 AND3_8( .ZN(g3997), .A1(g1250), .A2(g3425), .A3(g2849) );
  AND2_X1 AND2_194( .ZN(g4054), .A1(g3694), .A2(g69) );
  AND2_X1 AND2_195( .ZN(g6345), .A1(g6273), .A2(g6083) );
  AND2_X1 AND2_196( .ZN(g3132), .A1(g2306), .A2(g1206) );
  AND2_X1 AND2_197( .ZN(g3680), .A1(g2245), .A2(g2805) );
  AND2_X1 AND2_198( .ZN(g6637), .A1(g1842), .A2(g6549) );
  AND2_X1 AND2_199( .ZN(g3353), .A1(g3162), .A2(g2921) );
  AND2_X1 AND2_200( .ZN(g2142), .A1(g1793), .A2(g1777) );
  AND2_X1 AND2_201( .ZN(g2255), .A1(g1706), .A2(g736) );
  AND2_X1 AND2_202( .ZN(g6159), .A1(g3177), .A2(g6015) );
  AND2_X2 AND2_203( .ZN(g2081), .A1(g1094), .A2(g1546) );
  AND2_X2 AND2_204( .ZN(g3558), .A1(g338), .A2(g3199) );
  AND2_X1 AND2_205( .ZN(g5499), .A1(g5451), .A2(g3462) );
  AND2_X1 AND2_206( .ZN(g4389), .A1(g449), .A2(g3798) );
  AND2_X1 AND2_207( .ZN(g4171), .A1(g3956), .A2(g2104) );
  AND2_X1 AND2_208( .ZN(g6315), .A1(g3849), .A2(g6194) );
  AND2_X1 AND2_209( .ZN(g4371), .A1(g461), .A2(g3789) );
  AND3_X1 AND3_9( .ZN(g4429), .A1(g923), .A2(g4253), .A3(g2936) );
  AND2_X1 AND2_210( .ZN(g4787), .A1(g2937), .A2(g4628) );
  AND2_X1 AND2_211( .ZN(g6047), .A1(g5824), .A2(g1692) );
  AND2_X1 AND2_212( .ZN(g6874), .A1(g6873), .A2(g2060) );
  AND2_X1 AND2_213( .ZN(g2267), .A1(g1716), .A2(g791) );
  AND3_X1 AND3_10( .ZN(g5444), .A1(g4545), .A2(g5256), .A3(g1574) );
  AND2_X1 AND2_214( .ZN(g5269), .A1(g557), .A2(g5025) );
  AND2_X1 AND2_215( .ZN(g1407), .A1(g301), .A2(g866) );
  AND2_X1 AND2_216( .ZN(g4684), .A1(g4584), .A2(g1341) );
  AND2_X1 AND2_217( .ZN(g4791), .A1(g3936), .A2(g4636) );
  AND2_X1 AND2_218( .ZN(g6243), .A1(g500), .A2(g5890) );
  AND2_X1 AND2_219( .ZN(g6935), .A1(g6933), .A2(g3622) );
  AND2_X1 AND2_220( .ZN(g2746), .A1(g2473), .A2(g1954) );
  AND2_X1 AND2_221( .ZN(g4759), .A1(g536), .A2(g4500) );
  AND2_X1 AND2_222( .ZN(g6128), .A1(g5590), .A2(g5958) );
  AND2_X1 AND2_223( .ZN(g5414), .A1(g382), .A2(g5278) );
  AND2_X1 AND2_224( .ZN(g6130), .A1(g5720), .A2(g5958) );
  AND2_X1 AND2_225( .ZN(g5660), .A1(g4509), .A2(g5549) );
  AND2_X1 AND2_226( .ZN(g3375), .A1(g260), .A2(g2912) );
  AND2_X1 AND2_227( .ZN(g4449), .A1(g4266), .A2(g2887) );
  AND2_X1 AND2_228( .ZN(g3651), .A1(g3064), .A2(g2766) );
  AND2_X1 AND2_229( .ZN(g4865), .A1(g4776), .A2(g1849) );
  AND2_X1 AND2_230( .ZN(g2953), .A1(g2381), .A2(g293) );
  AND2_X2 AND2_231( .ZN(g2068), .A1(g1541), .A2(g1546) );
  AND2_X1 AND2_232( .ZN(g3285), .A1(g2195), .A2(g2653) );
  AND2_X1 AND2_233( .ZN(g4833), .A1(g4521), .A2(g4516) );
  AND2_X1 AND2_234( .ZN(g5178), .A1(g516), .A2(g4993) );
  AND2_X1 AND2_235( .ZN(g5679), .A1(g74), .A2(g5576) );
  AND2_X1 AND2_236( .ZN(g5378), .A1(g179), .A2(g5260) );
  AND2_X1 AND2_237( .ZN(g3339), .A1(g2734), .A2(g1914) );
  AND2_X1 AND2_238( .ZN(g1689), .A1(g766), .A2(g719) );
  AND2_X1 AND2_239( .ZN(g5182), .A1(g520), .A2(g4993) );
  AND2_X1 AND2_240( .ZN(g2699), .A1(g2397), .A2(g1905) );
  AND2_X1 AND2_241( .ZN(g2747), .A1(g2449), .A2(g1957) );
  AND2_X1 AND2_242( .ZN(g6090), .A1(g1161), .A2(g5742) );
  AND2_X1 AND2_243( .ZN(g4362), .A1(g3996), .A2(g3355) );
  AND2_X1 AND2_244( .ZN(g3672), .A1(g3136), .A2(g2800) );
  AND2_X1 AND2_245( .ZN(g4052), .A1(g418), .A2(g3388) );
  AND2_X1 AND2_246( .ZN(g3643), .A1(g2518), .A2(g3086) );
  AND2_X2 AND2_247( .ZN(g4452), .A1(g3820), .A2(g4227) );
  AND2_X2 AND2_248( .ZN(g6056), .A1(g5824), .A2(g1699) );
  AND2_X1 AND2_249( .ZN(g1826), .A1(g714), .A2(g710) );
  AND2_X1 AND2_250( .ZN(g6148), .A1(g3196), .A2(g6015) );
  AND2_X1 AND2_251( .ZN(g6348), .A1(g5869), .A2(g6211) );
  AND2_X1 AND2_252( .ZN(g5560), .A1(g5044), .A2(g5456) );
  AND2_X1 AND2_253( .ZN(g3634), .A1(g2179), .A2(g2744) );
  AND2_X1 AND2_254( .ZN(g6155), .A1(g2588), .A2(g5997) );
  AND2_X1 AND2_255( .ZN(g6851), .A1(g6846), .A2(g2293) );
  AND2_X1 AND2_256( .ZN(g3551), .A1(g2937), .A2(g938) );
  AND2_X1 AND2_257( .ZN(g3099), .A1(g218), .A2(g2350) );
  AND2_X1 AND2_258( .ZN(g3304), .A1(g2857), .A2(g1513) );
  AND2_X1 AND2_259( .ZN(g4486), .A1(g716), .A2(g4195) );
  AND2_X1 AND2_260( .ZN(g3499), .A1(g357), .A2(g2961) );
  AND2_X1 AND2_261( .ZN(g4730), .A1(g1423), .A2(g4565) );
  AND2_X1 AND2_262( .ZN(g5632), .A1(g4494), .A2(g5538) );
  AND2_X1 AND2_263( .ZN(g5095), .A1(g4794), .A2(g951) );
  AND2_X1 AND2_264( .ZN(g6260), .A1(g1703), .A2(g6048) );
  AND2_X1 AND2_265( .ZN(g4185), .A1(g398), .A2(g3906) );
  AND2_X1 AND2_266( .ZN(g1609), .A1(g760), .A2(g754) );
  AND2_X1 AND2_267( .ZN(g5495), .A1(g5444), .A2(g3456) );
  AND4_X1 AND4_1( .ZN(g2577), .A1(g1743), .A2(g1797), .A3(g1793), .A4(g1138) );
  AND2_X1 AND2_268( .ZN(g3613), .A1(g2604), .A2(g2312) );
  AND2_X1 AND2_269( .ZN(g6619), .A1(g6515), .A2(g6115) );
  AND2_X1 AND2_270( .ZN(g6318), .A1(g3865), .A2(g6212) );
  AND4_X1 AND4_2( .ZN(g2026), .A1(g1359), .A2(g1402), .A3(g1398), .A4(g901) );
  AND2_X1 AND2_271( .ZN(g5164), .A1(g437), .A2(g4877) );
  AND2_X1 AND2_272( .ZN(g5364), .A1(g574), .A2(g5194) );
  AND2_X1 AND2_273( .ZN(g5233), .A1(g551), .A2(g4980) );
  AND2_X1 AND2_274( .ZN(g2821), .A1(g1890), .A2(g910) );
  AND2_X1 AND2_275( .ZN(g3729), .A1(g327), .A2(g3441) );
  AND2_X1 AND2_276( .ZN(g5454), .A1(g5256), .A2(g4549) );
  AND2_X1 AND2_277( .ZN(g5553), .A1(g5012), .A2(g5440) );
  AND2_X1 AND2_278( .ZN(g6321), .A1(g3873), .A2(g6212) );
  AND2_X1 AND2_279( .ZN(g3660), .A1(g2568), .A2(g3110) );
  AND3_X1 AND3_11( .ZN(g6625), .A1(g2121), .A2(g1595), .A3(g6538) );
  AND2_X1 AND2_280( .ZN(g4045), .A1(g3425), .A2(g123) );
  AND2_X1 AND2_281( .ZN(g4445), .A1(g4235), .A2(g1854) );
  AND2_X2 AND2_282( .ZN(g6253), .A1(g508), .A2(g5896) );
  AND2_X1 AND2_283( .ZN(g4373), .A1(g4001), .A2(g3370) );
  AND2_X1 AND2_284( .ZN(g5189), .A1(g528), .A2(g4993) );
  AND2_X1 AND2_285( .ZN(g4491), .A1(g3554), .A2(g4215) );
  AND2_X1 AND2_286( .ZN(g6909), .A1(g6896), .A2(g6894) );
  AND2_X1 AND2_287( .ZN(g4169), .A1(g3966), .A2(g2099) );
  AND2_X1 AND2_288( .ZN(g5171), .A1(g406), .A2(g4950) );
  AND2_X1 AND2_289( .ZN(g4369), .A1(g3999), .A2(g3364) );
  AND2_X1 AND2_290( .ZN(g3679), .A1(g2245), .A2(g2803) );
  AND2_X1 AND2_291( .ZN(g4602), .A1(g4407), .A2(g4293) );
  AND2_X1 AND2_292( .ZN(g5371), .A1(g152), .A2(g5248) );
  AND2_X1 AND2_293( .ZN(g3378), .A1(g3136), .A2(g2932) );
  AND2_X1 AND2_294( .ZN(g5429), .A1(g398), .A2(g5304) );
  AND2_X1 AND2_295( .ZN(g4407), .A1(g4054), .A2(g74) );
  AND2_X1 AND2_296( .ZN(g5956), .A1(g5783), .A2(g5425) );
  AND2_X1 AND2_297( .ZN(g4868), .A1(g4774), .A2(g2891) );
  AND2_X1 AND2_298( .ZN(g5675), .A1(g64), .A2(g5574) );
  AND2_X1 AND2_299( .ZN(g3135), .A1(g2370), .A2(g2416) );
  AND2_X1 AND2_300( .ZN(g4459), .A1(g4245), .A2(g1899) );
  AND2_X1 AND2_301( .ZN(g3335), .A1(g230), .A2(g2884) );
  AND2_X1 AND2_302( .ZN(g3831), .A1(g2330), .A2(g3425) );
  AND2_X1 AND2_303( .ZN(g3182), .A1(g2473), .A2(g2512) );
  AND2_X2 AND2_304( .ZN(g3288), .A1(g2631), .A2(g2634) );
  AND2_X2 AND2_305( .ZN(g3382), .A1(g3136), .A2(g2934) );
  AND2_X1 AND2_306( .ZN(g4793), .A1(g4277), .A2(g4639) );
  AND2_X1 AND2_307( .ZN(g4015), .A1(g445), .A2(g3388) );
  AND2_X1 AND2_308( .ZN(g2107), .A1(g1583), .A2(g1543) );
  AND2_X1 AND2_309( .ZN(g6141), .A1(g3173), .A2(g5997) );
  AND2_X1 AND2_310( .ZN(g6341), .A1(g6261), .A2(g6074) );
  AND2_X1 AND2_311( .ZN(g6645), .A1(g6576), .A2(g6231) );
  AND2_X1 AND2_312( .ZN(g3632), .A1(g3043), .A2(g2743) );
  AND2_X1 AND2_313( .ZN(g3437), .A1(g837), .A2(g2853) );
  AND2_X1 AND2_314( .ZN(g3653), .A1(g2215), .A2(g2767) );
  AND2_X1 AND2_315( .ZN(g5201), .A1(g4859), .A2(g5084) );
  AND2_X1 AND2_316( .ZN(g3208), .A1(g895), .A2(g2551) );
  AND2_X1 AND2_317( .ZN(g3302), .A1(g212), .A2(g2867) );
  AND2_X1 AND2_318( .ZN(g6158), .A1(g2594), .A2(g6015) );
  AND2_X1 AND2_319( .ZN(g5449), .A1(g4545), .A2(g5246) );
  AND2_X1 AND2_320( .ZN(g5604), .A1(g5059), .A2(g5521) );
  AND2_X1 AND2_321( .ZN(g5098), .A1(g4021), .A2(g4837) );
  AND2_X1 AND2_322( .ZN(g5498), .A1(g5449), .A2(g3460) );
  AND2_X1 AND2_323( .ZN(g1585), .A1(g1017), .A2(g1011) );
  AND2_X1 AND2_324( .ZN(g6275), .A1(g1735), .A2(g6070) );
  AND2_X1 AND2_325( .ZN(g6311), .A1(g3837), .A2(g6194) );
  AND2_X1 AND2_326( .ZN(g4671), .A1(g4645), .A2(g4641) );
  AND3_X1 AND3_12( .ZN(g4247), .A1(g1764), .A2(g4007), .A3(g1628) );
  AND2_X1 AND2_327( .ZN(g3454), .A1(g2933), .A2(g1660) );
  AND2_X1 AND2_328( .ZN(g4826), .A1(g4209), .A2(g4463) );
  AND2_X1 AND2_329( .ZN(g5162), .A1(g5088), .A2(g2105) );
  AND2_X1 AND2_330( .ZN(g5362), .A1(g4437), .A2(g5174) );
  AND2_X1 AND2_331( .ZN(g3296), .A1(g3054), .A2(g2650) );
  AND2_X1 AND2_332( .ZN(g5419), .A1(g386), .A2(g5292) );
  AND2_X1 AND2_333( .ZN(g3725), .A1(g118), .A2(g3251) );
  AND2_X1 AND2_334( .ZN(g2935), .A1(g2291), .A2(g1788) );
  AND2_X1 AND2_335( .ZN(g5452), .A1(g5315), .A2(g4612) );
  AND2_X1 AND2_336( .ZN(g6559), .A1(g1612), .A2(g6474) );
  AND2_X1 AND2_337( .ZN(g5728), .A1(g5623), .A2(g3889) );
  AND2_X2 AND2_338( .ZN(g5486), .A1(g386), .A2(g5331) );
  AND2_X2 AND2_339( .ZN(g5185), .A1(g524), .A2(g4993) );
  AND2_X1 AND2_340( .ZN(g3171), .A1(g248), .A2(g2488) );
  AND2_X1 AND2_341( .ZN(g3371), .A1(g260), .A2(g2904) );
  AND3_X1 AND3_13( .ZN(g6628), .A1(g2138), .A2(g1612), .A3(g6540) );
  AND2_X1 AND2_342( .ZN(g4165), .A1(g3927), .A2(g1352) );
  AND2_X1 AND2_343( .ZN(g4048), .A1(g414), .A2(g3388) );
  AND2_X1 AND2_344( .ZN(g4448), .A1(g3815), .A2(g4225) );
  AND2_X1 AND2_345( .ZN(g3281), .A1(g2178), .A2(g2640) );
  AND2_X1 AND2_346( .ZN(g4827), .A1(g4520), .A2(g4515) );
  AND2_X1 AND2_347( .ZN(g4333), .A1(g3964), .A2(g3284) );
  AND3_X1 AND3_14( .ZN(I2566), .A1(g749), .A2(g743), .A3(g736) );
  AND2_X1 AND2_348( .ZN(g2166), .A1(g1633), .A2(g161) );
  AND2_X1 AND2_349( .ZN(g3684), .A1(g2268), .A2(g2817) );
  AND2_X1 AND2_350( .ZN(g4396), .A1(g422), .A2(g3801) );
  AND2_X1 AND2_351( .ZN(g3338), .A1(g3162), .A2(g2914) );
  AND2_X1 AND2_352( .ZN(g2056), .A1(g1672), .A2(g1675) );
  AND2_X2 AND2_353( .ZN(g5406), .A1(g374), .A2(g5270) );
  AND2_X2 AND2_354( .ZN(g3309), .A1(g2243), .A2(g2695) );
  AND2_X2 AND2_355( .ZN(g5635), .A1(g4498), .A2(g5542) );
  AND2_X2 AND2_356( .ZN(g5682), .A1(g84), .A2(g5578) );
  AND2_X2 AND2_357( .ZN(g5487), .A1(g390), .A2(g5331) );
  AND2_X2 AND2_358( .ZN(g6123), .A1(g5702), .A2(g5958) );
  AND2_X1 AND2_359( .ZN(g6323), .A1(g3877), .A2(g6194) );
  AND2_X1 AND2_360( .ZN(g3759), .A1(g2644), .A2(g3498) );
  AND2_X1 AND2_361( .ZN(g5226), .A1(g672), .A2(g5054) );
  AND2_X1 AND2_362( .ZN(g6151), .A1(g3209), .A2(g5997) );
  AND2_X1 AND2_363( .ZN(g3449), .A1(g128), .A2(g2946) );
  AND2_X1 AND2_364( .ZN(g6648), .A1(g6579), .A2(g6234) );
  AND2_X1 AND2_365( .ZN(g5173), .A1(g512), .A2(g4993) );
  AND2_X1 AND2_366( .ZN(g5373), .A1(g161), .A2(g5250) );
  AND2_X1 AND2_367( .ZN(g4181), .A1(g3939), .A2(g1381) );
  AND2_X1 AND2_368( .ZN(g2720), .A1(g2422), .A2(g1919) );
  AND2_X1 AND2_369( .ZN(g4685), .A1(g4591), .A2(g2079) );
  AND2_X1 AND2_370( .ZN(g5169), .A1(g5093), .A2(g1375) );
  AND2_X1 AND2_371( .ZN(g5369), .A1(g143), .A2(g5247) );
  AND2_X1 AND2_372( .ZN(g5602), .A1(g594), .A2(g5515) );
  AND4_X1 AND4_3( .ZN(g2834), .A1(g1263), .A2(g1257), .A3(g1270), .A4(I4040) );
  AND2_X1 AND2_373( .ZN(g3362), .A1(g3031), .A2(g2740) );
  AND2_X1 AND2_374( .ZN(g6343), .A1(g6268), .A2(g6078) );
  AND2_X1 AND2_375( .ZN(g2121), .A1(g1632), .A2(g754) );
  AND2_X1 AND2_376( .ZN(g2670), .A1(g2029), .A2(g1503) );
  AND2_X1 AND2_377( .ZN(g6693), .A1(g6618), .A2(g6617) );
  AND2_X1 AND2_378( .ZN(g1633), .A1(g716), .A2(g152) );
  AND2_X1 AND2_379( .ZN(g6334), .A1(g3858), .A2(g6212) );
  AND2_X1 AND2_380( .ZN(g3728), .A1(g326), .A2(g3441) );
  AND2_X1 AND2_381( .ZN(g6555), .A1(g1838), .A2(g6469) );
  AND2_X1 AND2_382( .ZN(g3730), .A1(g328), .A2(g3441) );
  AND2_X1 AND2_383( .ZN(g2909), .A1(g606), .A2(g2092) );
  AND2_X1 AND2_384( .ZN(g4041), .A1(g461), .A2(g3388) );
  AND2_X1 AND2_385( .ZN(g3425), .A1(g2296), .A2(g3208) );
  AND2_X1 AND2_386( .ZN(g6313), .A1(g3841), .A2(g6194) );
  AND2_X1 AND2_387( .ZN(g5940), .A1(g5115), .A2(g5794) );
  AND2_X2 AND2_388( .ZN(g4673), .A1(g4656), .A2(g4654) );
  AND2_X2 AND2_389( .ZN(g5188), .A1(g1043), .A2(g4894) );
  AND2_X1 AND2_390( .ZN(g6908), .A1(g6907), .A2(g3886) );
  AND2_X1 AND2_391( .ZN(g5216), .A1(g563), .A2(g5025) );
  AND2_X1 AND2_392( .ZN(g6094), .A1(g1177), .A2(g5753) );
  AND2_X1 AND2_393( .ZN(g4168), .A1(g3925), .A2(g1355) );
  AND2_X1 AND2_394( .ZN(g4368), .A1(g3998), .A2(g3363) );
  AND2_X1 AND2_395( .ZN(g5671), .A1(g54), .A2(g5572) );
  AND2_X1 AND2_396( .ZN(g3678), .A1(g2256), .A2(g2802) );
  AND2_X1 AND2_397( .ZN(g5428), .A1(g394), .A2(g5300) );
  AND2_X1 AND2_398( .ZN(g4058), .A1(g3424), .A2(g1246) );
  AND2_X1 AND2_399( .ZN(g3635), .A1(g2473), .A2(g3079) );
  AND2_X1 AND2_400( .ZN(g2860), .A1(g710), .A2(g2296) );
  AND2_X1 AND2_401( .ZN(g3682), .A1(g2772), .A2(g2430) );
  AND2_X1 AND2_402( .ZN(g3305), .A1(g2960), .A2(g2296) );
  AND2_X1 AND2_403( .ZN(g5910), .A1(g5816), .A2(g5667) );
  AND2_X1 AND2_404( .ZN(g3755), .A1(g2604), .A2(g3481) );
  AND2_X1 AND2_405( .ZN(g2659), .A1(g1686), .A2(g2296) );
  AND2_X1 AND2_406( .ZN(g5883), .A1(g5824), .A2(g3752) );
  AND2_X1 AND2_407( .ZN(g3373), .A1(g3118), .A2(g2927) );
  AND2_X1 AND2_408( .ZN(g5217), .A1(g4866), .A2(g5092) );
  AND2_X1 AND2_409( .ZN(g4863), .A1(g4777), .A2(g2874) );
  AND2_X1 AND2_410( .ZN(g3283), .A1(g2609), .A2(g2622) );
  AND2_X1 AND2_411( .ZN(g3602), .A1(g2688), .A2(g2663) );
  AND3_X1 AND3_15( .ZN(I2574), .A1(g804), .A2(g798), .A3(g791) );
  AND2_X1 AND2_412( .ZN(g5165), .A1(g508), .A2(g4993) );
  AND2_X1 AND2_413( .ZN(g6777), .A1(g6762), .A2(g3488) );
  AND3_X1 AND3_16( .ZN(g3718), .A1(g1743), .A2(g3140), .A3(g1157) );
  AND2_X1 AND2_414( .ZN(g3767), .A1(g2706), .A2(g3504) );
  AND2_X1 AND2_415( .ZN(g4688), .A1(g1474), .A2(g4568) );
  AND2_X1 AND2_416( .ZN(g1784), .A1(g858), .A2(g889) );
  AND2_X1 AND2_417( .ZN(g2853), .A1(g836), .A2(g2021) );
  AND2_X1 AND2_418( .ZN(g6799), .A1(g4948), .A2(g6782) );
  AND2_X1 AND2_419( .ZN(g2794), .A1(g2544), .A2(g1994) );
  AND2_X1 AND2_420( .ZN(g3203), .A1(g2497), .A2(g2565) );
  AND2_X1 AND2_421( .ZN(g6132), .A1(g3752), .A2(g5880) );
  AND2_X1 AND2_422( .ZN(g6238), .A1(g528), .A2(g5886) );
  AND2_X1 AND2_423( .ZN(g6153), .A1(g3216), .A2(g5997) );
  AND2_X1 AND2_424( .ZN(g4183), .A1(g3965), .A2(g1391) );
  AND2_X1 AND2_425( .ZN(g4383), .A1(g453), .A2(g3796) );
  AND2_X1 AND2_426( .ZN(g6558), .A1(g1842), .A2(g6474) );
  AND2_X1 AND2_427( .ZN(g5181), .A1(g449), .A2(g4877) );
  AND2_X1 AND2_428( .ZN(g3689), .A1(g3162), .A2(g2826) );
  AND2_X2 AND2_429( .ZN(g4588), .A1(g2419), .A2(g4273) );
  AND2_X2 AND2_430( .ZN(g5197), .A1(g465), .A2(g4967) );
  AND2_X1 AND2_431( .ZN(g4161), .A1(g3931), .A2(g2087) );
  AND2_X1 AND2_432( .ZN(g4361), .A1(g3995), .A2(g3354) );
  AND2_X1 AND2_433( .ZN(g3671), .A1(g2760), .A2(g2405) );
  AND2_X1 AND2_434( .ZN(g4051), .A1(g449), .A2(g3388) );
  AND2_X1 AND2_435( .ZN(g6092), .A1(g1123), .A2(g5731) );
  AND2_X1 AND2_436( .ZN(g4346), .A1(g157), .A2(g3773) );
  AND2_X1 AND2_437( .ZN(g2323), .A1(g471), .A2(g1358) );
  AND2_X1 AND2_438( .ZN(g5562), .A1(g5228), .A2(g5457) );
  AND2_X1 AND2_439( .ZN(g3910), .A1(g3546), .A2(g1049) );
  AND2_X1 AND2_440( .ZN(g3609), .A1(g2706), .A2(g2678) );
  AND2_X1 AND2_441( .ZN(g6262), .A1(g516), .A2(g5901) );
  AND3_X1 AND3_17( .ZN(g6736), .A1(g6712), .A2(g754), .A3(g5237) );
  AND2_X1 AND2_442( .ZN(g3758), .A1(g545), .A2(g3461) );
  AND2_X1 AND2_443( .ZN(g4043), .A1(g457), .A2(g3388) );
  AND2_X1 AND2_444( .ZN(g3365), .A1(g254), .A2(g2892) );
  AND3_X1 AND3_18( .ZN(g5441), .A1(g4537), .A2(g5251), .A3(g1558) );
  AND2_X1 AND2_445( .ZN(g5673), .A1(g59), .A2(g5573) );
  AND2_X1 AND2_446( .ZN(g4347), .A1(g3986), .A2(g3320) );
  AND2_X1 AND2_447( .ZN(g3133), .A1(g236), .A2(g2410) );
  AND2_X1 AND2_448( .ZN(g3333), .A1(g2264), .A2(g2728) );
  AND2_X1 AND2_449( .ZN(g3774), .A1(g3016), .A2(g3510) );
  AND2_X1 AND2_450( .ZN(g4697), .A1(g4589), .A2(g1363) );
  AND2_X1 AND2_451( .ZN(g3780), .A1(g3043), .A2(g3519) );
  AND3_X1 AND3_19( .ZN(g6737), .A1(g6714), .A2(g760), .A3(g5237) );
  AND2_X1 AND2_452( .ZN(g6077), .A1(g5824), .A2(g1735) );
  AND2_X1 AND2_453( .ZN(g3662), .A1(g2544), .A2(g3114) );
  AND2_X1 AND2_454( .ZN(g6643), .A1(g6574), .A2(g6229) );
  AND2_X1 AND2_455( .ZN(g3290), .A1(g2213), .A2(g2664) );
  AND2_X1 AND2_456( .ZN(g6634), .A1(g1595), .A2(g6545) );
  AND2_X1 AND2_457( .ZN(g3816), .A1(g3434), .A2(g861) );
  AND2_X1 AND2_458( .ZN(g2113), .A1(g1576), .A2(g1535) );
  AND2_X1 AND2_459( .ZN(g6099), .A1(g1222), .A2(g5753) );
  AND2_X1 AND2_460( .ZN(g6304), .A1(g5915), .A2(g6165) );
  AND2_X1 AND2_461( .ZN(g3181), .A1(g254), .A2(g2509) );
  AND2_X1 AND2_462( .ZN(g3381), .A1(g3128), .A2(g1998) );
  AND2_X1 AND2_463( .ZN(g3685), .A1(g2256), .A2(g2818) );
  AND2_X1 AND2_464( .ZN(g3700), .A1(g2276), .A2(g2837) );
  AND2_X1 AND2_465( .ZN(g3421), .A1(g622), .A2(g2846) );
  AND2_X1 AND2_466( .ZN(g5569), .A1(g5348), .A2(g3772) );
  AND2_X1 AND2_467( .ZN(g4460), .A1(g4218), .A2(g1539) );
  AND2_X1 AND2_468( .ZN(g4597), .A1(g3694), .A2(g4286) );
  AND2_X2 AND2_469( .ZN(g6613), .A1(g932), .A2(g6554) );
  AND2_X1 AND2_470( .ZN(g4739), .A1(g2850), .A2(g4579) );
  AND2_X1 AND2_471( .ZN(g6269), .A1(g524), .A2(g5908) );
  AND2_X1 AND2_472( .ZN(g4937), .A1(g166), .A2(g4732) );
  AND2_X1 AND2_473( .ZN(g4668), .A1(g4642), .A2(g4638) );
  AND2_X1 AND2_474( .ZN(g3631), .A1(g2631), .A2(g2324) );
  AND2_X1 AND2_475( .ZN(g2160), .A1(g1624), .A2(g929) );
  AND2_X1 AND2_476( .ZN(g4390), .A1(g418), .A2(g3799) );
  AND2_X1 AND2_477( .ZN(g3301), .A1(g218), .A2(g2866) );
  AND2_X1 AND2_478( .ZN(g4501), .A1(g4250), .A2(g1671) );
  AND2_X1 AND2_479( .ZN(g4156), .A1(g3926), .A2(g2078) );
  AND2_X1 AND2_480( .ZN(g4356), .A1(g175), .A2(g3779) );
  AND2_X1 AND2_481( .ZN(g4942), .A1(g175), .A2(g4736) );
  AND2_X1 AND2_482( .ZN(g5183), .A1(g418), .A2(g4950) );
  AND2_X1 AND2_483( .ZN(g4163), .A1(g374), .A2(g3892) );
  AND2_X1 AND2_484( .ZN(g5023), .A1(g3935), .A2(g4804) );
  AND2_X1 AND2_485( .ZN(g4363), .A1(g402), .A2(g3786) );
  AND2_X1 AND2_486( .ZN(g4032), .A1(g441), .A2(g3388) );
  AND2_X1 AND2_487( .ZN(g4053), .A1(g3387), .A2(g1415) );
  AND2_X1 AND2_488( .ZN(g4453), .A1(g4238), .A2(g1858) );
  AND2_X1 AND2_489( .ZN(g5161), .A1(g5095), .A2(g4535) );
  AND2_X1 AND2_490( .ZN(g3669), .A1(g2234), .A2(g2790) );
  AND2_X1 AND2_491( .ZN(g5361), .A1(g4435), .A2(g5168) );
  AND2_X1 AND2_492( .ZN(g3368), .A1(g2822), .A2(g2923) );
  AND2_X1 AND2_493( .ZN(g6135), .A1(g5584), .A2(g5958) );
  AND2_X1 AND2_494( .ZN(g5665), .A1(g361), .A2(g5570) );
  AND2_X1 AND2_495( .ZN(g6831), .A1(g6812), .A2(g5975) );
  AND2_X1 AND2_496( .ZN(g5451), .A1(g5251), .A2(g4544) );
  AND2_X1 AND2_497( .ZN(g6288), .A1(g5615), .A2(g6160) );
  AND2_X1 AND2_498( .ZN(g4157), .A1(g3830), .A2(g1533) );
  AND2_X1 AND2_499( .ZN(g4357), .A1(g3990), .A2(g3342) );
  AND2_X1 AND2_500( .ZN(g5146), .A1(g184), .A2(g5099) );
  AND2_X1 AND2_501( .ZN(g6916), .A1(g6903), .A2(g6901) );
  AND2_X1 AND2_502( .ZN(g5633), .A1(g4496), .A2(g5539) );
  AND2_X1 AND2_503( .ZN(g3505), .A1(g2924), .A2(g1749) );
  AND2_X1 AND2_504( .ZN(g6749), .A1(g6735), .A2(g6734) );
  AND2_X2 AND2_505( .ZN(g6798), .A1(g4946), .A2(g6781) );
  AND2_X2 AND2_506( .ZN(g5944), .A1(g5778), .A2(g5403) );
  AND2_X1 AND2_507( .ZN(g5240), .A1(g293), .A2(g4915) );
  AND2_X1 AND2_508( .ZN(g5043), .A1(g3941), .A2(g4805) );
  AND3_X1 AND3_20( .ZN(g5443), .A1(g4537), .A2(g5251), .A3(g2307) );
  AND2_X1 AND2_509( .ZN(g6302), .A1(g5740), .A2(g6164) );
  AND2_X1 AND2_510( .ZN(g6719), .A1(g4518), .A2(g6665) );
  AND2_X1 AND2_511( .ZN(g2092), .A1(g642), .A2(g1570) );
  AND2_X1 AND2_512( .ZN(g4683), .A1(g4585), .A2(g2066) );
  AND2_X1 AND2_513( .ZN(g5681), .A1(g79), .A2(g5577) );
  AND2_X1 AND2_514( .ZN(g3688), .A1(g2783), .A2(g2457) );
  AND2_X1 AND2_515( .ZN(g4735), .A1(g2018), .A2(g4577) );
  AND2_X1 AND2_516( .ZN(g6265), .A1(g520), .A2(g5903) );
  AND2_X1 AND2_517( .ZN(g4782), .A1(g1624), .A2(g4623) );
  AND2_X1 AND2_518( .ZN(g4661), .A1(g4637), .A2(g4634) );
  AND2_X1 AND2_519( .ZN(g4949), .A1(g193), .A2(g4753) );
  AND2_X1 AND2_520( .ZN(g3326), .A1(g2734), .A2(g1891) );
  AND2_X1 AND2_521( .ZN(g6770), .A1(g6754), .A2(g3482) );
  AND2_X1 AND2_522( .ZN(g3760), .A1(g548), .A2(g3465) );
  AND2_X2 AND2_523( .ZN(g5936), .A1(g5113), .A2(g5788) );
  AND2_X2 AND2_524( .ZN(g4039), .A1(g402), .A2(g3388) );
  AND2_X1 AND2_525( .ZN(g5317), .A1(g148), .A2(g4869) );
  AND2_X1 AND2_526( .ZN(g3383), .A1(g3128), .A2(g2004) );
  AND2_X1 AND2_527( .ZN(g5601), .A1(g5052), .A2(g5518) );
  AND2_X1 AND2_528( .ZN(g3608), .A1(g2599), .A2(g2308) );
  AND2_X1 AND2_529( .ZN(g3924), .A1(g3505), .A2(g471) );
  AND2_X1 AND2_530( .ZN(g4583), .A1(g1808), .A2(g4267) );
  AND2_X1 AND2_531( .ZN(g3161), .A1(g2397), .A2(g2470) );
  AND2_X1 AND2_532( .ZN(g2339), .A1(g1603), .A2(g197) );
  AND2_X1 AND2_533( .ZN(g3361), .A1(g3150), .A2(g1950) );
  AND2_X1 AND2_534( .ZN(g4616), .A1(g4231), .A2(g3761) );
  AND2_X1 AND2_535( .ZN(g3665), .A1(g2748), .A2(g2378) );
  AND2_X1 AND2_536( .ZN(g3127), .A1(g224), .A2(g2394) );
  AND2_X1 AND2_537( .ZN(g3327), .A1(g2772), .A2(g2906) );
  AND2_X1 AND2_538( .ZN(g3146), .A1(g2370), .A2(g2446) );
  AND2_X1 AND2_539( .ZN(g3633), .A1(g2497), .A2(g3076) );
  AND2_X1 AND2_540( .ZN(g5937), .A1(g5775), .A2(g5392) );
  AND2_X1 AND2_541( .ZN(g3103), .A1(g212), .A2(g2353) );
  AND2_X1 AND2_542( .ZN(g3303), .A1(g2722), .A2(g2890) );
  AND2_X1 AND2_543( .ZN(g5668), .A1(g49), .A2(g5571) );
  AND2_X1 AND2_544( .ZN(g6338), .A1(g6251), .A2(g6067) );
  AND2_X1 AND2_545( .ZN(g5190), .A1(g426), .A2(g4950) );
  AND2_X1 AND2_546( .ZN(g5501), .A1(g5454), .A2(g3478) );
  AND2_X1 AND2_547( .ZN(g2551), .A1(g715), .A2(g1826) );
  AND2_X1 AND2_548( .ZN(g5156), .A1(g434), .A2(g4877) );
  AND2_X1 AND2_549( .ZN(g5356), .A1(g5265), .A2(g1902) );
  AND2_X1 AND2_550( .ZN(g4277), .A1(g3936), .A2(g942) );
  AND2_X1 AND2_551( .ZN(g5942), .A1(g5117), .A2(g5797) );
  AND2_X1 AND2_552( .ZN(g4789), .A1(g3551), .A2(g4632) );
  AND2_X1 AND2_553( .ZN(g3316), .A1(g2748), .A2(g2894) );
  AND2_X1 AND2_554( .ZN(g3434), .A1(g2850), .A2(g857) );
  AND2_X1 AND2_555( .ZN(g5954), .A1(g5121), .A2(g5813) );
  AND2_X1 AND2_556( .ZN(g5163), .A1(g402), .A2(g4950) );
  AND2_X1 AND2_557( .ZN(g6098), .A1(g1209), .A2(g5753) );
  AND2_X1 AND2_558( .ZN(g3147), .A1(g2419), .A2(g59) );
  AND2_X1 AND2_559( .ZN(g5363), .A1(g4439), .A2(g5179) );
  AND2_X1 AND2_560( .ZN(g3681), .A1(g2234), .A2(g2806) );
  AND2_X1 AND2_561( .ZN(g5053), .A1(g4599), .A2(g4808) );
  AND2_X1 AND2_562( .ZN(g3697), .A1(g2796), .A2(g2481) );
  AND2_X1 AND2_563( .ZN(g5157), .A1(g496), .A2(g4904) );
  AND2_X1 AND2_564( .ZN(g5357), .A1(g398), .A2(g5220) );
  AND3_X1 AND3_21( .ZN(g4244), .A1(g1749), .A2(g4004), .A3(g1609) );
  AND2_X1 AND2_565( .ZN(g4340), .A1(g3972), .A2(g3291) );
  AND2_X2 AND2_566( .ZN(g3936), .A1(g3551), .A2(g940) );
  AND2_X1 AND2_567( .ZN(g3117), .A1(g218), .A2(g2367) );
  AND2_X1 AND2_568( .ZN(g3317), .A1(g2722), .A2(g2895) );
  AND2_X1 AND2_569( .ZN(g4035), .A1(g437), .A2(g3388) );
  AND2_X1 AND2_570( .ZN(g918), .A1(g610), .A2(g602) );
  AND2_X1 AND2_571( .ZN(g6086), .A1(g1143), .A2(g5742) );
  AND2_X1 AND2_572( .ZN(g4214), .A1(g1822), .A2(g4045) );
  AND2_X1 AND2_573( .ZN(g1620), .A1(g1056), .A2(g1084) );
  AND2_X1 AND2_574( .ZN(g3784), .A1(g114), .A2(g3251) );
  AND2_X1 AND2_575( .ZN(g2916), .A1(g1030), .A2(g2113) );
  AND2_X1 AND2_576( .ZN(g3479), .A1(g345), .A2(g2957) );
  AND2_X1 AND2_577( .ZN(g6131), .A1(g5593), .A2(g5975) );
  AND2_X1 AND2_578( .ZN(g3668), .A1(g2568), .A2(g3124) );
  AND2_X1 AND2_579( .ZN(g6331), .A1(g3891), .A2(g6212) );
  AND2_X1 AND2_580( .ZN(g4236), .A1(g654), .A2(g3907) );
  AND2_X1 AND2_581( .ZN(g3294), .A1(g139), .A2(g2870) );
  AND2_X1 AND2_582( .ZN(g5949), .A1(g5119), .A2(g5805) );
  AND2_X1 AND2_583( .ZN(g3190), .A1(g260), .A2(g2535) );
  AND2_X1 AND2_584( .ZN(g6766), .A1(g6750), .A2(g2986) );
  AND2_X1 AND2_585( .ZN(g3156), .A1(g242), .A2(g2464) );
  AND2_X1 AND2_586( .ZN(g3356), .A1(g248), .A2(g2888) );
  AND2_X1 AND2_587( .ZN(g5646), .A1(g4502), .A2(g5544) );
  AND2_X1 AND2_588( .ZN(g2873), .A1(g1845), .A2(g1861) );
  AND2_X1 AND2_589( .ZN(g6748), .A1(g6733), .A2(g6732) );
  AND2_X1 AND2_590( .ZN(g5603), .A1(g5504), .A2(g4911) );
  AND2_X1 AND2_591( .ZN(g5484), .A1(g378), .A2(g5331) );
  AND2_X1 AND2_592( .ZN(g4928), .A1(g148), .A2(g4723) );
  AND2_X1 AND2_593( .ZN(g3704), .A1(g2276), .A2(g2841) );
  AND2_X1 AND2_594( .ZN(g4464), .A1(g4272), .A2(g1937) );
  AND2_X1 AND2_595( .ZN(g4785), .A1(g2160), .A2(g4625) );
  AND2_X1 AND2_596( .ZN(g6091), .A1(g1161), .A2(g5753) );
  AND2_X1 AND2_597( .ZN(g3810), .A1(g625), .A2(g3421) );
  AND2_X1 AND2_598( .ZN(g5952), .A1(g5120), .A2(g5809) );
  AND2_X1 AND2_599( .ZN(g5616), .A1(g5505), .A2(g4929) );
  AND2_X1 AND2_600( .ZN(g6718), .A1(g4511), .A2(g6661) );
  AND2_X2 AND2_601( .ZN(g6767), .A1(g6754), .A2(g2986) );
  AND2_X2 AND2_602( .ZN(g3157), .A1(g2422), .A2(g2467) );
  AND2_X2 AND2_603( .ZN(g3357), .A1(g242), .A2(g2889) );
  AND2_X1 AND2_604( .ZN(g4489), .A1(g2166), .A2(g4206) );
  AND2_X1 AND2_605( .ZN(g2770), .A1(g2518), .A2(g1972) );
  AND2_X1 AND2_606( .ZN(g4471), .A1(g4253), .A2(g332) );
  AND2_X1 AND2_607( .ZN(g5503), .A1(g366), .A2(g5384) );
  AND2_X1 AND2_608( .ZN(g3626), .A1(g3031), .A2(g2727) );
  AND2_X1 AND2_609( .ZN(g4038), .A1(g430), .A2(g3388) );
  AND2_X1 AND2_610( .ZN(g5617), .A1(g5061), .A2(g5524) );
  AND2_X1 AND2_611( .ZN(g3683), .A1(g3150), .A2(g2813) );
  AND2_X1 AND2_612( .ZN(g4836), .A1(g4527), .A2(g4523) );
  AND2_X1 AND2_613( .ZN(g2138), .A1(g1639), .A2(g809) );
  AND2_X1 AND2_614( .ZN(g3661), .A1(g2234), .A2(g2778) );
  AND2_X1 AND2_615( .ZN(g6247), .A1(g504), .A2(g5893) );
  AND2_X1 AND2_616( .ZN(g3627), .A1(g2473), .A2(g3067) );
  AND2_X1 AND2_617( .ZN(g5945), .A1(g5118), .A2(g5801) );
  AND2_X1 AND2_618( .ZN(g2808), .A1(g2009), .A2(g1581) );
  AND2_X1 AND2_619( .ZN(g3292), .A1(g2214), .A2(g2667) );
  AND2_X1 AND2_620( .ZN(g3646), .A1(g2179), .A2(g2756) );
  AND2_X1 AND2_621( .ZN(g2759), .A1(g2473), .A2(g1966) );
  AND2_X1 AND2_622( .ZN(g6910), .A1(g6892), .A2(g6891) );
  AND2_X1 AND2_623( .ZN(g3603), .A1(g2370), .A2(g3019) );
  AND2_X1 AND2_624( .ZN(g3484), .A1(g349), .A2(g2958) );
  AND2_X1 AND2_625( .ZN(g5482), .A1(g370), .A2(g5331) );
  AND2_X1 AND2_626( .ZN(g3702), .A1(g2284), .A2(g2839) );
  AND2_X2 AND2_627( .ZN(g6066), .A1(g5824), .A2(g1721) );
  AND2_X1 AND2_628( .ZN(g5214), .A1(g562), .A2(g5025) );
  AND2_X1 AND2_629( .ZN(g3616), .A1(g2397), .A2(g3049) );
  AND2_X1 AND2_630( .ZN(g6055), .A1(g5824), .A2(g1696) );
  AND2_X1 AND2_631( .ZN(g6133), .A1(g5723), .A2(g5975) );
  AND2_X1 AND2_632( .ZN(g5663), .A1(g4513), .A2(g5550) );
  AND2_X1 AND2_633( .ZN(g6333), .A1(g3896), .A2(g6212) );
  AND2_X1 AND2_634( .ZN(g2419), .A1(g1808), .A2(g54) );
  AND2_X1 AND2_635( .ZN(g3764), .A1(g551), .A2(g3480) );
  AND2_X1 AND2_636( .ZN(g5402), .A1(g370), .A2(g5266) );
  AND2_X1 AND2_637( .ZN(g5236), .A1(g269), .A2(g4915) );
  AND2_X1 AND2_638( .ZN(g4708), .A1(g578), .A2(g4541) );
  AND2_X1 AND2_639( .ZN(g5556), .A1(g5015), .A2(g5445) );
  AND2_X1 AND2_640( .ZN(g4219), .A1(g3911), .A2(g1655) );
  AND2_X1 AND2_641( .ZN(g3277), .A1(g2174), .A2(g2625) );
  AND2_X1 AND2_642( .ZN(g3617), .A1(g2609), .A2(g2317) );
  AND2_X1 AND2_643( .ZN(g6093), .A1(g1177), .A2(g5742) );
  AND2_X2 AND2_644( .ZN(g2897), .A1(g1030), .A2(g2062) );
  AND2_X2 AND2_645( .ZN(g6256), .A1(g1696), .A2(g6040) );
  AND2_X1 AND2_646( .ZN(g4176), .A1(g386), .A2(g3901) );
  AND2_X1 AND2_647( .ZN(g6816), .A1(g6784), .A2(g3346) );
  AND2_X1 AND2_648( .ZN(g4829), .A1(g4526), .A2(g4522) );
  AND2_X1 AND2_649( .ZN(g6263), .A1(g1711), .A2(g6052) );
  AND2_X1 AND2_650( .ZN(g5194), .A1(g586), .A2(g4874) );
  AND2_X1 AND2_651( .ZN(g3709), .A1(g2284), .A2(g2845) );
  AND2_X1 AND2_652( .ZN(g5557), .A1(g5016), .A2(g5448) );
  AND2_X1 AND2_653( .ZN(g3340), .A1(g2772), .A2(g2915) );
  AND2_X1 AND2_654( .ZN(g6631), .A1(g1838), .A2(g6545) );
  AND2_X1 AND2_655( .ZN(g3907), .A1(g650), .A2(g3522) );
  AND2_X1 AND2_656( .ZN(g4177), .A1(g3933), .A2(g1372) );
  AND2_X1 AND2_657( .ZN(g5948), .A1(g5779), .A2(g5407) );
  AND2_X1 AND2_658( .ZN(g4377), .A1(g457), .A2(g3791) );
  AND2_X1 AND2_659( .ZN(g3690), .A1(g2276), .A2(g2827) );
  AND2_X1 AND2_660( .ZN(g5955), .A1(g5782), .A2(g5420) );
  AND2_X1 AND2_661( .ZN(g5350), .A1(g5325), .A2(g3453) );
  AND2_X1 AND2_662( .ZN(g4199), .A1(g628), .A2(g3810) );
  AND2_X1 AND2_663( .ZN(g5438), .A1(g5224), .A2(g3769) );
  AND2_X1 AND2_664( .ZN(g2868), .A1(g1316), .A2(g1861) );
  AND2_X1 AND2_665( .ZN(g3310), .A1(g224), .A2(g2871) );
  AND2_X1 AND2_666( .ZN(g4797), .A1(g4593), .A2(g4643) );
  AND2_X1 AND2_667( .ZN(g5212), .A1(g561), .A2(g5025) );
  AND2_X1 AND2_668( .ZN(g3663), .A1(g2215), .A2(g2779) );
  AND2_X1 AND2_669( .ZN(g2793), .A1(g2568), .A2(g1991) );
  AND2_X1 AND2_670( .ZN(g2015), .A1(g616), .A2(g1419) );
  AND2_X1 AND2_671( .ZN(g4344), .A1(g3981), .A2(g3306) );
  AND2_X1 AND2_672( .ZN(g5229), .A1(g545), .A2(g4980) );
  AND2_X1 AND2_673( .ZN(g6772), .A1(g6746), .A2(g3312) );
  AND2_X1 AND2_674( .ZN(g3762), .A1(g2672), .A2(g3500) );
  AND2_X1 AND2_675( .ZN(g4694), .A1(g1481), .A2(g4578) );
  AND2_X1 AND2_676( .ZN(g3657), .A1(g2734), .A2(g2357) );
  AND2_X1 AND2_677( .ZN(g2721), .A1(g2397), .A2(g1922) );
  AND2_X1 AND2_678( .ZN(g4488), .A1(g1633), .A2(g4202) );
  AND2_X1 AND2_679( .ZN(g4701), .A1(g4596), .A2(g1378) );
  AND2_X1 AND2_680( .ZN(g3928), .A1(g3512), .A2(g478) );
  AND3_X1 AND3_22( .ZN(g6474), .A1(g2138), .A2(g2036), .A3(g6397) );
  AND2_X1 AND2_681( .ZN(g3899), .A1(g323), .A2(g3441) );
  AND2_X1 AND2_682( .ZN(g3464), .A1(g341), .A2(g2956) );
  AND2_X1 AND2_683( .ZN(g5620), .A1(g5507), .A2(g4938) );
  AND2_X2 AND2_684( .ZN(g4870), .A1(g4779), .A2(g1884) );
  AND2_X2 AND2_685( .ZN(g3295), .A1(g2660), .A2(g2647) );
  AND2_X1 AND2_686( .ZN(g2671), .A1(g2263), .A2(g2296) );
  AND2_X1 AND2_687( .ZN(g1576), .A1(g1101), .A2(g1094) );
  AND2_X1 AND2_688( .ZN(g3844), .A1(g3540), .A2(g1665) );
  AND3_X1 AND3_23( .ZN(g1716), .A1(g821), .A2(g774), .A3(g784) );
  AND2_X1 AND2_689( .ZN(g3089), .A1(g212), .A2(g2336) );
  AND2_X1 AND2_690( .ZN(g3731), .A1(g331), .A2(g3441) );
  AND2_X1 AND2_691( .ZN(g3489), .A1(g2607), .A2(g1861) );
  AND2_X1 AND2_692( .ZN(g5192), .A1(g1046), .A2(g4894) );
  AND2_X1 AND2_693( .ZN(g5485), .A1(g382), .A2(g5331) );
  AND2_X1 AND2_694( .ZN(g5941), .A1(g5777), .A2(g5399) );
  AND2_X1 AND2_695( .ZN(g4230), .A1(g3756), .A2(g1861) );
  AND2_X1 AND2_696( .ZN(g6126), .A1(g5711), .A2(g5958) );
  AND2_X1 AND2_697( .ZN(g6326), .A1(g3833), .A2(g6194) );
  AND2_X1 AND2_698( .ZN(g4033), .A1(g426), .A2(g3388) );
  AND2_X2 AND2_699( .ZN(g3814), .A1(g913), .A2(g3546) );
  AND2_X2 AND2_700( .ZN(g2758), .A1(g2497), .A2(g1963) );
  AND2_X1 AND2_701( .ZN(g3350), .A1(g3150), .A2(g1928) );
  AND2_X1 AND2_702( .ZN(g2861), .A1(g2120), .A2(g1654) );
  AND2_X1 AND2_703( .ZN(g6924), .A1(g6920), .A2(g6919) );
  AND2_X1 AND2_704( .ZN(g5176), .A1(g410), .A2(g4950) );
  AND2_X1 AND2_705( .ZN(g4395), .A1(g445), .A2(g3800) );
  AND2_X1 AND2_706( .ZN(g5376), .A1(g170), .A2(g5255) );
  AND2_X1 AND2_707( .ZN(g5911), .A1(g5817), .A2(g5670) );
  AND2_X1 AND2_708( .ZN(g2846), .A1(g619), .A2(g2015) );
  AND2_X1 AND2_709( .ZN(g6127), .A1(g5714), .A2(g5975) );
  AND2_X1 AND2_710( .ZN(g6327), .A1(g3884), .A2(g6212) );
  AND2_X1 AND2_711( .ZN(g5225), .A1(g669), .A2(g5054) );
  AND2_X1 AND2_712( .ZN(g4342), .A1(g3978), .A2(g3299) );
  AND2_X1 AND2_713( .ZN(g6146), .A1(g3192), .A2(g5997) );
  AND2_X1 AND2_714( .ZN(g6346), .A1(g6274), .A2(g6087) );
  AND2_X1 AND2_715( .ZN(g2018), .A1(g1423), .A2(g1254) );
  AND2_X1 AND2_716( .ZN(g4354), .A1(g437), .A2(g3777) );
  AND4_X1 AND4_4( .ZN(I5352), .A1(g3529), .A2(g3531), .A3(g3535), .A4(g3538) );
  AND2_X1 AND2_717( .ZN(g5177), .A1(g445), .A2(g4877) );
  AND2_X1 AND2_718( .ZN(g6240), .A1(g4205), .A2(g5888) );
  AND2_X1 AND2_719( .ZN(g3620), .A1(g2422), .A2(g3060) );
  AND2_X1 AND2_720( .ZN(g1027), .A1(g598), .A2(g567) );
  AND2_X1 AND2_721( .ZN(g2685), .A1(g2370), .A2(g1887) );
  AND2_X1 AND2_722( .ZN(g2700), .A1(g2370), .A2(g1908) );
  AND2_X1 AND2_723( .ZN(g2021), .A1(g835), .A2(g1436) );
  AND2_X1 AND2_724( .ZN(g6316), .A1(g3855), .A2(g6194) );
  AND2_X1 AND2_725( .ZN(g5898), .A1(g5800), .A2(g5647) );
  AND2_X1 AND2_726( .ZN(g4401), .A1(g426), .A2(g3802) );
  AND2_X1 AND2_727( .ZN(g1514), .A1(g1017), .A2(g1011) );
  AND2_X1 AND2_728( .ZN(g5900), .A1(g5804), .A2(g5658) );
  AND2_X1 AND2_729( .ZN(g2950), .A1(g2156), .A2(g1612) );
  AND2_X1 AND2_730( .ZN(g4761), .A1(g4567), .A2(g1674) );
  AND2_X1 AND2_731( .ZN(g5245), .A1(g297), .A2(g4915) );
  AND2_X1 AND2_732( .ZN(g1763), .A1(g478), .A2(g1119) );
  AND2_X1 AND2_733( .ZN(g4828), .A1(g4510), .A2(g4508) );
  AND2_X2 AND2_734( .ZN(g3298), .A1(g2231), .A2(g2679) );
  AND2_X2 AND2_735( .ZN(g4830), .A1(g4529), .A2(g4525) );
  AND2_X2 AND2_736( .ZN(g5144), .A1(g166), .A2(g5099) );
  AND2_X2 AND2_737( .ZN(g4592), .A1(g3147), .A2(g4281) );
  AND2_X1 AND2_738( .ZN(g6914), .A1(g6895), .A2(g6893) );
  AND2_X1 AND2_739( .ZN(g2101), .A1(g1001), .A2(g1543) );
  AND2_X1 AND2_740( .ZN(g5488), .A1(g394), .A2(g5331) );
  AND2_X1 AND2_741( .ZN(g4932), .A1(g157), .A2(g4727) );
  AND2_X1 AND2_742( .ZN(g1416), .A1(g913), .A2(g266) );
  AND2_X1 AND2_743( .ZN(g5701), .A1(g5683), .A2(g3813) );
  AND2_X1 AND2_744( .ZN(g6317), .A1(g3862), .A2(g6194) );
  AND2_X1 AND2_745( .ZN(g5215), .A1(g4864), .A2(g5090) );
  AND2_X1 AND2_746( .ZN(g5951), .A1(g5780), .A2(g5411) );
  AND2_X1 AND2_747( .ZN(g4677), .A1(g4652), .A2(g4646) );
  AND2_X1 AND2_748( .ZN(g3176), .A1(g2422), .A2(g2494) );
  AND2_X1 AND2_749( .ZN(g3376), .A1(g3104), .A2(g1979) );
  AND2_X1 AND2_750( .ZN(g3286), .A1(g2196), .A2(g2656) );
  AND2_X1 AND2_751( .ZN(g3765), .A1(g554), .A2(g3485) );
  AND2_X1 AND2_752( .ZN(g4349), .A1(g441), .A2(g3775) );
  AND2_X1 AND2_753( .ZN(g6060), .A1(g5824), .A2(g1703) );
  AND4_X1 AND4_5( .ZN(g1595), .A1(g729), .A2(g719), .A3(g766), .A4(I2566) );
  AND4_X1 AND4_6( .ZN(I5359), .A1(g3518), .A2(g3521), .A3(g3526), .A4(g3530) );
  AND2_X1 AND2_754( .ZN(g3610), .A1(g2397), .A2(g3034) );
  AND3_X1 AND3_24( .ZN(g6739), .A1(g6715), .A2(g815), .A3(g5242) );
  AND4_X1 AND4_7( .ZN(g1612), .A1(g784), .A2(g774), .A3(g821), .A4(I2574) );
  AND2_X1 AND2_755( .ZN(g3324), .A1(g230), .A2(g2875) );
  AND2_X2 AND2_756( .ZN(g6079), .A1(g1236), .A2(g5753) );
  AND2_X2 AND2_757( .ZN(g5122), .A1(g193), .A2(g4662) );
  AND2_X1 AND2_758( .ZN(g3377), .A1(g3118), .A2(g2931) );
  AND2_X1 AND2_759( .ZN(g4352), .A1(g3988), .A2(g3331) );
  AND2_X1 AND2_760( .ZN(g4867), .A1(g4811), .A2(g3872) );
  AND2_X1 AND2_761( .ZN(g6156), .A1(g2591), .A2(g6015) );
  AND2_X1 AND2_762( .ZN(g3287), .A1(g135), .A2(g2865) );
  AND2_X1 AND2_763( .ZN(g5096), .A1(g4794), .A2(g4647) );
  AND2_X1 AND2_764( .ZN(g4186), .A1(g3973), .A2(g1395) );
  AND2_X1 AND2_765( .ZN(g5496), .A1(g5446), .A2(g3457) );
  AND2_X1 AND2_766( .ZN(g6250), .A1(g1692), .A2(g6036) );
  AND2_X1 AND2_767( .ZN(g4170), .A1(g382), .A2(g3900) );
  AND3_X1 AND3_25( .ZN(g4280), .A1(g2138), .A2(g1764), .A3(g4007) );
  AND2_X1 AND2_768( .ZN(g3144), .A1(g236), .A2(g2440) );
  AND2_X1 AND2_769( .ZN(g3344), .A1(g242), .A2(g2885) );
  AND2_X1 AND2_770( .ZN(g5142), .A1(g148), .A2(g5099) );
  AND2_X1 AND2_771( .ZN(g3819), .A1(g964), .A2(g3437) );
  AND2_X1 AND2_772( .ZN(g6912), .A1(g6899), .A2(g6897) );
  AND2_X1 AND2_773( .ZN(g3694), .A1(g3147), .A2(g64) );
  AND2_X1 AND2_774( .ZN(g6157), .A1(g3158), .A2(g5997) );
  AND2_X1 AND2_775( .ZN(g5481), .A1(g366), .A2(g5331) );
  AND2_X1 AND2_776( .ZN(g3701), .A1(g2268), .A2(g2838) );
  AND2_X1 AND2_777( .ZN(g5497), .A1(g5447), .A2(g3458) );
  AND2_X1 AND2_778( .ZN(g5154), .A1(g500), .A2(g4993) );
  AND2_X1 AND2_779( .ZN(g5354), .A1(g5249), .A2(g2903) );
  AND2_X1 AND2_780( .ZN(g4461), .A1(g4241), .A2(g2919) );
  AND2_X1 AND2_781( .ZN(g4756), .A1(g3816), .A2(g4587) );
  AND2_X1 AND2_782( .ZN(g4046), .A1(I5351), .A2(I5352) );
  AND2_X1 AND2_783( .ZN(g5218), .A1(g564), .A2(g5025) );
  AND2_X1 AND2_784( .ZN(g3650), .A1(g2660), .A2(g2347) );
  AND2_X1 AND2_785( .ZN(g4345), .A1(g3982), .A2(g3308) );
  AND2_X1 AND2_786( .ZN(g3336), .A1(g2760), .A2(g1911) );
  AND2_X1 AND2_787( .ZN(g3768), .A1(g3448), .A2(g1528) );
  AND2_X1 AND2_788( .ZN(g4159), .A1(g370), .A2(g3890) );
  AND2_X1 AND2_789( .ZN(g4359), .A1(g434), .A2(g3782) );
  AND2_X1 AND2_790( .ZN(g3806), .A1(g3384), .A2(g2024) );
  AND2_X1 AND2_791( .ZN(g4416), .A1(g3905), .A2(g1481) );
  AND2_X1 AND2_792( .ZN(g3887), .A1(g3276), .A2(g1861) );
  AND2_X1 AND2_793( .ZN(g3122), .A1(g2435), .A2(g1394) );
  AND2_X1 AND2_794( .ZN(g2732), .A1(g2449), .A2(g1940) );
  AND2_X1 AND2_795( .ZN(g4047), .A1(g453), .A2(g3388) );
  AND2_X1 AND2_796( .ZN(g6646), .A1(g6577), .A2(g6232) );
  AND3_X1 AND3_26( .ZN(g3433), .A1(g1359), .A2(g2831), .A3(g905) );
  AND2_X1 AND2_797( .ZN(g5953), .A1(g5781), .A2(g5415) );
  AND2_X1 AND2_798( .ZN(g6084), .A1(g1123), .A2(g5753) );
  AND2_X1 AND2_799( .ZN(g6603), .A1(g6581), .A2(g6236) );
  AND2_X1 AND2_800( .ZN(g4874), .A1(g582), .A2(g4708) );
  AND2_X1 AND2_801( .ZN(g5677), .A1(g69), .A2(g5575) );
  AND2_X1 AND2_802( .ZN(g3195), .A1(g2473), .A2(g2541) );
  AND2_X1 AND2_803( .ZN(g3337), .A1(g2796), .A2(g2913) );
  AND3_X1 AND3_27( .ZN(I4040), .A1(g1279), .A2(g2025), .A3(g1267) );
  AND2_X1 AND2_804( .ZN(g5149), .A1(g4910), .A2(g1480) );
  AND2_X1 AND2_805( .ZN(g5349), .A1(g5324), .A2(g3451) );
  AND2_X1 AND2_806( .ZN(g5198), .A1(g558), .A2(g5025) );
  AND2_X1 AND2_807( .ZN(g5398), .A1(g366), .A2(g5261) );
  AND2_X1 AND2_808( .ZN(g1570), .A1(g634), .A2(g1027) );
  AND2_X1 AND2_809( .ZN(g6647), .A1(g6578), .A2(g6233) );
  AND2_X1 AND2_810( .ZN(g1691), .A1(g821), .A2(g774) );
  AND2_X1 AND2_811( .ZN(g3692), .A1(g2268), .A2(g2829) );
  AND2_X1 AND2_812( .ZN(g3726), .A1(g119), .A2(g3251) );
  AND2_X1 AND2_813( .ZN(g3154), .A1(g2039), .A2(g1410) );
  AND2_X1 AND2_814( .ZN(g4800), .A1(g4648), .A2(g4296) );
  AND2_X1 AND2_815( .ZN(g5152), .A1(g430), .A2(g4950) );
  AND2_X1 AND2_816( .ZN(g6320), .A1(g3869), .A2(g6194) );
  AND2_X1 AND2_817( .ZN(g5211), .A1(g4860), .A2(g5086) );
  AND2_X1 AND2_818( .ZN(g5186), .A1(g422), .A2(g4950) );
  AND2_X1 AND2_819( .ZN(g5599), .A1(g5049), .A2(g5512) );
  AND2_X1 AND2_820( .ZN(g4490), .A1(g2941), .A2(g4210) );
  AND2_X1 AND2_821( .ZN(g3293), .A1(g212), .A2(g2864) );
  AND2_X1 AND2_822( .ZN(g6771), .A1(g6758), .A2(g3483) );
  AND2_X1 AND2_823( .ZN(g3329), .A1(g2748), .A2(g2907) );
  AND2_X1 AND2_824( .ZN(g5170), .A1(g5091), .A2(g2111) );
  AND2_X1 AND2_825( .ZN(g4456), .A1(g3829), .A2(g4229) );
  AND2_X1 AND2_826( .ZN(g6299), .A1(g5530), .A2(g6163) );
  AND2_X1 AND2_827( .ZN(g4348), .A1(g3987), .A2(g3322) );
  AND2_X1 AND2_828( .ZN(g3727), .A1(g122), .A2(g3251) );
  AND2_X1 AND2_829( .ZN(g2937), .A1(g2160), .A2(g931) );
  AND2_X1 AND2_830( .ZN(g4355), .A1(g430), .A2(g3778) );
  AND2_X1 AND2_831( .ZN(g5939), .A1(g5776), .A2(g5395) );
  AND3_X1 AND3_28( .ZN(g2294), .A1(g1716), .A2(g791), .A3(g798) );
  AND2_X1 AND2_832( .ZN(g4698), .A1(g4586), .A2(g2106) );
  AND2_X2 AND2_833( .ZN(g5483), .A1(g374), .A2(g5331) );
  AND2_X2 AND2_834( .ZN(g3703), .A1(g2284), .A2(g2840) );
  AND3_X1 AND3_29( .ZN(g6738), .A1(g6713), .A2(g809), .A3(g5242) );
  AND2_X1 AND2_835( .ZN(g2156), .A1(g815), .A2(g1642) );
  AND2_X1 AND2_836( .ZN(g6244), .A1(g4759), .A2(g5891) );
  AND2_X1 AND2_837( .ZN(g2356), .A1(g1603), .A2(g269) );
  AND2_X1 AND2_838( .ZN(g6140), .A1(g5587), .A2(g5975) );
  AND2_X1 AND2_839( .ZN(g3953), .A1(g3554), .A2(g188) );
  AND2_X1 AND2_840( .ZN(g6340), .A1(g6257), .A2(g6069) );
  AND2_X1 AND2_841( .ZN(g5187), .A1(g457), .A2(g4877) );
  AND2_X1 AND2_842( .ZN(g1628), .A1(g815), .A2(g809) );
  AND2_X1 AND2_843( .ZN(g4167), .A1(g378), .A2(g3898) );
  AND2_X1 AND2_844( .ZN(g6082), .A1(g1123), .A2(g5742) );
  AND2_X1 AND2_845( .ZN(g4367), .A1(g193), .A2(g3788) );
  AND2_X1 AND2_846( .ZN(g4872), .A1(g4760), .A2(g1549) );
  AND2_X1 AND2_847( .ZN(g4057), .A1(g422), .A2(g3388) );
  AND2_X1 AND2_848( .ZN(g5904), .A1(g5812), .A2(g5664) );
  AND2_X1 AND2_849( .ZN(g5200), .A1(g559), .A2(g5025) );
  AND2_X1 AND2_850( .ZN(g4457), .A1(g4261), .A2(g2902) );
  AND2_X1 AND2_851( .ZN(g5446), .A1(g4537), .A2(g5241) );
  AND2_X1 AND2_852( .ZN(g3349), .A1(g2783), .A2(g1925) );
  AND2_X1 AND2_853( .ZN(g2053), .A1(g1094), .A2(g1675) );
  AND2_X1 AND2_854( .ZN(g5145), .A1(g175), .A2(g5099) );
  AND2_X1 AND2_855( .ZN(g6915), .A1(g6906), .A2(g6905) );
  AND2_X1 AND2_856( .ZN(g4834), .A1(g4534), .A2(g4531) );
  AND2_X1 AND2_857( .ZN(g4686), .A1(g4590), .A2(g1348) );
  AND2_X1 AND2_858( .ZN(g5191), .A1(g461), .A2(g4877) );
  AND2_X1 AND2_859( .ZN(g3699), .A1(g2276), .A2(g2836) );
  AND2_X1 AND2_860( .ZN(g4598), .A1(g1978), .A2(g4253) );
  AND2_X1 AND2_861( .ZN(g5637), .A1(g4499), .A2(g5543) );
  AND2_X1 AND2_862( .ZN(g5159), .A1(g536), .A2(g4967) );
  AND2_X1 AND2_863( .ZN(g5359), .A1(g4428), .A2(g5155) );
  AND2_X1 AND2_864( .ZN(g4253), .A1(g1861), .A2(g3819) );
  AND2_X1 AND2_865( .ZN(g3644), .A1(g2197), .A2(g2755) );
  AND2_X1 AND2_866( .ZN(g3319), .A1(g2688), .A2(g2675) );
  AND2_X1 AND2_867( .ZN(g3352), .A1(g2796), .A2(g2920) );
  AND2_X1 AND2_868( .ZN(g5047), .A1(g3954), .A2(g4806) );
  AND3_X1 AND3_30( .ZN(g5447), .A1(g4545), .A2(g5256), .A3(g2311) );
  AND2_X1 AND2_869( .ZN(g4687), .A1(g4493), .A2(g1542) );
  AND2_X1 AND2_870( .ZN(g3186), .A1(g2449), .A2(g2515) );
  AND2_X1 AND2_871( .ZN(g3170), .A1(g254), .A2(g2485) );
  AND2_X1 AND2_872( .ZN(g3614), .A1(g2998), .A2(g2691) );
  AND2_X1 AND2_873( .ZN(g3325), .A1(g224), .A2(g2876) );
  AND2_X2 AND2_874( .ZN(g4341), .A1(g3977), .A2(g3297) );
  AND2_X2 AND2_875( .ZN(g2782), .A1(g2518), .A2(g1985) );
  AND2_X2 AND2_876( .ZN(g6295), .A1(g5379), .A2(g6162) );
  AND2_X1 AND2_877( .ZN(g3280), .A1(g2177), .A2(g2637) );
  AND2_X1 AND2_878( .ZN(g5017), .A1(g4784), .A2(g1679) );
  AND2_X1 AND2_879( .ZN(g4691), .A1(g4581), .A2(g2098) );
  AND2_X1 AND2_880( .ZN(g5935), .A1(g5112), .A2(g5784) );
  AND2_X1 AND2_881( .ZN(g2949), .A1(g830), .A2(g1861) );
  AND4_X1 AND4_8( .ZN(I5351), .A1(g3511), .A2(g3517), .A3(g3520), .A4(g3525) );
  AND2_X1 AND2_882( .ZN(g5234), .A1(g197), .A2(g4915) );
  AND2_X1 AND2_883( .ZN(g3636), .A1(g2701), .A2(g2327) );
  AND3_X1 AND3_31( .ZN(g2292), .A1(g1706), .A2(g736), .A3(g743) );
  AND2_X1 AND2_884( .ZN(g6089), .A1(g1143), .A2(g5731) );
  AND2_X1 AND2_885( .ZN(g6731), .A1(g6717), .A2(g4427) );
  AND2_X1 AND2_886( .ZN(g6557), .A1(g1595), .A2(g6469) );
  AND2_X1 AND2_887( .ZN(g4358), .A1(g3991), .A2(g3343) );
  AND2_X1 AND2_888( .ZN(g2084), .A1(g1577), .A2(g1563) );
  AND2_X1 AND2_889( .ZN(g2850), .A1(g2018), .A2(g1255) );
  AND2_X1 AND2_890( .ZN(g5213), .A1(g4862), .A2(g5087) );
  AND2_X1 AND2_891( .ZN(g6254), .A1(g532), .A2(g5897) );
  AND2_X1 AND2_892( .ZN(g6150), .A1(g3204), .A2(g6015) );
  AND2_X1 AND2_893( .ZN(g5902), .A1(g5808), .A2(g5661) );
  AND2_X1 AND2_894( .ZN(g3145), .A1(g2397), .A2(g2443) );
  AND2_X1 AND2_895( .ZN(g3345), .A1(g236), .A2(g2886) );
  AND2_X1 AND2_896( .ZN(g6773), .A1(g6762), .A2(g2986) );
  AND2_X1 AND2_897( .ZN(g3763), .A1(g3064), .A2(g3501) );
  AND2_X1 AND2_898( .ZN(g3191), .A1(g2497), .A2(g2538) );
  AND2_X1 AND2_899( .ZN(g4180), .A1(g3929), .A2(g2119) );
  AND2_X1 AND2_900( .ZN(g5166), .A1(g541), .A2(g4967) );
  AND2_X1 AND2_901( .ZN(g3637), .A1(g2822), .A2(g2752) );
  AND2_X1 AND2_902( .ZN(g4832), .A1(g4517), .A2(g4512) );
  AND2_X1 AND2_903( .ZN(g6769), .A1(g6758), .A2(g2986) );
  AND2_X1 AND2_904( .ZN(g3307), .A1(g2242), .A2(g2692) );
  AND2_X1 AND2_905( .ZN(g3359), .A1(g2822), .A2(g2922) );
  AND2_X1 AND2_906( .ZN(g4794), .A1(g4593), .A2(g949) );
  AND2_X1 AND2_907( .ZN(g3757), .A1(g2619), .A2(g3487) );
  AND2_X1 AND2_908( .ZN(g3522), .A1(g646), .A2(g2909) );
  AND2_X1 AND2_909( .ZN(g3315), .A1(g2701), .A2(g1875) );
  AND2_X1 AND2_910( .ZN(g3642), .A1(g3054), .A2(g2754) );
  AND2_X1 AND2_911( .ZN(g3654), .A1(g2518), .A2(g3100) );
  AND2_X1 AND2_912( .ZN(g5619), .A1(g5064), .A2(g5527) );
  AND2_X2 AND2_913( .ZN(g5167), .A1(g5011), .A2(g1556) );
  OR2_X1 OR2_0( .ZN(g3880), .A1(g3658), .A2(g3665) );
  OR2_X1 OR2_1( .ZN(g4440), .A1(g4371), .A2(g4038) );
  OR2_X1 OR2_2( .ZN(g3978), .A1(g3655), .A2(g3117) );
  OR2_X1 OR2_3( .ZN(g6788), .A1(g3760), .A2(g6767) );
  OR2_X1 OR2_4( .ZN(g3935), .A1(g3464), .A2(g2868) );
  OR2_X1 OR2_5( .ZN(g3982), .A1(g3663), .A2(g3127) );
  OR4_X1 OR4_0( .ZN(I8376), .A1(g6315), .A2(g6126), .A3(g6129), .A4(g6146) );
  OR2_X1 OR2_6( .ZN(g5625), .A1(g5495), .A2(g3281) );
  OR2_X1 OR2_7( .ZN(g6298), .A1(g6255), .A2(g6093) );
  OR3_X1 OR3_0( .ZN(g6485), .A1(I8393), .A2(I8394), .A3(I8395) );
  OR2_X1 OR2_8( .ZN(g4655), .A1(g4368), .A2(g3660) );
  OR2_X1 OR2_9( .ZN(g6252), .A1(g5905), .A2(g2381) );
  OR2_X1 OR2_10( .ZN(g6176), .A1(g6068), .A2(g6033) );
  OR4_X1 OR4_1( .ZN(I8377), .A1(g6150), .A2(g6324), .A3(g5180), .A4(g5181) );
  OR2_X1 OR2_11( .ZN(g6286), .A1(g6238), .A2(g6079) );
  OR2_X1 OR2_12( .ZN(g3851), .A1(g3681), .A2(g3146) );
  OR2_X1 OR2_13( .ZN(g3964), .A1(g3634), .A2(g3089) );
  OR2_X1 OR2_14( .ZN(g5659), .A1(g5551), .A2(g5398) );
  OR2_X1 OR2_15( .ZN(g2928), .A1(g2100), .A2(g1582) );
  OR2_X1 OR2_16( .ZN(g6287), .A1(g6241), .A2(g6082) );
  OR2_X1 OR2_17( .ZN(g3989), .A1(g3679), .A2(g3144) );
  OR2_X1 OR2_18( .ZN(g5374), .A1(g5215), .A2(g4947) );
  OR2_X1 OR2_19( .ZN(g3971), .A1(g3644), .A2(g3099) );
  OR2_X1 OR2_20( .ZN(g6781), .A1(g6718), .A2(g6748) );
  OR2_X1 OR2_21( .ZN(g3598), .A1(g2808), .A2(g2821) );
  OR2_X2 OR2_22( .ZN(g4641), .A1(g4347), .A2(g3627) );
  OR2_X1 OR2_23( .ZN(g4450), .A1(g4389), .A2(g4047) );
  OR2_X1 OR2_24( .ZN(g3740), .A1(g3335), .A2(g2747) );
  OR4_X1 OR4_2( .ZN(I8136), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_25( .ZN(g5628), .A1(g5498), .A2(g3292) );
  OR2_X1 OR2_26( .ZN(g5630), .A1(g5501), .A2(g3309) );
  OR2_X1 OR2_27( .ZN(g6114), .A1(g5904), .A2(g5604) );
  OR2_X1 OR2_28( .ZN(g5323), .A1(g5098), .A2(g4802) );
  OR2_X1 OR2_29( .ZN(g5666), .A1(g5555), .A2(g5406) );
  OR4_X1 OR4_3( .ZN(I8137), .A1(g4894), .A2(g4904), .A3(g4993), .A4(g4967) );
  OR3_X1 OR3_1( .ZN(I8395), .A1(g5182), .A2(g5200), .A3(g6280) );
  OR2_X1 OR2_30( .ZN(g3879), .A1(g3704), .A2(g3195) );
  OR4_X1 OR4_4( .ZN(I9057), .A1(g6320), .A2(g6828), .A3(g6830), .A4(g6153) );
  OR2_X1 OR2_31( .ZN(g4092), .A1(g3311), .A2(g2721) );
  OR4_X1 OR4_5( .ZN(I8081), .A1(g4894), .A2(g4904), .A3(g4993), .A4(g4967) );
  OR2_X1 OR2_32( .ZN(g4864), .A1(g4744), .A2(g4490) );
  OR3_X1 OR3_2( .ZN(g6845), .A1(I9064), .A2(I9065), .A3(I9066) );
  OR2_X2 OR2_33( .ZN(g5372), .A1(g5213), .A2(g4942) );
  OR2_X1 OR2_34( .ZN(g5693), .A1(g5632), .A2(g5481) );
  OR2_X1 OR2_35( .ZN(g5804), .A1(g5371), .A2(g5603) );
  OR2_X1 OR2_36( .ZN(g6142), .A1(g5909), .A2(g3806) );
  OR2_X1 OR2_37( .ZN(I8129), .A1(g4915), .A2(g5025) );
  OR4_X1 OR4_6( .ZN(g6481), .A1(I8367), .A2(I8368), .A3(I8369), .A4(I8370) );
  OR2_X1 OR2_38( .ZN(g4651), .A1(g4357), .A2(g3643) );
  OR2_X1 OR2_39( .ZN(g4285), .A1(g3490), .A2(g3887) );
  OR2_X1 OR2_40( .ZN(g4500), .A1(g4243), .A2(g2010) );
  OR3_X1 OR3_3( .ZN(g5202), .A1(g4904), .A2(g4914), .A3(g4894) );
  OR2_X1 OR2_41( .ZN(g3750), .A1(g3372), .A2(g2794) );
  OR2_X1 OR2_42( .ZN(g6267), .A1(g2953), .A2(g5884) );
  OR2_X1 OR2_43( .ZN(g4231), .A1(g3997), .A2(g4000) );
  OR2_X1 OR2_44( .ZN(g6676), .A1(g6631), .A2(g6555) );
  OR2_X1 OR2_45( .ZN(g6293), .A1(g6244), .A2(g6085) );
  OR2_X1 OR2_46( .ZN(g4205), .A1(g3843), .A2(g541) );
  OR2_X1 OR2_47( .ZN(g4634), .A1(g4341), .A2(g3615) );
  OR4_X1 OR4_7( .ZN(I8349), .A1(I8345), .A2(I8346), .A3(I8347), .A4(I8348) );
  OR2_X1 OR2_48( .ZN(g6703), .A1(g6692), .A2(g4831) );
  OR2_X1 OR2_49( .ZN(g3884), .A1(g3666), .A2(g3671) );
  OR2_X1 OR2_50( .ZN(g4444), .A1(g4378), .A2(g4042) );
  OR2_X1 OR2_51( .ZN(g4862), .A1(g4739), .A2(g4489) );
  OR4_X1 OR4_8( .ZN(I8119), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR2_X1 OR2_52( .ZN(g3988), .A1(g3678), .A2(g3143) );
  OR2_X1 OR2_53( .ZN(g5674), .A1(g5558), .A2(g5419) );
  OR2_X1 OR2_54( .ZN(g6747), .A1(g6614), .A2(g6731) );
  OR2_X2 OR2_55( .ZN(g6855), .A1(g6851), .A2(g2085) );
  OR2_X2 OR2_56( .ZN(I8211), .A1(g4915), .A2(g5025) );
  OR4_X1 OR4_9( .ZN(I8386), .A1(g6152), .A2(g6327), .A3(g5183), .A4(g5177) );
  OR2_X1 OR2_57( .ZN(g5680), .A1(g5562), .A2(g5429) );
  OR2_X1 OR2_58( .ZN(g4946), .A1(g4830), .A2(g4833) );
  OR2_X1 OR2_59( .ZN(I8370), .A1(g5214), .A2(g6358) );
  OR2_X1 OR2_60( .ZN(g4436), .A1(g4359), .A2(g4035) );
  OR3_X1 OR3_4( .ZN(I8387), .A1(g5178), .A2(g5209), .A3(g6281) );
  OR2_X1 OR2_61( .ZN(g6274), .A1(g5682), .A2(g5956) );
  OR2_X1 OR2_62( .ZN(g6426), .A1(g6288), .A2(g6119) );
  OR2_X1 OR2_63( .ZN(g6170), .A1(g6061), .A2(g6014) );
  OR2_X1 OR2_64( .ZN(g3996), .A1(g3691), .A2(g3171) );
  OR4_X1 OR4_10( .ZN(I8345), .A1(g6326), .A2(g6135), .A3(g6140), .A4(g6157) );
  OR2_X1 OR2_65( .ZN(g5623), .A1(g5503), .A2(g5357) );
  OR3_X1 OR3_5( .ZN(g6483), .A1(I8385), .A2(I8386), .A3(I8387) );
  OR2_X1 OR2_66( .ZN(g4653), .A1(g4361), .A2(g3652) );
  OR2_X1 OR2_67( .ZN(g3878), .A1(g3703), .A2(g3191) );
  OR2_X1 OR2_68( .ZN(g6790), .A1(g3765), .A2(g6773) );
  OR4_X1 OR4_11( .ZN(I8359), .A1(g5232), .A2(g5236), .A3(g5216), .A4(g5226) );
  OR2_X1 OR2_69( .ZN(g4752), .A1(g4452), .A2(g4155) );
  OR2_X1 OR2_70( .ZN(g6461), .A1(g6353), .A2(g6351) );
  OR2_X1 OR2_71( .ZN(g3981), .A1(g3661), .A2(g3123) );
  OR2_X1 OR2_72( .ZN(g5024), .A1(g4793), .A2(g4600) );
  OR2_X1 OR2_73( .ZN(g4233), .A1(g3912), .A2(g471) );
  OR2_X1 OR2_74( .ZN(g4454), .A1(g4395), .A2(g4051) );
  OR2_X1 OR2_75( .ZN(g5672), .A1(g5557), .A2(g5414) );
  OR2_X1 OR2_76( .ZN(g5077), .A1(g1612), .A2(g4694) );
  OR2_X1 OR2_77( .ZN(g5231), .A1(g5048), .A2(g672) );
  OR2_X1 OR2_78( .ZN(g6307), .A1(g6262), .A2(g6096) );
  OR2_X1 OR2_79( .ZN(g3744), .A1(g3345), .A2(g2759) );
  OR2_X1 OR2_80( .ZN(g6251), .A1(g5668), .A2(g5939) );
  OR2_X1 OR2_81( .ZN(g6447), .A1(g6340), .A2(g5938) );
  OR4_X2 OR4_12( .ZN(I8128), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR2_X1 OR2_82( .ZN(g3864), .A1(g3693), .A2(g3176) );
  OR2_X1 OR2_83( .ZN(g5044), .A1(g4797), .A2(g4602) );
  OR2_X1 OR2_84( .ZN(g4745), .A1(g4468), .A2(g4569) );
  OR2_X1 OR2_85( .ZN(g6272), .A1(g5679), .A2(g5953) );
  OR2_X1 OR2_86( .ZN(g5014), .A1(g4785), .A2(g4583) );
  OR2_X1 OR2_87( .ZN(g3871), .A1(g3701), .A2(g3186) );
  OR4_X1 OR4_13( .ZN(I7970), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR4_X1 OR4_14( .ZN(I8348), .A1(g5229), .A2(g5234), .A3(g5218), .A4(g5225) );
  OR2_X1 OR2_88( .ZN(g6554), .A1(g6337), .A2(g6466) );
  OR4_X1 OR4_15( .ZN(I7987), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_89( .ZN(g5916), .A1(g5728), .A2(g3781) );
  OR4_X1 OR4_16( .ZN(I8118), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR4_X1 OR4_17( .ZN(I8367), .A1(g6313), .A2(g6124), .A3(g6127), .A4(g6144) );
  OR2_X1 OR2_90( .ZN(g6456), .A1(g6346), .A2(g5954) );
  OR4_X1 OR4_18( .ZN(I8393), .A1(g6317), .A2(g6130), .A3(g6133), .A4(g6151) );
  OR2_X1 OR2_91( .ZN(g4086), .A1(g3310), .A2(g2720) );
  OR2_X1 OR2_92( .ZN(g1589), .A1(g1059), .A2(g1045) );
  OR2_X1 OR2_93( .ZN(g6118), .A1(g5911), .A2(g5619) );
  OR2_X1 OR2_94( .ZN(g6167), .A1(g6056), .A2(g6039) );
  OR2_X1 OR2_95( .ZN(g3862), .A1(g3632), .A2(g3641) );
  OR2_X1 OR2_96( .ZN(g6457), .A1(g6352), .A2(g6347) );
  OR2_X1 OR2_97( .ZN(g4635), .A1(g4342), .A2(g3616) );
  OR2_X1 OR2_98( .ZN(g6549), .A1(g6473), .A2(g4247) );
  OR2_X1 OR2_99( .ZN(g6686), .A1(g6259), .A2(g6645) );
  OR2_X1 OR2_100( .ZN(g5532), .A1(g5350), .A2(g3278) );
  OR4_X1 OR4_19( .ZN(g6670), .A1(g6557), .A2(g6634), .A3(g4410), .A4(g2948) );
  OR2_X1 OR2_101( .ZN(g5012), .A1(g4782), .A2(g4580) );
  OR2_X1 OR2_102( .ZN(g4059), .A1(g3466), .A2(g3425) );
  OR2_X1 OR2_103( .ZN(g5281), .A1(g5074), .A2(g5124) );
  OR4_X1 OR4_20( .ZN(I8358), .A1(g5192), .A2(g5153), .A3(g5158), .A4(g5197) );
  OR2_X2 OR2_104( .ZN(g6687), .A1(g6260), .A2(g6646) );
  OR2_X2 OR2_105( .ZN(g3749), .A1(g3371), .A2(g2793) );
  OR2_X2 OR2_106( .ZN(g5808), .A1(g5373), .A2(g5616) );
  OR2_X1 OR2_107( .ZN(g6691), .A1(g6275), .A2(g6603) );
  OR2_X1 OR2_108( .ZN(g3873), .A1(g3649), .A2(g3657) );
  OR2_X1 OR2_109( .ZN(g3869), .A1(g3642), .A2(g3650) );
  OR2_X1 OR2_110( .ZN(g6659), .A1(g6634), .A2(g6631) );
  OR2_X1 OR2_111( .ZN(g4430), .A1(g4349), .A2(g4015) );
  OR2_X1 OR2_112( .ZN(g6239), .A1(g2339), .A2(g6073) );
  OR2_X1 OR2_113( .ZN(g6545), .A1(g6468), .A2(g4244) );
  OR2_X1 OR2_114( .ZN(g4638), .A1(g4345), .A2(g3620) );
  OR2_X1 OR2_115( .ZN(g6794), .A1(g6777), .A2(g3333) );
  OR2_X1 OR2_116( .ZN(g6931), .A1(g6741), .A2(g6929) );
  OR2_X1 OR2_117( .ZN(g3990), .A1(g3684), .A2(g3155) );
  OR2_X1 OR2_118( .ZN(g5385), .A1(g3992), .A2(g5318) );
  OR2_X1 OR2_119( .ZN(g3888), .A1(g3672), .A2(g3682) );
  OR2_X1 OR2_120( .ZN(g5470), .A1(g5359), .A2(g5142) );
  OR2_X1 OR2_121( .ZN(g6300), .A1(g6253), .A2(g6091) );
  OR2_X1 OR2_122( .ZN(g4455), .A1(g4396), .A2(g4052) );
  OR3_X1 OR3_6( .ZN(g6750), .A1(g6670), .A2(g6625), .A3(g6736) );
  OR2_X1 OR2_123( .ZN(g5678), .A1(g5560), .A2(g5428) );
  OR2_X1 OR2_124( .ZN(g3745), .A1(g3356), .A2(g2770) );
  OR2_X1 OR2_125( .ZN(g6440), .A1(g6336), .A2(g5935) );
  OR2_X1 OR2_126( .ZN(g3865), .A1(g3637), .A2(g3648) );
  OR2_X1 OR2_127( .ZN(g3833), .A1(g3602), .A2(g3608) );
  OR2_X1 OR2_128( .ZN(g4021), .A1(g3558), .A2(g2949) );
  OR2_X1 OR2_129( .ZN(g3896), .A1(g3689), .A2(g3697) );
  OR2_X1 OR2_130( .ZN(g5535), .A1(g5353), .A2(g3300) );
  OR2_X1 OR2_131( .ZN(g5015), .A1(g4787), .A2(g4588) );
  OR2_X1 OR2_132( .ZN(g4631), .A1(g4340), .A2(g3611) );
  OR2_X1 OR2_133( .ZN(g5246), .A1(g5077), .A2(g2080) );
  OR2_X1 OR2_134( .ZN(g6792), .A1(g6770), .A2(g3321) );
  OR4_X2 OR4_21( .ZN(I7980), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR4_X1 OR4_22( .ZN(I8360), .A1(I8356), .A2(I8357), .A3(I8358), .A4(I8359) );
  OR2_X1 OR2_135( .ZN(g4441), .A1(g4372), .A2(g4039) );
  OR2_X1 OR2_136( .ZN(g6113), .A1(g5902), .A2(g5601) );
  OR3_X1 OR3_7( .ZN(g5388), .A1(g5318), .A2(g1589), .A3(g3491) );
  OR2_X1 OR2_137( .ZN(I8379), .A1(g5212), .A2(g6357) );
  OR2_X1 OR2_138( .ZN(g5430), .A1(g5161), .A2(g4873) );
  OR2_X1 OR2_139( .ZN(g4458), .A1(g4401), .A2(g4057) );
  OR2_X1 OR2_140( .ZN(g3748), .A1(g3366), .A2(g2782) );
  OR2_X1 OR2_141( .ZN(g6264), .A1(g5675), .A2(g5948) );
  OR2_X1 OR2_142( .ZN(g4074), .A1(g3301), .A2(g2699) );
  OR2_X1 OR2_143( .ZN(g6450), .A1(g6341), .A2(g5940) );
  OR2_X1 OR2_144( .ZN(g4080), .A1(g3302), .A2(g2700) );
  OR2_X1 OR2_145( .ZN(g5066), .A1(g4668), .A2(g4672) );
  OR2_X1 OR2_146( .ZN(g6179), .A1(g6077), .A2(g6051) );
  OR4_X1 OR4_23( .ZN(I8209), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_147( .ZN(g6289), .A1(g6240), .A2(g6081) );
  OR2_X1 OR2_148( .ZN(g6658), .A1(g6132), .A2(g6620) );
  OR2_X1 OR2_149( .ZN(g6271), .A1(g2955), .A2(g5885) );
  OR2_X1 OR2_150( .ZN(g5662), .A1(g5553), .A2(g5402) );
  OR2_X1 OR2_151( .ZN(g5018), .A1(g4791), .A2(g4597) );
  OR2_X1 OR2_152( .ZN(I7972), .A1(g4915), .A2(g5025) );
  OR3_X1 OR3_8( .ZN(g5467), .A1(g3868), .A2(g5318), .A3(g3992) );
  OR2_X1 OR2_153( .ZN(g5816), .A1(g5378), .A2(g5620) );
  OR2_X2 OR2_154( .ZN(g5700), .A1(g5663), .A2(g5488) );
  OR2_X2 OR2_155( .ZN(g4451), .A1(g4390), .A2(g4048) );
  OR2_X1 OR2_156( .ZN(g6864), .A1(g6852), .A2(g2089) );
  OR2_X1 OR2_157( .ZN(g5817), .A1(g5380), .A2(g5621) );
  OR2_X1 OR2_158( .ZN(g3883), .A1(g3709), .A2(g3203) );
  OR2_X1 OR2_159( .ZN(g5605), .A1(g3575), .A2(g5500) );
  OR3_X1 OR3_9( .ZN(I9059), .A1(g5185), .A2(g5198), .A3(g6279) );
  OR2_X1 OR2_160( .ZN(g4443), .A1(g4377), .A2(g4041) );
  OR2_X1 OR2_161( .ZN(g4434), .A1(g4355), .A2(g4033) );
  OR2_X1 OR2_162( .ZN(g5669), .A1(g5556), .A2(g5410) );
  OR2_X1 OR2_163( .ZN(g5368), .A1(g5201), .A2(g4932) );
  OR4_X1 OR4_24( .ZN(I7979), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_164( .ZN(g5531), .A1(g5349), .A2(g3275) );
  OR2_X1 OR2_165( .ZN(g5458), .A1(g3466), .A2(g5311) );
  OR2_X1 OR2_166( .ZN(g6795), .A1(g4867), .A2(g6772) );
  OR2_X1 OR2_167( .ZN(g4936), .A1(g4827), .A2(g4828) );
  OR2_X1 OR2_168( .ZN(g5074), .A1(g4792), .A2(g4598) );
  OR2_X1 OR2_169( .ZN(g5474), .A1(g5363), .A2(g5146) );
  OR2_X1 OR2_170( .ZN(g6926), .A1(g6798), .A2(g6923) );
  OR3_X1 OR3_10( .ZN(g6754), .A1(g6676), .A2(g6625), .A3(g6737) );
  OR2_X1 OR2_171( .ZN(g6273), .A1(g5681), .A2(g5955) );
  OR2_X1 OR2_172( .ZN(g6444), .A1(g6338), .A2(g5936) );
  OR4_X1 OR4_25( .ZN(I8378), .A1(g5173), .A2(g5166), .A3(g5235), .A4(g5245) );
  OR4_X1 OR4_26( .ZN(I8135), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR3_X1 OR3_11( .ZN(g5326), .A1(g5069), .A2(g4410), .A3(g3012) );
  OR3_X1 OR3_12( .ZN(I9066), .A1(g5189), .A2(g5269), .A3(g6400) );
  OR2_X1 OR2_173( .ZN(g6927), .A1(g6799), .A2(g6924) );
  OR2_X1 OR2_174( .ZN(g3751), .A1(g3375), .A2(g2807) );
  OR2_X1 OR2_175( .ZN(g6660), .A1(g6640), .A2(g6637) );
  OR2_X1 OR2_176( .ZN(g6679), .A1(g6637), .A2(g6558) );
  OR4_X1 OR4_27( .ZN(I8208), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_177( .ZN(g6182), .A1(g6047), .A2(g6034) );
  OR3_X2 OR3_13( .ZN(g5327), .A1(g5077), .A2(g4416), .A3(g3028) );
  OR2_X1 OR2_178( .ZN(g3743), .A1(g3344), .A2(g2758) );
  OR2_X1 OR2_179( .ZN(g3856), .A1(g3686), .A2(g3157) );
  OR2_X1 OR2_180( .ZN(g5303), .A1(g5053), .A2(g4768) );
  OR2_X1 OR2_181( .ZN(g5696), .A1(g5637), .A2(g5484) );
  OR2_X1 OR2_182( .ZN(g3992), .A1(g1555), .A2(g3559) );
  OR2_X1 OR2_183( .ZN(g5472), .A1(g5361), .A2(g5144) );
  OR2_X1 OR2_184( .ZN(g3863), .A1(g3692), .A2(g3172) );
  OR2_X1 OR2_185( .ZN(g6437), .A1(g6302), .A2(g6121) );
  OR2_X1 OR2_186( .ZN(g6917), .A1(g6909), .A2(g6910) );
  OR2_X1 OR2_187( .ZN(g3857), .A1(g3687), .A2(g3161) );
  OR2_X1 OR2_188( .ZN(g5533), .A1(g5351), .A2(g3290) );
  OR2_X1 OR2_189( .ZN(g5697), .A1(g5646), .A2(g5485) );
  OR2_X1 OR2_190( .ZN(g5013), .A1(g4826), .A2(g4621) );
  OR2_X1 OR2_191( .ZN(g4627), .A1(g4333), .A2(g3603) );
  OR2_X1 OR2_192( .ZN(g6454), .A1(g6344), .A2(g5949) );
  OR2_X1 OR2_193( .ZN(g6296), .A1(g6247), .A2(g6088) );
  OR2_X1 OR2_194( .ZN(g4646), .A1(g4353), .A2(g3635) );
  OR4_X1 OR4_28( .ZN(I8138), .A1(g4980), .A2(g4915), .A3(g5025), .A4(g5054) );
  OR2_X1 OR2_195( .ZN(g6189), .A1(g6060), .A2(g6035) );
  OR2_X1 OR2_196( .ZN(g3977), .A1(g3653), .A2(g3113) );
  OR4_X1 OR4_29( .ZN(I9058), .A1(g6156), .A2(g6331), .A3(g5190), .A4(g5164) );
  OR2_X1 OR2_197( .ZN(g6787), .A1(g3758), .A2(g6766) );
  OR2_X1 OR2_198( .ZN(g5060), .A1(g3491), .A2(g4819) );
  OR2_X1 OR2_199( .ZN(g6297), .A1(g6248), .A2(g6089) );
  OR2_X1 OR2_200( .ZN(g3999), .A1(g3699), .A2(g3181) );
  OR2_X2 OR2_201( .ZN(g6684), .A1(g6250), .A2(g6643) );
  OR4_X1 OR4_30( .ZN(I7978), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X2 OR2_202( .ZN(g6109), .A1(g5900), .A2(g5599) );
  OR2_X1 OR2_203( .ZN(g6791), .A1(g6768), .A2(g3307) );
  OR2_X1 OR2_204( .ZN(g6309), .A1(g6265), .A2(g6098) );
  OR2_X1 OR2_205( .ZN(g3732), .A1(g3324), .A2(g2732) );
  OR2_X1 OR2_206( .ZN(g3533), .A1(g3154), .A2(g3166) );
  OR4_X1 OR4_31( .ZN(I8385), .A1(g6316), .A2(g6128), .A3(g6131), .A4(g6149) );
  OR2_X1 OR2_207( .ZN(g6268), .A1(g5677), .A2(g5951) );
  OR2_X1 OR2_208( .ZN(g3820), .A1(g3287), .A2(g2671) );
  OR2_X1 OR2_209( .ZN(g6452), .A1(g6342), .A2(g5942) );
  OR2_X1 OR2_210( .ZN(g5626), .A1(g5496), .A2(g3285) );
  OR2_X1 OR2_211( .ZN(g4656), .A1(g4369), .A2(g3662) );
  OR2_X1 OR2_212( .ZN(g6185), .A1(g6055), .A2(g5995) );
  OR2_X1 OR2_213( .ZN(g3739), .A1(g3334), .A2(g2746) );
  OR4_X1 OR4_32( .ZN(I7989), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR2_X1 OR2_214( .ZN(g3995), .A1(g3690), .A2(g3170) );
  OR4_X1 OR4_33( .ZN(I8369), .A1(g5165), .A2(g5159), .A3(g5233), .A4(g5240) );
  OR4_X1 OR4_34( .ZN(I7971), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR2_X1 OR2_215( .ZN(g5627), .A1(g5497), .A2(g3286) );
  OR3_X1 OR3_14( .ZN(g6682), .A1(g6478), .A2(g6624), .A3(g6623) );
  OR2_X1 OR2_216( .ZN(g3942), .A1(g3215), .A2(g3575) );
  OR2_X1 OR2_217( .ZN(g5583), .A1(g5569), .A2(g4020) );
  OR2_X1 OR2_218( .ZN(g6173), .A1(g6066), .A2(g6043) );
  OR2_X1 OR2_219( .ZN(g3954), .A1(g3484), .A2(g3489) );
  OR2_X1 OR2_220( .ZN(g6920), .A1(g6915), .A2(g6916) );
  OR2_X1 OR2_221( .ZN(g6261), .A1(g5673), .A2(g5944) );
  OR2_X1 OR2_222( .ZN(g6793), .A1(g6771), .A2(g3323) );
  OR2_X1 OR2_223( .ZN(g4948), .A1(g4834), .A2(g4836) );
  OR2_X1 OR2_224( .ZN(g6246), .A1(g5665), .A2(g5937) );
  OR2_X1 OR2_225( .ZN(g5224), .A1(g5123), .A2(g3630) );
  OR2_X1 OR2_226( .ZN(g5277), .A1(g5023), .A2(g4763) );
  OR2_X1 OR2_227( .ZN(g4438), .A1(g4363), .A2(g4037) );
  OR2_X1 OR2_228( .ZN(g4773), .A1(g4495), .A2(g4220) );
  OR2_X1 OR2_229( .ZN(g6689), .A1(g6266), .A2(g6648) );
  OR2_X2 OR2_230( .ZN(g3998), .A1(g3698), .A2(g3180) );
  OR4_X1 OR4_35( .ZN(I8774), .A1(g6655), .A2(g6653), .A3(g6651), .A4(g6649) );
  OR2_X1 OR2_231( .ZN(g3850), .A1(g3680), .A2(g3145) );
  OR2_X1 OR2_232( .ZN(g6108), .A1(g5898), .A2(g5598) );
  OR3_X1 OR3_15( .ZN(g6758), .A1(g6673), .A2(g6628), .A3(g6738) );
  OR2_X1 OR2_233( .ZN(g2896), .A1(g2323), .A2(g1763) );
  OR2_X1 OR2_234( .ZN(g6455), .A1(g6345), .A2(g5952) );
  OR2_X1 OR2_235( .ZN(g3986), .A1(g3667), .A2(g3133) );
  OR2_X1 OR2_236( .ZN(g6846), .A1(g5860), .A2(g6834) );
  OR2_X1 OR2_237( .ZN(g3503), .A1(g3122), .A2(g3132) );
  OR4_X1 OR4_36( .ZN(I7969), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_238( .ZN(g4941), .A1(g4829), .A2(g4832) );
  OR2_X1 OR2_239( .ZN(g6290), .A1(g6245), .A2(g6086) );
  OR2_X1 OR2_240( .ZN(g3987), .A1(g3669), .A2(g3134) );
  OR2_X1 OR2_241( .ZN(g6847), .A1(g5861), .A2(g6837) );
  OR2_X1 OR2_242( .ZN(g6685), .A1(g6256), .A2(g6644) );
  OR2_X1 OR2_243( .ZN(g5295), .A1(g5047), .A2(g4766) );
  OR2_X1 OR2_244( .ZN(g4473), .A1(g3575), .A2(g4253) );
  OR2_X1 OR2_245( .ZN(g3991), .A1(g3685), .A2(g3156) );
  OR4_X1 OR4_37( .ZN(I7988), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_246( .ZN(g5471), .A1(g5360), .A2(g5143) );
  OR4_X1 OR4_38( .ZN(I8368), .A1(g6148), .A2(g6321), .A3(g5176), .A4(g5184) );
  OR2_X1 OR2_247( .ZN(g6257), .A1(g5671), .A2(g5941) );
  OR2_X1 OR2_248( .ZN(g6301), .A1(g6254), .A2(g6092) );
  OR4_X1 OR4_39( .ZN(g6673), .A1(g6559), .A2(g6640), .A3(g4416), .A4(g2950) );
  OR4_X1 OR4_40( .ZN(I8080), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_249( .ZN(g6669), .A1(g6613), .A2(g4679) );
  OR2_X1 OR2_250( .ZN(g3877), .A1(g3651), .A2(g3659) );
  OR4_X1 OR4_41( .ZN(I8126), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_251( .ZN(g5062), .A1(g4661), .A2(g4666) );
  OR2_X1 OR2_252( .ZN(g6480), .A1(I8360), .A2(g6359) );
  OR4_X2 OR4_42( .ZN(I8779), .A1(g6605), .A2(g6656), .A3(g6654), .A4(g6652) );
  OR2_X1 OR2_253( .ZN(g6688), .A1(g6263), .A2(g6647) );
  OR2_X1 OR2_254( .ZN(g5085), .A1(g4694), .A2(g4280) );
  OR2_X1 OR2_255( .ZN(I7981), .A1(g4915), .A2(g5025) );
  OR4_X1 OR4_43( .ZN(I8127), .A1(g6015), .A2(g6212), .A3(g4950), .A4(g4877) );
  OR2_X1 OR2_256( .ZN(g4433), .A1(g4354), .A2(g4032) );
  OR4_X1 OR4_44( .ZN(I8346), .A1(g6159), .A2(g6334), .A3(g5163), .A4(g5191) );
  OR2_X1 OR2_257( .ZN(g5812), .A1(g5376), .A2(g5618) );
  OR2_X1 OR2_258( .ZN(g4859), .A1(g4730), .A2(g4486) );
  OR2_X1 OR2_259( .ZN(g6665), .A1(I8778), .A2(I8779) );
  OR2_X1 OR2_260( .ZN(g5473), .A1(g5362), .A2(g5145) );
  OR4_X1 OR4_45( .ZN(I8347), .A1(g5188), .A2(g5157), .A3(g5154), .A4(g5193) );
  OR2_X1 OR2_261( .ZN(g6303), .A1(g6258), .A2(g6094) );
  OR2_X1 OR2_262( .ZN(g5069), .A1(g1595), .A2(g4688) );
  OR4_X1 OR4_46( .ZN(I9064), .A1(g6323), .A2(g6829), .A3(g6831), .A4(g6155) );
  OR2_X1 OR2_263( .ZN(g4497), .A1(g4166), .A2(g3784) );
  OR4_X1 OR4_47( .ZN(I8210), .A1(g5202), .A2(g4993), .A3(g4967), .A4(g4980) );
  OR2_X1 OR2_264( .ZN(g5377), .A1(g5217), .A2(g4949) );
  OR2_X1 OR2_265( .ZN(g3837), .A1(g3609), .A2(g3613) );
  OR2_X1 OR2_266( .ZN(g6116), .A1(g5910), .A2(g5617) );
  OR4_X1 OR4_48( .ZN(I8117), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_267( .ZN(g4001), .A1(g3702), .A2(g3190) );
  OR2_X2 OR2_268( .ZN(g3842), .A1(g3670), .A2(g3135) );
  OR2_X1 OR2_269( .ZN(g5291), .A1(g5043), .A2(g4764) );
  OR2_X1 OR2_270( .ZN(g3941), .A1(g3479), .A2(g2873) );
  OR2_X1 OR2_271( .ZN(g5694), .A1(g5633), .A2(g5482) );
  OR2_X1 OR2_272( .ZN(g6936), .A1(g5438), .A2(g6935) );
  OR2_X1 OR2_273( .ZN(g4068), .A1(g3293), .A2(g2685) );
  OR4_X1 OR4_49( .ZN(I8079), .A1(g6194), .A2(g5958), .A3(g5975), .A4(g5997) );
  OR2_X1 OR2_274( .ZN(g4468), .A1(g4214), .A2(g3831) );
  OR2_X1 OR2_275( .ZN(g4866), .A1(g4756), .A2(g4491) );
  OR2_X1 OR2_276( .ZN(g3829), .A1(g3294), .A2(g3305) );
  OR4_X1 OR4_50( .ZN(I8356), .A1(g6311), .A2(g6123), .A3(g6125), .A4(g6141) );
  OR2_X1 OR2_277( .ZN(g3733), .A1(g3325), .A2(g2733) );
  OR2_X1 OR2_278( .ZN(g6937), .A1(g4616), .A2(g6934) );
  OR2_X1 OR2_279( .ZN(g6479), .A1(I8349), .A2(g6335) );
  OR2_X1 OR2_280( .ZN(g6294), .A1(g6249), .A2(g6090) );
  OR2_X1 OR2_281( .ZN(g5065), .A1(g4667), .A2(g4671) );
  OR2_X1 OR2_282( .ZN(g5228), .A1(g5096), .A2(g4800) );
  OR4_X1 OR4_51( .ZN(I8357), .A1(g6145), .A2(g6318), .A3(g5171), .A4(g5187) );
  OR2_X1 OR2_283( .ZN(g3849), .A1(g3618), .A2(g3625) );
  OR2_X1 OR2_284( .ZN(g6704), .A1(g6660), .A2(g492) );
  OR2_X1 OR2_285( .ZN(g4599), .A1(g3499), .A2(g4230) );
  OR2_X1 OR2_286( .ZN(g6453), .A1(g6343), .A2(g5945) );
  OR2_X1 OR2_287( .ZN(g4544), .A1(g4410), .A2(g2995) );
  OR4_X1 OR4_52( .ZN(I8778), .A1(g6612), .A2(g6611), .A3(g6609), .A4(g6607) );
  OR2_X1 OR2_288( .ZN(g2924), .A1(g2095), .A2(g1573) );
  OR2_X1 OR2_289( .ZN(g4427), .A1(g4373), .A2(g3668) );
  OR2_X1 OR2_290( .ZN(g4446), .A1(g4383), .A2(g4043) );
  OR2_X1 OR2_291( .ZN(g3870), .A1(g3700), .A2(g3182) );
  OR3_X1 OR3_16( .ZN(g6683), .A1(g6465), .A2(g6622), .A3(g6621) );
  OR2_X1 OR2_292( .ZN(g5676), .A1(g5559), .A2(g5424) );
  OR2_X1 OR2_293( .ZN(g4637), .A1(g4344), .A2(g3619) );
  OR2_X1 OR2_294( .ZN(g3972), .A1(g3646), .A2(g3103) );
  OR2_X1 OR2_295( .ZN(g6782), .A1(g6719), .A2(g6749) );
  OR2_X1 OR2_296( .ZN(g6661), .A1(I8773), .A2(I8774) );
  OR2_X2 OR2_297( .ZN(g4757), .A1(g4456), .A2(g4158) );
  OR2_X2 OR2_298( .ZN(g6292), .A1(g6243), .A2(g6084) );
  OR2_X1 OR2_299( .ZN(g4811), .A1(g4429), .A2(g4432) );
  OR2_X1 OR2_300( .ZN(g4642), .A1(g4348), .A2(g3628) );
  OR2_X1 OR2_301( .ZN(g4447), .A1(g4384), .A2(g4044) );
  OR2_X1 OR2_302( .ZN(g5624), .A1(g5494), .A2(g3280) );
  OR2_X1 OR2_303( .ZN(g5068), .A1(g4673), .A2(g4677) );
  OR2_X1 OR2_304( .ZN(g4654), .A1(g4362), .A2(g3654) );
  OR2_X1 OR2_305( .ZN(g3891), .A1(g3683), .A2(g3688) );
  OR2_X1 OR2_306( .ZN(g3913), .A1(g3449), .A2(g2860) );
  OR2_X1 OR2_307( .ZN(I7990), .A1(g4915), .A2(g5025) );
  OR2_X1 OR2_308( .ZN(g6702), .A1(g6659), .A2(g496) );
  OR2_X1 OR2_309( .ZN(g6919), .A1(g6912), .A2(g6914) );
  OR2_X1 OR2_310( .ZN(I8120), .A1(g4915), .A2(g5025) );
  OR2_X1 OR2_311( .ZN(g4243), .A1(g4053), .A2(g4058) );
  OR2_X1 OR2_312( .ZN(g5699), .A1(g5660), .A2(g5487) );
  OR2_X1 OR2_313( .ZN(g5241), .A1(g5069), .A2(g2067) );
  OR2_X1 OR2_314( .ZN(g4234), .A1(g3921), .A2(g478) );
  OR2_X1 OR2_315( .ZN(g3815), .A1(g3282), .A2(g2659) );
  OR2_X1 OR2_316( .ZN(g5386), .A1(g5227), .A2(g669) );
  OR2_X1 OR2_317( .ZN(g6789), .A1(g3764), .A2(g6769) );
  OR4_X1 OR4_53( .ZN(I8082), .A1(g4980), .A2(g4915), .A3(g5025), .A4(g5054) );
  OR2_X1 OR2_318( .ZN(g5370), .A1(g5211), .A2(g4937) );
  OR2_X2 OR2_319( .ZN(g3828), .A1(g3304), .A2(g1351) );
  OR4_X1 OR4_54( .ZN(I9065), .A1(g6158), .A2(g6333), .A3(g5152), .A4(g5156) );
  OR2_X1 OR2_320( .ZN(g3746), .A1(g3357), .A2(g2771) );
  OR2_X1 OR2_321( .ZN(g5083), .A1(g4688), .A2(g4271) );
  OR2_X1 OR2_322( .ZN(g6907), .A1(g6874), .A2(g3358) );
  OR2_X1 OR2_323( .ZN(g5622), .A1(g5492), .A2(g3277) );
  OR2_X1 OR2_324( .ZN(g6690), .A1(g6270), .A2(g6650) );
  OR4_X1 OR4_55( .ZN(g6482), .A1(I8376), .A2(I8377), .A3(I8378), .A4(I8379) );
  OR2_X1 OR2_325( .ZN(g4652), .A1(g4358), .A2(g3645) );
  OR2_X1 OR2_326( .ZN(g4549), .A1(g4416), .A2(g3013) );
  OR2_X1 OR2_327( .ZN(g3747), .A1(g3365), .A2(g2781) );
  OR2_X1 OR2_328( .ZN(g3855), .A1(g3626), .A2(g3631) );
  OR2_X1 OR2_329( .ZN(g5695), .A1(g5635), .A2(g5483) );
  OR2_X1 OR2_330( .ZN(g6110), .A1(g5883), .A2(g5996) );
  OR2_X1 OR2_331( .ZN(g6310), .A1(g6269), .A2(g6099) );
  OR2_X1 OR2_332( .ZN(g5016), .A1(g4789), .A2(g4592) );
  OR3_X1 OR3_17( .ZN(g6762), .A1(g6679), .A2(g6628), .A3(g6739) );
  OR2_X1 OR2_333( .ZN(g4740), .A1(g4448), .A2(g4154) );
  OR4_X1 OR4_56( .ZN(I8394), .A1(g6154), .A2(g6329), .A3(g5186), .A4(g5172) );
  OR2_X1 OR2_334( .ZN(g6556), .A1(g6339), .A2(g6467) );
  OR2_X1 OR2_335( .ZN(g6930), .A1(g6740), .A2(g6928) );
  OR2_X1 OR2_336( .ZN(g3599), .A1(g2935), .A2(g1637) );
  OR2_X2 OR2_337( .ZN(g3821), .A1(g2951), .A2(g3466) );
  OR2_X1 OR2_338( .ZN(g4860), .A1(g4735), .A2(g4488) );
  OR2_X1 OR2_339( .ZN(g6237), .A1(g5912), .A2(g2381) );
  OR2_X1 OR2_340( .ZN(g4645), .A1(g4352), .A2(g3633) );
  OR3_X2 OR3_18( .ZN(g6844), .A1(I9057), .A2(I9058), .A3(I9059) );
  OR4_X2 OR4_57( .ZN(I8773), .A1(g6610), .A2(g6608), .A3(g6606), .A4(g6604) );
  OR2_X1 OR2_341( .ZN(g5629), .A1(g5499), .A2(g3298) );
  OR2_X1 OR2_342( .ZN(g4607), .A1(g4232), .A2(g3899) );
  OR2_X1 OR2_343( .ZN(g6705), .A1(g6693), .A2(g4835) );
  OR2_X1 OR2_344( .ZN(g5800), .A1(g5369), .A2(g5600) );
  OR2_X1 OR2_345( .ZN(g6242), .A1(g2356), .A2(g6075) );
  OR2_X1 OR2_346( .ZN(g3841), .A1(g3614), .A2(g3617) );
  OR2_X1 OR2_347( .ZN(g6918), .A1(g6911), .A2(g6913) );
  OR2_X1 OR2_348( .ZN(g5348), .A1(g5317), .A2(g5122) );
  OR2_X1 OR2_349( .ZN(g3858), .A1(g3629), .A2(g3636) );
  OR2_X1 OR2_350( .ZN(g5698), .A1(g5648), .A2(g5486) );
  OR2_X1 OR2_351( .ZN(g4630), .A1(g4339), .A2(g3610) );
  OR2_X1 OR2_352( .ZN(g6921), .A1(g6908), .A2(g6816) );
  OR2_X1 OR2_353( .ZN(g5367), .A1(g5199), .A2(g4928) );
  NAND3_X1 NAND3_0( .ZN(g1777), .A1(g1060), .A2(g102), .A3(g89) );
  NAND2_X2 NAND2_0( .ZN(I7217), .A1(g152), .A2(I7216) );
  NAND2_X1 NAND2_1( .ZN(I7571), .A1(g5678), .A2(I7569) );
  NAND4_X4 NAND4_0( .ZN(g5686), .A1(g5546), .A2(g1017), .A3(g1551), .A4(g2916) );
  NAND2_X1 NAND2_2( .ZN(I2073), .A1(g15), .A2(I2072) );
  NAND2_X1 NAND2_3( .ZN(I2796), .A1(g804), .A2(I2795) );
  NAND2_X1 NAND2_4( .ZN(g948), .A1(I2014), .A2(I2015) );
  NAND2_X1 NAND2_5( .ZN(I4205), .A1(g743), .A2(I4203) );
  NAND2_X1 NAND2_6( .ZN(I3875), .A1(g285), .A2(I3874) );
  NAND3_X1 NAND3_1( .ZN(g3330), .A1(g1815), .A2(g1797), .A3(g3109) );
  NAND2_X1 NAND2_7( .ZN(g4151), .A1(I5536), .A2(I5537) );
  NAND3_X2 NAND3_2( .ZN(g2435), .A1(g1138), .A2(g1777), .A3(g1157) );
  NAND2_X1 NAND2_8( .ZN(I5658), .A1(g3983), .A2(I5657) );
  NAND2_X1 NAND2_9( .ZN(g1558), .A1(I2527), .A2(I2528) );
  NAND2_X1 NAND2_10( .ZN(I4444), .A1(g2092), .A2(g606) );
  NAND2_X1 NAND2_11( .ZN(I5271), .A1(g3710), .A2(I5269) );
  NAND2_X1 NAND2_12( .ZN(I2898), .A1(g1027), .A2(I2897) );
  NAND2_X1 NAND2_13( .ZN(I2797), .A1(g798), .A2(I2795) );
  NAND2_X1 NAND2_14( .ZN(I2245), .A1(g567), .A2(I2244) );
  NAND2_X1 NAND2_15( .ZN(I3988), .A1(g291), .A2(g2544) );
  NAND2_X1 NAND2_16( .ZN(g1574), .A1(I2543), .A2(I2544) );
  NAND4_X1 NAND4_1( .ZN(g3529), .A1(g3200), .A2(g2215), .A3(g2976), .A4(g2968) );
  NAND2_X1 NAND2_17( .ZN(I1963), .A1(g242), .A2(I1961) );
  NAND2_X1 NAND2_18( .ZN(I5209), .A1(g3271), .A2(I5207) );
  NAND2_X1 NAND2_19( .ZN(I7562), .A1(g74), .A2(g5676) );
  NAND2_X1 NAND2_20( .ZN(g5506), .A1(I7231), .A2(I7232) );
  NAND2_X1 NAND2_21( .ZN(g5111), .A1(I6744), .A2(I6745) );
  NAND2_X1 NAND2_22( .ZN(I4182), .A1(g2292), .A2(g749) );
  NAND2_X1 NAND2_23( .ZN(I6186), .A1(g4301), .A2(I6185) );
  NAND2_X1 NAND2_24( .ZN(I7441), .A1(g594), .A2(I7439) );
  NAND2_X1 NAND2_25( .ZN(I6026), .A1(g4223), .A2(g4221) );
  NAND2_X1 NAND2_26( .ZN(I2768), .A1(g743), .A2(I2766) );
  NAND2_X1 NAND2_27( .ZN(I3933), .A1(g288), .A2(g2473) );
  NAND3_X1 NAND3_3( .ZN(g5853), .A1(g5638), .A2(g2053), .A3(g1076) );
  NAND2_X1 NAND2_28( .ZN(g2731), .A1(I3894), .A2(I3895) );
  NAND2_X1 NAND2_29( .ZN(g5507), .A1(I7238), .A2(I7239) );
  NAND2_X1 NAND2_30( .ZN(g2966), .A1(I4160), .A2(I4161) );
  NAND2_X1 NAND2_31( .ZN(I2934), .A1(g1436), .A2(I2933) );
  NAND2_X1 NAND2_32( .ZN(I3179), .A1(g736), .A2(I3177) );
  NAND2_X1 NAND2_33( .ZN(I6187), .A1(g3955), .A2(I6185) );
  NAND2_X1 NAND2_34( .ZN(I6027), .A1(g4223), .A2(I6026) );
  NAND3_X2 NAND3_4( .ZN(g2009), .A1(g901), .A2(g1387), .A3(g905) );
  NAND2_X1 NAND2_35( .ZN(I4233), .A1(g2267), .A2(g798) );
  NAND2_X1 NAND2_36( .ZN(g2769), .A1(I3953), .A2(I3954) );
  NAND2_X1 NAND2_37( .ZN(g1044), .A1(I2081), .A2(I2082) );
  NAND4_X1 NAND4_2( .ZN(g4674), .A1(g4550), .A2(g1514), .A3(g2107), .A4(g2897) );
  NAND2_X1 NAND2_38( .ZN(I7569), .A1(g79), .A2(g5678) );
  NAND2_X1 NAND2_39( .ZN(I6391), .A1(g4504), .A2(I6390) );
  NAND4_X1 NAND4_3( .ZN(g3525), .A1(g3192), .A2(g3002), .A3(g2197), .A4(g2179) );
  NAND4_X1 NAND4_4( .ZN(g4680), .A1(g4550), .A2(g1514), .A3(g1006), .A4(g2897) );
  NAND2_X1 NAND2_40( .ZN(I2081), .A1(g25), .A2(I2080) );
  NAND2_X1 NAND2_41( .ZN(I8195), .A1(g471), .A2(I8194) );
  NAND2_X1 NAND2_42( .ZN(g1534), .A1(I2498), .A2(I2499) );
  NAND2_X1 NAND2_43( .ZN(I2497), .A1(g1042), .A2(g1036) );
  NAND2_X1 NAND2_44( .ZN(g939), .A1(I1987), .A2(I1988) );
  NAND2_X1 NAND2_45( .ZN(I5269), .A1(g3705), .A2(g3710) );
  NAND3_X2 NAND3_5( .ZN(g3985), .A1(g1138), .A2(g3718), .A3(g2142) );
  NAND2_X1 NAND2_46( .ZN(g1036), .A1(I2061), .A2(I2062) );
  NAND2_X1 NAND2_47( .ZN(I2676), .A1(g131), .A2(I2674) );
  NAND2_X1 NAND2_48( .ZN(g1749), .A1(I2767), .A2(I2768) );
  NAND2_X1 NAND2_49( .ZN(g6097), .A1(g2954), .A2(g5857) );
  NAND3_X1 NAND3_6( .ZN(g6783), .A1(g6747), .A2(g5068), .A3(g5066) );
  NAND2_X1 NAND2_50( .ZN(g5776), .A1(I7528), .A2(I7529) );
  NAND2_X1 NAND2_51( .ZN(I7434), .A1(g5554), .A2(I7432) );
  NAND2_X1 NAND2_52( .ZN(g1042), .A1(I2073), .A2(I2074) );
  NAND2_X1 NAND2_53( .ZN(I7210), .A1(g5367), .A2(I7208) );
  NAND4_X1 NAND4_5( .ZN(g3530), .A1(g3204), .A2(g3023), .A3(g2197), .A4(g2179) );
  NAND2_X1 NAND2_54( .ZN(I6964), .A1(g586), .A2(I6962) );
  NAND2_X1 NAND2_55( .ZN(I5208), .A1(g3267), .A2(I5207) );
  NAND2_X1 NAND2_56( .ZN(I5302), .A1(g3505), .A2(I5300) );
  NAND2_X1 NAND2_57( .ZN(g5777), .A1(I7535), .A2(I7536) );
  NAND2_X1 NAND2_58( .ZN(g4613), .A1(I6195), .A2(I6196) );
  NAND2_X1 NAND2_59( .ZN(I2544), .A1(g774), .A2(I2542) );
  NAND2_X1 NAND2_60( .ZN(g1138), .A1(g102), .A2(g98) );
  NAND2_X1 NAND2_61( .ZN(I1994), .A1(g504), .A2(g218) );
  NAND2_X1 NAND2_62( .ZN(I4445), .A1(g2092), .A2(I4444) );
  NAND2_X1 NAND2_63( .ZN(I2061), .A1(g7), .A2(I2060) );
  NAND2_X1 NAND2_64( .ZN(I5189), .A1(g3593), .A2(I5187) );
  NAND2_X1 NAND2_65( .ZN(g4903), .A1(g4717), .A2(g858) );
  NAND2_X1 NAND2_66( .ZN(I3178), .A1(g1706), .A2(I3177) );
  NAND2_X1 NAND2_67( .ZN(I4920), .A1(g3522), .A2(I4919) );
  NAND2_X1 NAND2_68( .ZN(g2951), .A1(g2142), .A2(g1797) );
  NAND4_X1 NAND4_6( .ZN(g3518), .A1(g3177), .A2(g3023), .A3(g3007), .A4(g2981) );
  NAND2_X1 NAND2_69( .ZN(I2003), .A1(g500), .A2(g212) );
  NAND3_X2 NAND3_7( .ZN(g6717), .A1(g6669), .A2(g5065), .A3(g5062) );
  NAND2_X1 NAND2_70( .ZN(I3916), .A1(g2449), .A2(I3914) );
  NAND4_X1 NAND4_7( .ZN(g5864), .A1(g5649), .A2(g1529), .A3(g1088), .A4(g2068) );
  NAND3_X1 NAND3_8( .ZN(g2008), .A1(g866), .A2(g873), .A3(g1784) );
  NAND2_X1 NAND2_71( .ZN(I5309), .A1(g3512), .A2(I5307) );
  NAND2_X1 NAND2_72( .ZN(I7432), .A1(g111), .A2(g5554) );
  NAND2_X1 NAND2_73( .ZN(I4203), .A1(g2255), .A2(g743) );
  NAND4_X1 NAND4_8( .ZN(g3521), .A1(g3187), .A2(g3023), .A3(g3007), .A4(g2179) );
  NAND2_X1 NAND2_74( .ZN(I5759), .A1(g3836), .A2(g3503) );
  NAND2_X1 NAND2_75( .ZN(I6962), .A1(g4874), .A2(g586) );
  NAND2_X1 NAND2_76( .ZN(I6659), .A1(g4762), .A2(g3541) );
  NAND2_X1 NAND2_77( .ZN(I4940), .A1(g3437), .A2(I4939) );
  NAND2_X1 NAND2_78( .ZN(I2935), .A1(g345), .A2(I2933) );
  NAND2_X1 NAND2_79( .ZN(g2266), .A1(I3412), .A2(I3413) );
  NAND2_X1 NAND2_80( .ZN(I2542), .A1(g821), .A2(g774) );
  NAND2_X1 NAND2_81( .ZN(I3412), .A1(g1419), .A2(I3411) );
  NAND2_X1 NAND2_82( .ZN(I3189), .A1(g1716), .A2(I3188) );
  NAND2_X1 NAND2_83( .ZN(g5634), .A1(g5563), .A2(g4767) );
  NAND2_X1 NAND2_84( .ZN(I3990), .A1(g2544), .A2(I3988) );
  NAND2_X1 NAND2_85( .ZN(g2960), .A1(I4151), .A2(I4152) );
  NAND2_X1 NAND2_86( .ZN(g5926), .A1(g5741), .A2(g639) );
  NAND4_X1 NAND4_9( .ZN(g3511), .A1(g3158), .A2(g3002), .A3(g2976), .A4(g2968) );
  NAND2_X1 NAND2_87( .ZN(I7439), .A1(g5515), .A2(g594) );
  NAND2_X1 NAND2_88( .ZN(I2090), .A1(g33), .A2(I2089) );
  NAND4_X1 NAND4_10( .ZN(g5862), .A1(g5649), .A2(g1529), .A3(g1535), .A4(g2068) );
  NAND2_X1 NAND2_89( .ZN(I9050), .A1(g6832), .A2(g3598) );
  NAND2_X1 NAND2_90( .ZN(I5766), .A1(g3961), .A2(g3957) );
  NAND3_X1 NAND3_9( .ZN(g1582), .A1(g784), .A2(g774), .A3(g821) );
  NAND2_X1 NAND2_91( .ZN(g1793), .A1(g94), .A2(g1084) );
  NAND2_X1 NAND2_92( .ZN(g3968), .A1(I5227), .A2(I5228) );
  NAND2_X1 NAND2_93( .ZN(I7527), .A1(g49), .A2(g5662) );
  NAND2_X1 NAND2_94( .ZN(I5226), .A1(g3259), .A2(g3263) );
  NAND2_X1 NAND2_95( .ZN(g4049), .A1(g3677), .A2(g3425) );
  NAND2_X1 NAND2_96( .ZN(I7224), .A1(g161), .A2(I7223) );
  NAND2_X1 NAND2_97( .ZN(I5767), .A1(g3961), .A2(I5766) );
  NAND2_X1 NAND2_98( .ZN(I5535), .A1(g3907), .A2(g654) );
  NAND2_X1 NAND2_99( .ZN(I5227), .A1(g3259), .A2(I5226) );
  NAND2_X1 NAND2_100( .ZN(g5947), .A1(g5821), .A2(g2944) );
  NAND2_X1 NAND2_101( .ZN(g3742), .A1(I4920), .A2(I4921) );
  NAND4_X2 NAND4_11( .ZN(g5873), .A1(g5649), .A2(g1017), .A3(g1564), .A4(g2113) );
  NAND2_X1 NAND2_102( .ZN(g4504), .A1(I6027), .A2(I6028) );
  NAND2_X1 NAND2_103( .ZN(I7244), .A1(g188), .A2(g5377) );
  NAND3_X1 NAND3_10( .ZN(g5869), .A1(g5649), .A2(g1076), .A3(g2081) );
  NAND2_X1 NAND2_104( .ZN(I5188), .A1(g3589), .A2(I5187) );
  NAND2_X1 NAND2_105( .ZN(g3983), .A1(I5270), .A2(I5271) );
  NAND4_X1 NAND4_12( .ZN(g4678), .A1(g2897), .A2(g2101), .A3(g1514), .A4(g4550) );
  NAND2_X1 NAND2_106( .ZN(g6843), .A1(I9051), .A2(I9052) );
  NAND2_X1 NAND2_107( .ZN(g3961), .A1(I5208), .A2(I5209) );
  NAND2_X1 NAND2_108( .ZN(I5308), .A1(g478), .A2(I5307) );
  NAND2_X1 NAND2_109( .ZN(I2506), .A1(g1047), .A2(g1044) );
  NAND2_X1 NAND2_110( .ZN(I3445), .A1(g1689), .A2(g729) );
  NAND2_X1 NAND2_111( .ZN(g2061), .A1(I3169), .A2(I3170) );
  NAND2_X1 NAND2_112( .ZN(I3169), .A1(g1540), .A2(I3168) );
  NAND3_X1 NAND3_11( .ZN(g6740), .A1(g6703), .A2(g6457), .A3(g4936) );
  NAND2_X1 NAND2_113( .ZN(I7556), .A1(g69), .A2(I7555) );
  NAND2_X1 NAND2_114( .ZN(g4007), .A1(I5308), .A2(I5309) );
  NAND2_X1 NAND2_115( .ZN(I5196), .A1(g3567), .A2(I5195) );
  NAND2_X1 NAND2_116( .ZN(I7563), .A1(g74), .A2(I7562) );
  NAND2_X1 NAND2_117( .ZN(g5684), .A1(I7440), .A2(I7441) );
  NAND2_X1 NAND2_118( .ZN(I2507), .A1(g1047), .A2(I2506) );
  NAND2_X1 NAND2_119( .ZN(I1995), .A1(g504), .A2(I1994) );
  NAND2_X1 NAND2_120( .ZN(g2307), .A1(I3446), .A2(I3447) );
  NAND2_X1 NAND2_121( .ZN(I7237), .A1(g179), .A2(g5374) );
  NAND2_X1 NAND2_122( .ZN(g2858), .A1(g1815), .A2(g2577) );
  NAND2_X1 NAND2_123( .ZN(g2757), .A1(I3934), .A2(I3935) );
  NAND2_X1 NAND2_124( .ZN(I6744), .A1(g4708), .A2(I6743) );
  NAND2_X1 NAND2_125( .ZN(I4183), .A1(g2292), .A2(I4182) );
  NAND2_X1 NAND2_126( .ZN(I7557), .A1(g5674), .A2(I7555) );
  NAND2_X1 NAND2_127( .ZN(I2300), .A1(g830), .A2(I2299) );
  NAND2_X1 NAND2_128( .ZN(I3188), .A1(g1716), .A2(g791) );
  NAND4_X1 NAND4_13( .ZN(g5865), .A1(g5649), .A2(g1088), .A3(g1076), .A4(g2068) );
  NAND2_X1 NAND2_129( .ZN(I5197), .A1(g3571), .A2(I5195) );
  NAND2_X1 NAND2_130( .ZN(I4161), .A1(g619), .A2(I4159) );
  NAND2_X1 NAND2_131( .ZN(I3741), .A1(g349), .A2(I3739) );
  NAND2_X1 NAND2_132( .ZN(g5019), .A1(I6660), .A2(I6661) );
  NAND2_X1 NAND2_133( .ZN(I5257), .A1(g3714), .A2(g3719) );
  NAND4_X1 NAND4_14( .ZN(g3532), .A1(g3212), .A2(g2215), .A3(g3007), .A4(g2981) );
  NAND2_X1 NAND2_134( .ZN(I2528), .A1(g719), .A2(I2526) );
  NAND2_X1 NAND2_135( .ZN(I5301), .A1(g471), .A2(I5300) );
  NAND2_X1 NAND2_136( .ZN(g1743), .A1(g1064), .A2(g94) );
  NAND2_X1 NAND2_137( .ZN(g1411), .A1(g314), .A2(g873) );
  NAND2_X1 NAND2_138( .ZN(g3012), .A1(I4204), .A2(I4205) );
  NAND2_X1 NAND2_139( .ZN(g5504), .A1(I7217), .A2(I7218) );
  NAND2_X1 NAND2_140( .ZN(I6175), .A1(g4236), .A2(g571) );
  NAND2_X1 NAND2_141( .ZN(I3455), .A1(g1691), .A2(g784) );
  NAND2_X1 NAND2_142( .ZN(I6500), .A1(g4504), .A2(I6499) );
  NAND3_X2 NAND3_12( .ZN(g1573), .A1(g729), .A2(g719), .A3(g766) );
  NAND2_X1 NAND2_143( .ZN(I3846), .A1(g284), .A2(g2370) );
  NAND2_X1 NAND2_144( .ZN(I4210), .A1(g2294), .A2(g804) );
  NAND2_X1 NAND2_145( .ZN(g4803), .A1(I6474), .A2(I6475) );
  NAND2_X1 NAND2_146( .ZN(g3109), .A1(g2360), .A2(g1064) );
  NAND2_X1 NAND2_147( .ZN(g2698), .A1(I3847), .A2(I3848) );
  NAND2_X1 NAND2_148( .ZN(g3957), .A1(I5196), .A2(I5197) );
  NAND2_X1 NAND2_149( .ZN(I6499), .A1(g4504), .A2(g3541) );
  NAND4_X1 NAND4_15( .ZN(g4816), .A1(g996), .A2(g4550), .A3(g1518), .A4(g2073) );
  NAND2_X1 NAND2_150( .ZN(I3847), .A1(g284), .A2(I3846) );
  NAND2_X1 NAND2_151( .ZN(I7520), .A1(g361), .A2(g5659) );
  NAND2_X1 NAND2_152( .ZN(I4784), .A1(g622), .A2(I4782) );
  NAND2_X1 NAND2_153( .ZN(I1952), .A1(g524), .A2(I1951) );
  NAND4_X1 NAND4_16( .ZN(g3539), .A1(g2591), .A2(g2215), .A3(g2197), .A4(g2981) );
  NAND2_X1 NAND2_154( .ZN(I8202), .A1(g478), .A2(I8201) );
  NAND2_X1 NAND2_155( .ZN(I1986), .A1(g508), .A2(g224) );
  NAND2_X1 NAND2_156( .ZN(I2933), .A1(g1436), .A2(g345) );
  NAND2_X1 NAND2_157( .ZN(I5760), .A1(g3836), .A2(I5759) );
  NAND2_X2 NAND2_158( .ZN(g4301), .A1(I5767), .A2(I5768) );
  NAND2_X2 NAND2_159( .ZN(I1970), .A1(g516), .A2(I1969) );
  NAND2_X2 NAND2_160( .ZN(I7225), .A1(g5370), .A2(I7223) );
  NAND2_X2 NAND2_161( .ZN(I6660), .A1(g4762), .A2(I6659) );
  NAND2_X2 NAND2_162( .ZN(g5502), .A1(I7209), .A2(I7210) );
  NAND2_X2 NAND2_163( .ZN(I3168), .A1(g1540), .A2(g1534) );
  NAND2_X2 NAND2_164( .ZN(I1987), .A1(g508), .A2(I1986) );
  NAND2_X2 NAND2_165( .ZN(g1316), .A1(I2300), .A2(I2301) );
  NAND2_X1 NAND2_166( .ZN(I2674), .A1(g710), .A2(g131) );
  NAND4_X1 NAND4_17( .ZN(g4669), .A1(g4550), .A2(g1017), .A3(g1680), .A4(g2897) );
  NAND2_X1 NAND2_167( .ZN(I3411), .A1(g1419), .A2(g616) );
  NAND2_X1 NAND2_168( .ZN(I7245), .A1(g188), .A2(I7244) );
  NAND2_X1 NAND2_169( .ZN(g2607), .A1(I3740), .A2(I3741) );
  NAND2_X1 NAND2_170( .ZN(g5308), .A1(I6963), .A2(I6964) );
  NAND2_X1 NAND2_171( .ZN(g2311), .A1(I3456), .A2(I3457) );
  NAND4_X1 NAND4_18( .ZN(g3535), .A1(g3216), .A2(g2215), .A3(g2197), .A4(g2968) );
  NAND2_X1 NAND2_172( .ZN(g5455), .A1(g2330), .A2(g5311) );
  NAND2_X1 NAND2_173( .ZN(I4782), .A1(g2846), .A2(g622) );
  NAND2_X1 NAND2_174( .ZN(I9052), .A1(g3598), .A2(I9050) );
  NAND2_X1 NAND2_175( .ZN(I3126), .A1(g1279), .A2(I3125) );
  NAND2_X1 NAND2_176( .ZN(I3400), .A1(g135), .A2(I3398) );
  NAND2_X1 NAND2_177( .ZN(I4526), .A1(g2909), .A2(g646) );
  NAND2_X1 NAND2_178( .ZN(g5780), .A1(I7556), .A2(I7557) );
  NAND2_X1 NAND2_179( .ZN(g3246), .A1(I4527), .A2(I4528) );
  NAND3_X2 NAND3_13( .ZN(g3502), .A1(g1411), .A2(g1402), .A3(g2795) );
  NAND2_X1 NAND2_180( .ZN(g4608), .A1(I6176), .A2(I6177) );
  NAND2_X1 NAND2_181( .ZN(I4919), .A1(g3522), .A2(g650) );
  NAND3_X1 NAND3_14( .ZN(g2100), .A1(g1588), .A2(g804), .A3(g791) );
  NAND2_X1 NAND2_182( .ZN(I7230), .A1(g170), .A2(g5372) );
  NAND2_X1 NAND2_183( .ZN(I7433), .A1(g111), .A2(I7432) );
  NAND2_X1 NAND2_184( .ZN(I3127), .A1(g1276), .A2(I3125) );
  NAND2_X1 NAND2_185( .ZN(g3028), .A1(I4234), .A2(I4235) );
  NAND2_X1 NAND2_186( .ZN(I2795), .A1(g804), .A2(g798) );
  NAND2_X1 NAND2_187( .ZN(I5784), .A1(g628), .A2(I5782) );
  NAND2_X1 NAND2_188( .ZN(I4527), .A1(g2909), .A2(I4526) );
  NAND2_X1 NAND2_189( .ZN(I7550), .A1(g5672), .A2(I7548) );
  NAND2_X1 NAND2_190( .ZN(I4546), .A1(g2853), .A2(I4545) );
  NAND2_X1 NAND2_191( .ZN(I6745), .A1(g582), .A2(I6743) );
  NAND2_X1 NAND2_192( .ZN(I5294), .A1(g625), .A2(I5292) );
  NAND2_X1 NAND2_193( .ZN(I6963), .A1(g4874), .A2(I6962) );
  NAND3_X1 NAND3_15( .ZN(g3741), .A1(g901), .A2(g3433), .A3(g2340) );
  NAND2_X1 NAND2_194( .ZN(g1157), .A1(g89), .A2(g107) );
  NAND2_X1 NAND2_195( .ZN(I2499), .A1(g1036), .A2(I2497) );
  NAND2_X1 NAND2_196( .ZN(g937), .A1(I1979), .A2(I1980) );
  NAND2_X1 NAND2_197( .ZN(g4472), .A1(g3380), .A2(g4253) );
  NAND3_X1 NAND3_16( .ZN(g2010), .A1(g1473), .A2(g1470), .A3(g1459) );
  NAND2_X1 NAND2_198( .ZN(g928), .A1(I1962), .A2(I1963) );
  NAND2_X1 NAND2_199( .ZN(I7097), .A1(g5194), .A2(g574) );
  NAND2_X1 NAND2_200( .ZN(I4547), .A1(g353), .A2(I4545) );
  NAND2_X1 NAND2_201( .ZN(I3697), .A1(g1570), .A2(g642) );
  NAND2_X1 NAND2_202( .ZN(I3914), .A1(g287), .A2(g2449) );
  NAND2_X1 NAND2_203( .ZN(I2543), .A1(g821), .A2(I2542) );
  NAND2_X1 NAND2_204( .ZN(I3413), .A1(g616), .A2(I3411) );
  NAND2_X1 NAND2_205( .ZN(I7218), .A1(g5368), .A2(I7216) );
  NAND2_X1 NAND2_206( .ZN(I7312), .A1(g5364), .A2(I7311) );
  NAND4_X1 NAND4_19( .ZN(g3538), .A1(g2588), .A2(g2215), .A3(g2197), .A4(g2179) );
  NAND2_X1 NAND2_207( .ZN(g5505), .A1(I7224), .A2(I7225) );
  NAND2_X1 NAND2_208( .ZN(g1075), .A1(I2109), .A2(I2110) );
  NAND2_X1 NAND2_209( .ZN(I2014), .A1(g532), .A2(I2013) );
  NAND2_X1 NAND2_210( .ZN(g2804), .A1(I4009), .A2(I4010) );
  NAND3_X1 NAND3_17( .ZN(g6742), .A1(g6683), .A2(g932), .A3(g6716) );
  NAND2_X1 NAND2_211( .ZN(I6185), .A1(g4301), .A2(g3955) );
  NAND4_X1 NAND4_20( .ZN(g5863), .A1(g5649), .A2(g1076), .A3(g1535), .A4(g2068) );
  NAND2_X1 NAND2_212( .ZN(I3739), .A1(g2021), .A2(g349) );
  NAND2_X1 NAND2_213( .ZN(I2022), .A1(g528), .A2(I2021) );
  NAND2_X2 NAND2_214( .ZN(I5782), .A1(g3810), .A2(g628) );
  NAND2_X2 NAND2_215( .ZN(I7576), .A1(g84), .A2(g5680) );
  NAND4_X1 NAND4_21( .ZN(g5688), .A1(g5546), .A2(g1585), .A3(g2084), .A4(g2916) );
  NAND4_X1 NAND4_22( .ZN(g5857), .A1(g5638), .A2(g1552), .A3(g1017), .A4(g2062) );
  NAND2_X2 NAND2_216( .ZN(I3190), .A1(g791), .A2(I3188) );
  NAND2_X2 NAND2_217( .ZN(I5292), .A1(g3421), .A2(g625) );
  NAND2_X2 NAND2_218( .ZN(g1764), .A1(I2796), .A2(I2797) );
  NAND2_X2 NAND2_219( .ZN(I3954), .A1(g2497), .A2(I3952) );
  NAND2_X2 NAND2_220( .ZN(g5779), .A1(I7549), .A2(I7550) );
  NAND2_X2 NAND2_221( .ZN(I7577), .A1(g84), .A2(I7576) );
  NAND2_X2 NAND2_222( .ZN(I5647), .A1(g3974), .A2(g3968) );
  NAND4_X1 NAND4_23( .ZN(g3531), .A1(g3209), .A2(g2215), .A3(g2976), .A4(g2179) );
  NAND2_X2 NAND2_223( .ZN(I1980), .A1(g230), .A2(I1978) );
  NAND2_X2 NAND2_224( .ZN(g5508), .A1(I7245), .A2(I7246) );
  NAND2_X1 NAND2_225( .ZN(I4150), .A1(g2551), .A2(g139) );
  NAND2_X1 NAND2_226( .ZN(g6873), .A1(g6848), .A2(g3621) );
  NAND2_X1 NAND2_227( .ZN(g6095), .A1(g2952), .A2(g5854) );
  NAND2_X1 NAND2_228( .ZN(I4009), .A1(g292), .A2(I4008) );
  NAND2_X1 NAND2_229( .ZN(I2675), .A1(g710), .A2(I2674) );
  NAND2_X1 NAND2_230( .ZN(g926), .A1(I1952), .A2(I1953) );
  NAND2_X1 NAND2_231( .ZN(I3894), .A1(g286), .A2(I3893) );
  NAND2_X1 NAND2_232( .ZN(I4212), .A1(g804), .A2(I4210) );
  NAND2_X1 NAND2_233( .ZN(g5565), .A1(I7312), .A2(I7313) );
  NAND2_X1 NAND2_234( .ZN(I6028), .A1(g4221), .A2(I6026) );
  NAND2_X1 NAND2_235( .ZN(I2109), .A1(g602), .A2(I2108) );
  NAND2_X1 NAND2_236( .ZN(I5244), .A1(g3247), .A2(I5242) );
  NAND3_X1 NAND3_18( .ZN(g1402), .A1(g310), .A2(g866), .A3(g873) );
  NAND2_X1 NAND2_237( .ZN(I4921), .A1(g650), .A2(I4919) );
  NAND2_X1 NAND2_238( .ZN(I7536), .A1(g5666), .A2(I7534) );
  NAND2_X1 NAND2_239( .ZN(I7223), .A1(g161), .A2(g5370) );
  NAND2_X2 NAND2_240( .ZN(I2498), .A1(g1042), .A2(I2497) );
  NAND2_X2 NAND2_241( .ZN(I1951), .A1(g524), .A2(g248) );
  NAND2_X2 NAND2_242( .ZN(I7522), .A1(g5659), .A2(I7520) );
  NAND2_X2 NAND2_243( .ZN(I3952), .A1(g289), .A2(g2497) );
  NAND2_X1 NAND2_244( .ZN(g5775), .A1(I7521), .A2(I7522) );
  NAND2_X1 NAND2_245( .ZN(I8201), .A1(g478), .A2(g6192) );
  NAND2_X1 NAND2_246( .ZN(g2024), .A1(I3126), .A2(I3127) );
  NAND2_X1 NAND2_247( .ZN(g2795), .A1(g1997), .A2(g866) );
  NAND2_X1 NAND2_248( .ZN(g4004), .A1(I5301), .A2(I5302) );
  NAND2_X1 NAND2_249( .ZN(I6196), .A1(g631), .A2(I6194) );
  NAND2_X1 NAND2_250( .ZN(I3970), .A1(g290), .A2(g2518) );
  NAND2_X1 NAND2_251( .ZN(I4941), .A1(g357), .A2(I4939) );
  NAND2_X1 NAND2_252( .ZN(I5657), .A1(g3983), .A2(g3979) );
  NAND2_X1 NAND2_253( .ZN(I7542), .A1(g59), .A2(I7541) );
  NAND2_X1 NAND2_254( .ZN(I2897), .A1(g1027), .A2(g634) );
  NAND2_X1 NAND2_255( .ZN(I2682), .A1(g918), .A2(I2681) );
  NAND2_X1 NAND2_256( .ZN(I2766), .A1(g749), .A2(g743) );
  NAND2_X1 NAND2_257( .ZN(g3013), .A1(I4211), .A2(I4212) );
  NAND2_X1 NAND2_258( .ZN(I5242), .A1(g3242), .A2(g3247) );
  NAND2_X1 NAND2_259( .ZN(I7529), .A1(g5662), .A2(I7527) );
  NAND2_X1 NAND2_260( .ZN(g1822), .A1(g1070), .A2(g1084) );
  NAND2_X1 NAND2_261( .ZN(I3876), .A1(g2397), .A2(I3874) );
  NAND2_X1 NAND2_262( .ZN(I2091), .A1(g29), .A2(I2089) );
  NAND2_X1 NAND2_263( .ZN(I3915), .A1(g287), .A2(I3914) );
  NAND2_X1 NAND2_264( .ZN(I9051), .A1(g6832), .A2(I9050) );
  NAND2_X1 NAND2_265( .ZN(I2767), .A1(g749), .A2(I2766) );
  NAND2_X1 NAND2_266( .ZN(I1979), .A1(g512), .A2(I1978) );
  NAND2_X1 NAND2_267( .ZN(g3597), .A1(I4783), .A2(I4784) );
  NAND3_X1 NAND3_19( .ZN(g2831), .A1(g2007), .A2(g862), .A3(g1784) );
  NAND2_X1 NAND2_268( .ZN(g5683), .A1(I7433), .A2(I7434) );
  NAND2_X1 NAND2_269( .ZN(g5778), .A1(I7542), .A2(I7543) );
  NAND2_X2 NAND2_270( .ZN(I2015), .A1(g260), .A2(I2013) );
  NAND2_X2 NAND2_271( .ZN(g930), .A1(I1970), .A2(I1971) );
  NAND2_X1 NAND2_272( .ZN(g5782), .A1(I7570), .A2(I7571) );
  NAND2_X1 NAND2_273( .ZN(g4002), .A1(I5293), .A2(I5294) );
  NAND2_X1 NAND2_274( .ZN(I2246), .A1(g598), .A2(I2244) );
  NAND2_X1 NAND2_275( .ZN(I6743), .A1(g4708), .A2(g582) );
  NAND2_X1 NAND2_276( .ZN(I7549), .A1(g64), .A2(I7548) );
  NAND2_X1 NAND2_277( .ZN(g2947), .A1(g1411), .A2(g2026) );
  NAND2_X1 NAND2_278( .ZN(g4762), .A1(I6391), .A2(I6392) );
  NAND3_X1 NAND3_20( .ZN(g2095), .A1(g1584), .A2(g749), .A3(g736) );
  NAND2_X1 NAND2_279( .ZN(g944), .A1(I2004), .A2(I2005) );
  NAND2_X1 NAND2_280( .ZN(I6474), .A1(g4541), .A2(I6473) );
  NAND2_X1 NAND2_281( .ZN(I7232), .A1(g5372), .A2(I7230) );
  NAND2_X1 NAND2_282( .ZN(I1953), .A1(g248), .A2(I1951) );
  NAND2_X1 NAND2_283( .ZN(g2719), .A1(I3875), .A2(I3876) );
  NAND2_X1 NAND2_284( .ZN(I8203), .A1(g6192), .A2(I8201) );
  NAND2_X1 NAND2_285( .ZN(I4008), .A1(g292), .A2(g2568) );
  NAND2_X1 NAND2_286( .ZN(g4237), .A1(g4049), .A2(g4017) );
  NAND2_X1 NAND2_287( .ZN(g1829), .A1(I2898), .A2(I2899) );
  NAND2_X1 NAND2_288( .ZN(g901), .A1(g314), .A2(g310) );
  NAND2_X1 NAND2_289( .ZN(g941), .A1(I1995), .A2(I1996) );
  NAND2_X1 NAND2_290( .ZN(I7570), .A1(g79), .A2(I7569) );
  NAND2_X1 NAND2_291( .ZN(I2108), .A1(g602), .A2(g610) );
  NAND2_X1 NAND2_292( .ZN(g1540), .A1(I2507), .A2(I2508) );
  NAND4_X1 NAND4_24( .ZN(g4814), .A1(g4550), .A2(g1575), .A3(g1550), .A4(g2073) );
  NAND2_X1 NAND2_293( .ZN(I7311), .A1(g5364), .A2(g590) );
  NAND2_X1 NAND2_294( .ZN(I5270), .A1(g3705), .A2(I5269) );
  NAND2_X1 NAND2_295( .ZN(g2745), .A1(I3915), .A2(I3916) );
  NAND3_X1 NAND3_21( .ZN(g1797), .A1(g98), .A2(g1064), .A3(g1070) );
  NAND2_X1 NAND2_296( .ZN(g2791), .A1(I3989), .A2(I3990) );
  NAND2_X1 NAND2_297( .ZN(I7239), .A1(g5374), .A2(I7237) );
  NAND4_X1 NAND4_25( .ZN(g3526), .A1(g3196), .A2(g3023), .A3(g2197), .A4(g2981) );
  NAND3_X1 NAND3_22( .ZN(g6741), .A1(g6705), .A2(g6461), .A3(g4941) );
  NAND2_X1 NAND2_298( .ZN(I8196), .A1(g6188), .A2(I8194) );
  NAND2_X1 NAND2_299( .ZN(I3895), .A1(g2422), .A2(I3893) );
  NAND2_X2 NAND2_300( .ZN(I4783), .A1(g2846), .A2(I4782) );
  NAND2_X1 NAND2_301( .ZN(I2021), .A1(g528), .A2(g254) );
  NAND2_X1 NAND2_302( .ZN(g905), .A1(g301), .A2(g319) );
  NAND2_X1 NAND2_303( .ZN(g3276), .A1(I4546), .A2(I4547) );
  NAND2_X1 NAND2_304( .ZN(g6774), .A1(g6754), .A2(g6750) );
  NAND2_X1 NAND2_305( .ZN(I5207), .A1(g3267), .A2(g3271) );
  NAND2_X1 NAND2_306( .ZN(I2301), .A1(g341), .A2(I2299) );
  NAND2_X1 NAND2_307( .ZN(I5259), .A1(g3719), .A2(I5257) );
  NAND2_X1 NAND2_308( .ZN(I7440), .A1(g5515), .A2(I7439) );
  NAND2_X1 NAND2_309( .ZN(I7528), .A1(g49), .A2(I7527) );
  NAND2_X1 NAND2_310( .ZN(g4640), .A1(g4402), .A2(g1056) );
  NAND4_X1 NAND4_26( .ZN(g4812), .A1(g4550), .A2(g1560), .A3(g1559), .A4(g2073) );
  NAND2_X2 NAND2_311( .ZN(g1845), .A1(I2934), .A2(I2935) );
  NAND2_X2 NAND2_312( .ZN(g6397), .A1(I8202), .A2(I8203) );
  NAND2_X1 NAND2_313( .ZN(I5768), .A1(g3957), .A2(I5766) );
  NAND2_X1 NAND2_314( .ZN(I1978), .A1(g512), .A2(g230) );
  NAND2_X1 NAND2_315( .ZN(g4610), .A1(I6186), .A2(I6187) );
  NAND2_X1 NAND2_316( .ZN(I5228), .A1(g3263), .A2(I5226) );
  NAND2_X1 NAND2_317( .ZN(I2074), .A1(g11), .A2(I2072) );
  NAND3_X1 NAND3_23( .ZN(g3140), .A1(g2409), .A2(g1060), .A3(g1620) );
  NAND2_X1 NAND2_318( .ZN(I6390), .A1(g4504), .A2(g4610) );
  NAND2_X1 NAND2_319( .ZN(I3177), .A1(g1706), .A2(g736) );
  NAND2_X1 NAND2_320( .ZN(I4152), .A1(g139), .A2(I4150) );
  NAND2_X1 NAND2_321( .ZN(I6501), .A1(g3541), .A2(I6499) );
  NAND2_X1 NAND2_322( .ZN(I7548), .A1(g64), .A2(g5672) );
  NAND2_X1 NAND2_323( .ZN(g1815), .A1(g102), .A2(g1070) );
  NAND2_X1 NAND2_324( .ZN(I7555), .A1(g69), .A2(g5674) );
  NAND4_X1 NAND4_27( .ZN(g3517), .A1(g3173), .A2(g3002), .A3(g2976), .A4(g2179) );
  NAND2_X1 NAND2_325( .ZN(I2080), .A1(g25), .A2(g19) );
  NAND2_X1 NAND2_326( .ZN(I4211), .A1(g2294), .A2(I4210) );
  NAND2_X1 NAND2_327( .ZN(I3399), .A1(g1826), .A2(I3398) );
  NAND2_X1 NAND2_328( .ZN(I5195), .A1(g3567), .A2(g3571) );
  NAND2_X1 NAND2_329( .ZN(I7313), .A1(g590), .A2(I7311) );
  NAND2_X1 NAND2_330( .ZN(g2582), .A1(I3698), .A2(I3699) );
  NAND2_X1 NAND2_331( .ZN(I4939), .A1(g3437), .A2(g357) );
  NAND2_X1 NAND2_332( .ZN(g950), .A1(I2022), .A2(I2023) );
  NAND2_X1 NAND2_333( .ZN(g4819), .A1(I6500), .A2(I6501) );
  NAND2_X1 NAND2_334( .ZN(I7521), .A1(g361), .A2(I7520) );
  NAND2_X1 NAND2_335( .ZN(I2023), .A1(g254), .A2(I2021) );
  NAND2_X1 NAND2_336( .ZN(I4446), .A1(g606), .A2(I4444) );
  NAND2_X1 NAND2_337( .ZN(I5783), .A1(g3810), .A2(I5782) );
  NAND2_X1 NAND2_338( .ZN(g2940), .A1(g197), .A2(g2381) );
  NAND2_X1 NAND2_339( .ZN(g4825), .A1(g4472), .A2(g4465) );
  NAND2_X1 NAND2_340( .ZN(I5293), .A1(g3421), .A2(I5292) );
  NAND2_X1 NAND2_341( .ZN(I5761), .A1(g3503), .A2(I5759) );
  NAND2_X1 NAND2_342( .ZN(I1971), .A1(g236), .A2(I1969) );
  NAND2_X1 NAND2_343( .ZN(I3972), .A1(g2518), .A2(I3970) );
  NAND2_X1 NAND2_344( .ZN(I4159), .A1(g2015), .A2(g619) );
  NAND2_X1 NAND2_345( .ZN(I6661), .A1(g3541), .A2(I6659) );
  NAND2_X1 NAND2_346( .ZN(g1398), .A1(g306), .A2(g889) );
  NAND2_X1 NAND2_347( .ZN(I6475), .A1(g578), .A2(I6473) );
  NAND2_X1 NAND2_348( .ZN(I3934), .A1(g288), .A2(I3933) );
  NAND2_X1 NAND2_349( .ZN(I7541), .A1(g59), .A2(g5669) );
  NAND2_X1 NAND2_350( .ZN(I2508), .A1(g1044), .A2(I2506) );
  NAND4_X1 NAND4_28( .ZN(g5854), .A1(g5638), .A2(g1683), .A3(g1552), .A4(g2062) );
  NAND2_X1 NAND2_351( .ZN(g4465), .A1(g319), .A2(g4253) );
  NAND2_X1 NAND2_352( .ZN(I2072), .A1(g15), .A2(g11) );
  NAND2_X2 NAND2_353( .ZN(I7238), .A1(g179), .A2(I7237) );
  NAND2_X2 NAND2_354( .ZN(g3955), .A1(I5188), .A2(I5189) );
  NAND2_X2 NAND2_355( .ZN(I7209), .A1(g143), .A2(I7208) );
  NAND2_X2 NAND2_356( .ZN(g5431), .A1(I7098), .A2(I7099) );
  NAND2_X1 NAND2_357( .ZN(I2681), .A1(g918), .A2(g613) );
  NAND2_X1 NAND2_358( .ZN(I2013), .A1(g532), .A2(g260) );
  NAND2_X1 NAND2_359( .ZN(I4234), .A1(g2267), .A2(I4233) );
  NAND2_X1 NAND2_360( .ZN(g2780), .A1(I3971), .A2(I3972) );
  NAND2_X1 NAND2_361( .ZN(g2067), .A1(I3178), .A2(I3179) );
  NAND2_X1 NAND2_362( .ZN(I1962), .A1(g520), .A2(I1961) );
  NAND2_X1 NAND2_363( .ZN(I5258), .A1(g3714), .A2(I5257) );
  NAND3_X1 NAND3_24( .ZN(g1387), .A1(g862), .A2(g314), .A3(g301) );
  NAND2_X1 NAND2_364( .ZN(I2060), .A1(g7), .A2(g3) );
  NAND2_X1 NAND2_365( .ZN(g5781), .A1(I7563), .A2(I7564) );
  NAND2_X1 NAND2_366( .ZN(g2263), .A1(I3399), .A2(I3400) );
  NAND2_X1 NAND2_367( .ZN(g4221), .A1(I5648), .A2(I5649) );
  NAND2_X1 NAND2_368( .ZN(g1359), .A1(g866), .A2(g306) );
  NAND2_X1 NAND2_369( .ZN(I7231), .A1(g170), .A2(I7230) );
  NAND2_X1 NAND2_370( .ZN(I3953), .A1(g289), .A2(I3952) );
  NAND2_X1 NAND2_371( .ZN(I5187), .A1(g3589), .A2(g3593) );
  NAND3_X1 NAND3_25( .ZN(g5852), .A1(g5638), .A2(g2053), .A3(g1661) );
  NAND4_X1 NAND4_29( .ZN(g3520), .A1(g3183), .A2(g3002), .A3(g2197), .A4(g2968) );
  NAND2_X2 NAND2_372( .ZN(g1047), .A1(I2090), .A2(I2091) );
  NAND2_X2 NAND2_373( .ZN(I7099), .A1(g574), .A2(I7097) );
  NAND2_X2 NAND2_374( .ZN(I3848), .A1(g2370), .A2(I3846) );
  NAND2_X1 NAND2_375( .ZN(I3699), .A1(g642), .A2(I3697) );
  NAND2_X1 NAND2_376( .ZN(I3398), .A1(g1826), .A2(g135) );
  NAND2_X1 NAND2_377( .ZN(I1969), .A1(g516), .A2(g236) );
  NAND2_X1 NAND2_378( .ZN(I5307), .A1(g478), .A2(g3512) );
  NAND2_X1 NAND2_379( .ZN(g3974), .A1(I5243), .A2(I5244) );
  NAND2_X1 NAND2_380( .ZN(I5536), .A1(g3907), .A2(I5535) );
  NAND2_X1 NAND2_381( .ZN(g1417), .A1(g873), .A2(g889) );
  NAND2_X1 NAND2_382( .ZN(I7543), .A1(g5669), .A2(I7541) );
  NAND2_X1 NAND2_383( .ZN(g5943), .A1(g5818), .A2(g2940) );
  NAND2_X1 NAND2_384( .ZN(I7534), .A1(g54), .A2(g5666) );
  NAND2_X1 NAND2_385( .ZN(g4319), .A1(I5783), .A2(I5784) );
  NAND2_X1 NAND2_386( .ZN(I3893), .A1(g286), .A2(g2422) );
  NAND2_X1 NAND2_387( .ZN(g2080), .A1(I3189), .A2(I3190) );
  NAND2_X1 NAND2_388( .ZN(I2683), .A1(g613), .A2(I2681) );
  NAND2_X1 NAND2_389( .ZN(I5537), .A1(g654), .A2(I5535) );
  NAND2_X1 NAND2_390( .ZN(I3170), .A1(g1534), .A2(I3168) );
  NAND2_X1 NAND2_391( .ZN(I3125), .A1(g1279), .A2(g1276) );
  NAND2_X1 NAND2_392( .ZN(I5243), .A1(g3242), .A2(I5242) );
  NAND2_X1 NAND2_393( .ZN(I1988), .A1(g224), .A2(I1986) );
  NAND2_X1 NAND2_394( .ZN(I6194), .A1(g4199), .A2(g631) );
  NAND2_X2 NAND2_395( .ZN(g3207), .A1(I4445), .A2(I4446) );
  NAND2_X2 NAND2_396( .ZN(I2526), .A1(g766), .A2(g719) );
  NAND2_X2 NAND2_397( .ZN(g6929), .A1(g4536), .A2(g6927) );
  NAND2_X1 NAND2_398( .ZN(g3215), .A1(g2340), .A2(g1402) );
  NAND2_X1 NAND2_399( .ZN(I3446), .A1(g1689), .A2(I3445) );
  NAND2_X1 NAND2_400( .ZN(I7208), .A1(g143), .A2(g5367) );
  NAND2_X1 NAND2_401( .ZN(g5783), .A1(I7577), .A2(I7578) );
  NAND2_X1 NAND2_402( .ZN(I4545), .A1(g2853), .A2(g353) );
  NAND2_X2 NAND2_403( .ZN(I2004), .A1(g500), .A2(I2003) );
  NAND2_X2 NAND2_404( .ZN(I2527), .A1(g766), .A2(I2526) );
  NAND2_X1 NAND2_405( .ZN(I5649), .A1(g3968), .A2(I5647) );
  NAND2_X1 NAND2_406( .ZN(g6778), .A1(g6762), .A2(g6758) );
  NAND2_X1 NAND2_407( .ZN(g1686), .A1(I2675), .A2(I2676) );
  NAND2_X1 NAND2_408( .ZN(g4223), .A1(I5658), .A2(I5659) );
  NAND2_X1 NAND2_409( .ZN(I1996), .A1(g218), .A2(I1994) );
  NAND2_X1 NAND2_410( .ZN(I3447), .A1(g729), .A2(I3445) );
  NAND2_X1 NAND2_411( .ZN(I4204), .A1(g2255), .A2(I4203) );
  NAND2_X1 NAND2_412( .ZN(I3874), .A1(g285), .A2(g2397) );
  NAND2_X1 NAND2_413( .ZN(g2944), .A1(g269), .A2(g2381) );
  NAND2_X1 NAND2_414( .ZN(g1253), .A1(I2245), .A2(I2246) );
  NAND3_X1 NAND3_26( .ZN(g2434), .A1(g1064), .A2(g1070), .A3(g1620) );
  NAND2_X1 NAND2_415( .ZN(I2299), .A1(g830), .A2(g341) );
  NAND3_X1 NAND3_27( .ZN(g5866), .A1(g5649), .A2(g1529), .A3(g2081) );
  NAND2_X1 NAND2_416( .ZN(g1687), .A1(I2682), .A2(I2683) );
  NAND2_X1 NAND2_417( .ZN(I3935), .A1(g2473), .A2(I3933) );
  NAND2_X1 NAND2_418( .ZN(g4017), .A1(g107), .A2(g3425) );
  NAND2_X1 NAND2_419( .ZN(I4528), .A1(g646), .A2(I4526) );
  NAND2_X1 NAND2_420( .ZN(I2244), .A1(g567), .A2(g598) );
  NAND2_X1 NAND2_421( .ZN(I4151), .A1(g2551), .A2(I4150) );
  NAND2_X1 NAND2_422( .ZN(I6392), .A1(g4610), .A2(I6390) );
  NAND2_X1 NAND2_423( .ZN(I4010), .A1(g2568), .A2(I4008) );
  NAND2_X1 NAND2_424( .ZN(I2082), .A1(g19), .A2(I2080) );
  NAND4_X1 NAND4_30( .ZN(g5818), .A1(g5638), .A2(g2056), .A3(g1666), .A4(g1661) );
  NAND2_X1 NAND2_425( .ZN(g3979), .A1(I5258), .A2(I5259) );
  NAND2_X1 NAND2_426( .ZN(I6176), .A1(g4236), .A2(I6175) );
  NAND2_X1 NAND2_427( .ZN(I4235), .A1(g798), .A2(I4233) );
  NAND2_X1 NAND2_428( .ZN(I2110), .A1(g610), .A2(I2108) );
  NAND2_X1 NAND2_429( .ZN(I7098), .A1(g5194), .A2(I7097) );
  NAND2_X1 NAND2_430( .ZN(I3456), .A1(g1691), .A2(I3455) );
  NAND4_X1 NAND4_31( .ZN(g5821), .A1(g5638), .A2(g2056), .A3(g1076), .A4(g1666) );
  NAND2_X1 NAND2_431( .ZN(I3698), .A1(g1570), .A2(I3697) );
  NAND2_X1 NAND2_432( .ZN(g2995), .A1(I4183), .A2(I4184) );
  NAND2_X1 NAND2_433( .ZN(I6473), .A1(g4541), .A2(g578) );
  NAND2_X1 NAND2_434( .ZN(I5659), .A1(g3979), .A2(I5657) );
  NAND2_X1 NAND2_435( .ZN(g5636), .A1(g5564), .A2(g4769) );
  NAND2_X1 NAND2_436( .ZN(I6177), .A1(g571), .A2(I6175) );
  NAND2_X1 NAND2_437( .ZN(I2899), .A1(g634), .A2(I2897) );
  NAND2_X1 NAND2_438( .ZN(I3457), .A1(g784), .A2(I3455) );
  NAND2_X1 NAND2_439( .ZN(I3989), .A1(g291), .A2(I3988) );
  NAND2_X1 NAND2_440( .ZN(I3971), .A1(g290), .A2(I3970) );
  NAND2_X1 NAND2_441( .ZN(I4160), .A1(g2015), .A2(I4159) );
  NAND2_X1 NAND2_442( .ZN(I2089), .A1(g33), .A2(g29) );
  NAND2_X2 NAND2_443( .ZN(g4670), .A1(g4611), .A2(g3528) );
  NAND4_X1 NAND4_32( .ZN(g4813), .A1(g4550), .A2(g965), .A3(g1560), .A4(g2073) );
  NAND2_X2 NAND2_444( .ZN(I3740), .A1(g2021), .A2(I3739) );
  NAND2_X1 NAND2_445( .ZN(I8194), .A1(g471), .A2(g6188) );
  NAND2_X1 NAND2_446( .ZN(I5300), .A1(g471), .A2(g3505) );
  NAND3_X1 NAND3_28( .ZN(g3893), .A1(g3664), .A2(g3656), .A3(g3647) );
  NAND2_X1 NAND2_447( .ZN(g6928), .A1(g4532), .A2(g6926) );
  NAND2_X1 NAND2_448( .ZN(I7578), .A1(g5680), .A2(I7576) );
  NAND2_X1 NAND2_449( .ZN(I7535), .A1(g54), .A2(I7534) );
  NAND2_X1 NAND2_450( .ZN(I1961), .A1(g520), .A2(g242) );
  NAND4_X1 NAND4_33( .ZN(g3544), .A1(g2594), .A2(g2215), .A3(g2197), .A4(g2179) );
  NAND2_X1 NAND2_451( .ZN(g6394), .A1(I8195), .A2(I8196) );
  NAND2_X1 NAND2_452( .ZN(I5648), .A1(g3974), .A2(I5647) );
  NAND2_X1 NAND2_453( .ZN(I7246), .A1(g5377), .A2(I7244) );
  NAND2_X1 NAND2_454( .ZN(g3756), .A1(I4940), .A2(I4941) );
  NAND2_X1 NAND2_455( .ZN(I2062), .A1(g3), .A2(I2060) );
  NAND2_X1 NAND2_456( .ZN(I6195), .A1(g4199), .A2(I6194) );
  NAND2_X1 NAND2_457( .ZN(I7216), .A1(g152), .A2(g5368) );
  NAND4_X1 NAND4_34( .ZN(g3536), .A1(g3219), .A2(g2215), .A3(g3007), .A4(g2179) );
  NAND2_X1 NAND2_458( .ZN(I7564), .A1(g5676), .A2(I7562) );
  NAND2_X1 NAND2_459( .ZN(g4300), .A1(I5760), .A2(I5761) );
  NAND2_X1 NAND2_460( .ZN(I4184), .A1(g749), .A2(I4182) );
  NAND2_X1 NAND2_461( .ZN(I2005), .A1(g212), .A2(I2003) );
  NAND2_X1 NAND2_462( .ZN(g5318), .A1(g676), .A2(g5060) );
  NAND4_X1 NAND4_35( .ZN(g5872), .A1(g5649), .A2(g1557), .A3(g1564), .A4(g2113) );
  NOR2_X2 NOR2_0( .ZN(g5552), .A1(g5354), .A2(g5356) );
  NOR2_X2 NOR2_1( .ZN(g4235), .A1(g3780), .A2(g3362) );
  NOR2_X1 NOR2_2( .ZN(g6073), .A1(g197), .A2(g5862) );
  NOR2_X1 NOR2_3( .ZN(g4776), .A1(g4449), .A2(g4453) );
  NOR2_X1 NOR2_4( .ZN(g4777), .A1(g4457), .A2(g4459) );
  NOR2_X1 NOR2_5( .ZN(g4238), .A1(g3755), .A2(g3279) );
  NOR3_X1 NOR4_0_A( .ZN(extra0), .A1(g6385), .A2(g3733), .A3(g4092) );
  NOR2_X1 NOR4_0( .ZN(g6433), .A1(extra0), .A2(g4314) );
  NOR2_X1 NOR2_6( .ZN(g6496), .A1(g952), .A2(g6354) );
  NOR2_X1 NOR2_7( .ZN(g1422), .A1(g1039), .A2(g913) );
  NOR2_X1 NOR2_8( .ZN(g3931), .A1(g3353), .A2(g3361) );
  NOR2_X1 NOR2_9( .ZN(g1560), .A1(g996), .A2(g980) );
  NOR2_X1 NOR2_10( .ZN(g3905), .A1(g3512), .A2(g478) );
  NOR2_X1 NOR2_11( .ZN(g5094), .A1(g4685), .A2(g4686) );
  NOR2_X1 NOR2_12( .ZN(g3973), .A1(g3368), .A2(g3374) );
  NOR2_X1 NOR2_13( .ZN(g3528), .A1(g1802), .A2(g3167) );
  NOR2_X1 NOR2_14( .ZN(g5541), .A1(g5388), .A2(g1880) );
  NOR2_X1 NOR2_15( .ZN(g3621), .A1(g1407), .A2(g2842) );
  NOR2_X1 NOR2_16( .ZN(g1449), .A1(g489), .A2(g1048) );
  NOR2_X2 NOR2_17( .ZN(g3965), .A1(g3359), .A2(g3367) );
  NOR2_X2 NOR2_18( .ZN(g3933), .A1(g3327), .A2(g3336) );
  NOR3_X2 NOR4_1_A( .ZN(extra1), .A1(I7978), .A2(I7979), .A3(I7980) );
  NOR2_X2 NOR4_1( .ZN(g6280), .A1(extra1), .A2(I7981) );
  NOR2_X1 NOR2_19( .ZN(g2433), .A1(g1418), .A2(g1449) );
  NOR3_X1 NOR3_0( .ZN(g1470), .A1(g937), .A2(g930), .A3(g928) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(g6376), .A2(g4086), .A3(g4074) );
  NOR2_X1 NOR4_2( .ZN(g6427), .A1(extra2), .A2(g4068) );
  NOR3_X1 NOR4_3_A( .ZN(extra3), .A1(g6385), .A2(g4334), .A3(g4092) );
  NOR2_X1 NOR4_3( .ZN(g6446), .A1(extra3), .A2(g4314) );
  NOR3_X1 NOR4_4_A( .ZN(extra4), .A1(I8135), .A2(I8136), .A3(I8137) );
  NOR2_X1 NOR4_4( .ZN(g6359), .A1(extra4), .A2(I8138) );
  NOR3_X1 NOR3_1( .ZN(g1459), .A1(g926), .A2(g950), .A3(g948) );
  NOR2_X1 NOR2_20( .ZN(g4584), .A1(g4164), .A2(g4168) );
  NOR2_X1 NOR2_21( .ZN(g3926), .A1(g3338), .A2(g3350) );
  NOR3_X1 NOR4_5_A( .ZN(extra5), .A1(I7969), .A2(I7970), .A3(I7971) );
  NOR2_X1 NOR4_5( .ZN(g6279), .A1(extra5), .A2(I7972) );
  NOR2_X1 NOR2_22( .ZN(g5265), .A1(g4863), .A2(g4865) );
  NOR2_X1 NOR2_23( .ZN(g3927), .A1(g3382), .A2(g3383) );
  NOR2_X1 NOR2_24( .ZN(g3903), .A1(g3505), .A2(g471) );
  NOR2_X1 NOR2_25( .ZN(g1418), .A1(g486), .A2(g943) );
  NOR2_X1 NOR2_26( .ZN(g4578), .A1(g4234), .A2(g3928) );
  NOR2_X1 NOR2_27( .ZN(g4261), .A1(g3762), .A2(g3295) );
  NOR3_X1 NOR4_6_A( .ZN(extra6), .A1(I8126), .A2(I8127), .A3(I8128) );
  NOR2_X1 NOR4_6( .ZN(g6358), .A1(extra6), .A2(I8129) );
  NOR2_X1 NOR2_28( .ZN(g4589), .A1(g4180), .A2(g4183) );
  NOR2_X1 NOR2_29( .ZN(g1474), .A1(g760), .A2(g754) );
  NOR2_X1 NOR2_30( .ZN(g3956), .A1(g3337), .A2(g3349) );
  NOR2_X1 NOR2_31( .ZN(g4774), .A1(g4442), .A2(g4445) );
  NOR2_X1 NOR2_32( .ZN(g5091), .A1(g4698), .A2(g4701) );
  NOR2_X1 NOR2_33( .ZN(g4950), .A1(g1472), .A2(g4680) );
  NOR2_X1 NOR2_34( .ZN(g5227), .A1(g5019), .A2(g3559) );
  NOR2_X1 NOR2_35( .ZN(g4585), .A1(g4171), .A2(g4177) );
  NOR2_X1 NOR2_36( .ZN(g6494), .A1(g952), .A2(g6348) );
  NOR3_X1 NOR3_2( .ZN(g5048), .A1(g4819), .A2(g3491), .A3(g3559) );
  NOR3_X1 NOR3_3( .ZN(g3664), .A1(g2804), .A2(g2791), .A3(g2780) );
  NOR2_X1 NOR2_37( .ZN(g4000), .A1(g1250), .A2(g3425) );
  NOR2_X1 NOR2_38( .ZN(g5418), .A1(g5162), .A2(g5169) );
  NOR2_X1 NOR2_39( .ZN(g5093), .A1(g4683), .A2(g4684) );
  NOR2_X1 NOR2_40( .ZN(g4779), .A1(g4461), .A2(g4464) );
  NOR2_X1 NOR2_41( .ZN(g6492), .A1(g6348), .A2(g1734) );
  NOR3_X1 NOR3_4( .ZN(g4240), .A1(g1589), .A2(g1879), .A3(g3793) );
  NOR2_X1 NOR2_42( .ZN(g4596), .A1(g4184), .A2(g4186) );
  NOR2_X1 NOR2_43( .ZN(g1603), .A1(g1039), .A2(g658) );
  NOR3_X1 NOR3_5( .ZN(g2908), .A1(g536), .A2(g2010), .A3(g541) );
  NOR2_X1 NOR2_44( .ZN(g4581), .A1(g4156), .A2(g4160) );
  NOR2_X1 NOR2_45( .ZN(g5423), .A1(g5170), .A2(g5175) );
  NOR2_X1 NOR2_46( .ZN(g4432), .A1(g923), .A2(g4253) );
  NOR3_X1 NOR4_7_A( .ZN(extra7), .A1(g6385), .A2(g3733), .A3(g4328) );
  NOR2_X1 NOR4_7( .ZN(g6436), .A1(extra7), .A2(g4080) );
  NOR2_X1 NOR2_47( .ZN(g4568), .A1(g4233), .A2(g3924) );
  NOR3_X1 NOR4_8_A( .ZN(extra8), .A1(I8079), .A2(I8080), .A3(I8081) );
  NOR2_X1 NOR4_8( .ZN(g6335), .A1(extra8), .A2(I8082) );
  NOR2_X1 NOR2_48( .ZN(g5753), .A1(g1477), .A2(g5688) );
  NOR2_X1 NOR2_49( .ZN(g6495), .A1(g6354), .A2(g1775) );
  NOR3_X1 NOR4_9_A( .ZN(extra9), .A1(g6376), .A2(g4323), .A3(g4074) );
  NOR2_X1 NOR4_9( .ZN(g6442), .A1(extra9), .A2(g4302) );
  NOR3_X1 NOR4_10_A( .ZN(extra10), .A1(g6376), .A2(g4086), .A3(g4074) );
  NOR2_X1 NOR4_10( .ZN(g6429), .A1(extra10), .A2(g4302) );
  NOR3_X1 NOR4_11_A( .ZN(extra11), .A1(I7987), .A2(I7988), .A3(I7989) );
  NOR2_X1 NOR4_11( .ZN(g6281), .A1(extra11), .A2(I7990) );
  NOR3_X1 NOR4_12_A( .ZN(extra12), .A1(g6385), .A2(g4334), .A3(g4328) );
  NOR2_X1 NOR4_12( .ZN(g6449), .A1(extra12), .A2(g4080) );
  NOR2_X1 NOR2_50( .ZN(g4590), .A1(g4169), .A2(g4172) );
  NOR2_X1 NOR2_51( .ZN(g4877), .A1(g952), .A2(g4680) );
  NOR3_X1 NOR4_13_A( .ZN(extra13), .A1(g6376), .A2(g4323), .A3(g4309) );
  NOR2_X1 NOR4_13( .ZN(g6445), .A1(extra13), .A2(g4068) );
  NOR3_X1 NOR4_14_A( .ZN(extra14), .A1(g5391), .A2(g1589), .A3(g3793) );
  NOR2_X1 NOR4_14( .ZN(g5561), .A1(extra14), .A2(g1880) );
  NOR2_X1 NOR2_52( .ZN(g3929), .A1(g3373), .A2(g3376) );
  NOR3_X1 NOR3_6( .ZN(g1473), .A1(g944), .A2(g941), .A3(g939) );
  NOR2_X1 NOR2_53( .ZN(g4967), .A1(g4674), .A2(g952) );
  NOR3_X1 NOR4_15_A( .ZN(extra15), .A1(g6385), .A2(g3733), .A3(g4092) );
  NOR2_X1 NOR4_15( .ZN(g6430), .A1(extra15), .A2(g4080) );
  NOR2_X1 NOR2_54( .ZN(g4993), .A1(g4674), .A2(g1477) );
  NOR3_X1 NOR4_16_A( .ZN(extra16), .A1(g6376), .A2(g4323), .A3(g4309) );
  NOR2_X1 NOR4_16( .ZN(g6448), .A1(extra16), .A2(g4302) );
  NOR3_X1 NOR3_7( .ZN(g3647), .A1(g2731), .A2(g2719), .A3(g2698) );
  NOR2_X1 NOR2_55( .ZN(g3925), .A1(g3303), .A2(g3315) );
  NOR2_X1 NOR2_56( .ZN(g5731), .A1(g952), .A2(g5688) );
  NOR2_X1 NOR2_57( .ZN(g3959), .A1(g3352), .A2(g3360) );
  NOR2_X1 NOR2_58( .ZN(g1481), .A1(g815), .A2(g809) );
  NOR3_X1 NOR3_8( .ZN(g3656), .A1(g2769), .A2(g2757), .A3(g2745) );
  NOR2_X1 NOR2_59( .ZN(g4245), .A1(g3759), .A2(g3288) );
  NOR2_X1 NOR2_60( .ZN(g3930), .A1(g3317), .A2(g3328) );
  NOR2_X1 NOR2_61( .ZN(g5249), .A1(g4868), .A2(g4870) );
  NOR2_X1 NOR2_62( .ZN(g3966), .A1(g3329), .A2(g3339) );
  NOR3_X1 NOR4_17_A( .ZN(extra17), .A1(I8208), .A2(I8209), .A3(I8210) );
  NOR2_X1 NOR4_17( .ZN(g6400), .A1(extra17), .A2(I8211) );
  NOR2_X1 NOR2_63( .ZN(g4266), .A1(g3757), .A2(g3283) );
  NOR3_X2 NOR4_18_A( .ZN(extra18), .A1(g6385), .A2(g4334), .A3(g4328) );
  NOR2_X2 NOR4_18( .ZN(g6451), .A1(extra18), .A2(g4314) );
  NOR3_X2 NOR3_9( .ZN(g5324), .A1(g5069), .A2(g4410), .A3(g766) );
  NOR3_X1 NOR4_19_A( .ZN(extra19), .A1(g6385), .A2(g4334), .A3(g4092) );
  NOR2_X1 NOR4_19( .ZN(g6443), .A1(extra19), .A2(g4080) );
  NOR2_X1 NOR2_64( .ZN(g5088), .A1(g4691), .A2(g4697) );
  NOR2_X1 NOR2_65( .ZN(g3958), .A1(g3316), .A2(g3326) );
  NOR2_X1 NOR2_66( .ZN(g4241), .A1(g3774), .A2(g3341) );
  NOR3_X1 NOR4_20_A( .ZN(extra20), .A1(g6376), .A2(g4086), .A3(g4309) );
  NOR2_X1 NOR4_20( .ZN(g6432), .A1(extra20), .A2(g4068) );
  NOR3_X1 NOR4_21_A( .ZN(extra21), .A1(I8117), .A2(I8118), .A3(I8119) );
  NOR2_X1 NOR4_21( .ZN(g6357), .A1(extra21), .A2(I8120) );
  NOR2_X1 NOR2_67( .ZN(g3923), .A1(g3378), .A2(g3381) );
  NOR2_X1 NOR2_68( .ZN(g6075), .A1(g269), .A2(g5863) );
  NOR2_X1 NOR2_69( .ZN(g3934), .A1(g3377), .A2(g3379) );
  NOR3_X1 NOR4_22_A( .ZN(extra22), .A1(g6385), .A2(g3733), .A3(g4328) );
  NOR2_X1 NOR4_22( .ZN(g6439), .A1(extra22), .A2(g4314) );
  NOR2_X1 NOR2_70( .ZN(g4272), .A1(g3767), .A2(g3319) );
  NOR2_X1 NOR2_71( .ZN(g1879), .A1(g1603), .A2(g1416) );
  NOR3_X1 NOR3_10( .ZN(g5325), .A1(g5077), .A2(g4416), .A3(g821) );
  NOR3_X1 NOR4_23_A( .ZN(extra23), .A1(g6376), .A2(g4086), .A3(g4309) );
  NOR2_X1 NOR4_23( .ZN(g6435), .A1(extra23), .A2(g4302) );
  NOR2_X1 NOR2_72( .ZN(g4586), .A1(g4161), .A2(g4165) );
  NOR2_X1 NOR2_73( .ZN(g3939), .A1(g3340), .A2(g3351) );
  NOR3_X1 NOR4_24_A( .ZN(extra24), .A1(g6376), .A2(g4323), .A3(g4074) );
  NOR2_X1 NOR4_24( .ZN(g6438), .A1(extra24), .A2(g4068) );
  NOR2_X1 NOR2_74( .ZN(g1518), .A1(g980), .A2(g965) );
  NOR2_X2 NOR2_75( .ZN(g4239), .A1(g3763), .A2(g3296) );
  NOR2_X1 NOR2_76( .ZN(g4591), .A1(g4178), .A2(g4181) );

endmodule
