//# 3 inputs
//# 6 outputs
//# 14 D-type flipflops
//# 44 inverters
//# 75 gates (31 ANDs + 9 NANDs + 16 ORs + 19 NORs)

module s298(CK,G0,G1,G117,G118,G132,G133,G2,G66,G67);
input CK,G0,G1,G2;
output G117,G132,G66,G118,G133,G67;

  wire G10,G29,G11,G30,G12,G34,G13,G39,G14,G44,G15,G56,G16,G86,G17,G92,
    G18,G98,G19,G102,G20,G107,G21,G113,G22,G119,G23,G125,G28,G130,G38,G40,
    G45,G46,G50,G51,G54,G55,G59,G60,G64,II155,II158,G76,G82,G87,G91,G93,
    G96,G99,G103,G108,G112,G114,II210,II213,G120,G124,G121,II221,G126,G131,G127,II229,
    II232,II235,II238,G26,G27,G31,G32,G33,G35,G36,G37,G42,G41,G48,G47,G49,
    G52,G57,G61,G58,G65,G62,G63,G74,G75,G88,G89,G90,G94,G95,G100,G105,
    G104,G110,G109,G111,G115,G122,G123,G128,G129,G24,G25,G68,G69,G70,G71,G72,
    G73,G77,G78,G79,G80,G81,G83,G84,G85,G43,G97,G101,G106,G116,G53,extra0,
    extra1,extra2;

  DFF_X1 DFF_0( .CK(CK), .Q(G10), .D(G29) );
  DFF_X1 DFF_1( .CK(CK), .Q(G11), .D(G30) );
  DFF_X2 DFF_2( .CK(CK), .Q(G12), .D(G34) );
  DFF_X2 DFF_3( .CK(CK), .Q(G13), .D(G39) );
  DFF_X1 DFF_4( .CK(CK), .Q(G14), .D(G44) );
  DFF_X1 DFF_5( .CK(CK), .Q(G15), .D(G56) );
  DFF_X1 DFF_6( .CK(CK), .Q(G16), .D(G86) );
  DFF_X1 DFF_7( .CK(CK), .Q(G17), .D(G92) );
  DFF_X1 DFF_8( .CK(CK), .Q(G18), .D(G98) );
  DFF_X1 DFF_9( .CK(CK), .Q(G19), .D(G102) );
  DFF_X1 DFF_10( .CK(CK), .Q(G20), .D(G107) );
  DFF_X1 DFF_11( .CK(CK), .Q(G21), .D(G113) );
  DFF_X2 DFF_12( .CK(CK), .Q(G22), .D(G119) );
  DFF_X1 DFF_13( .CK(CK), .Q(G23), .D(G125) );
  INV_X1 NOT_0( .ZN(G28), .A(G130) );
  INV_X1 NOT_1( .ZN(G38), .A(G10) );
  INV_X1 NOT_2( .ZN(G40), .A(G13) );
  INV_X1 NOT_3( .ZN(G45), .A(G12) );
  INV_X1 NOT_4( .ZN(G46), .A(G11) );
  INV_X1 NOT_5( .ZN(G50), .A(G14) );
  INV_X1 NOT_6( .ZN(G51), .A(G23) );
  INV_X1 NOT_7( .ZN(G54), .A(G11) );
  INV_X1 NOT_8( .ZN(G55), .A(G13) );
  INV_X1 NOT_9( .ZN(G59), .A(G12) );
  INV_X1 NOT_10( .ZN(G60), .A(G22) );
  INV_X1 NOT_11( .ZN(G64), .A(G15) );
  INV_X1 NOT_12( .ZN(II155), .A(G16) );
  INV_X1 NOT_13( .ZN(G66), .A(II155) );
  INV_X1 NOT_14( .ZN(II158), .A(G17) );
  INV_X1 NOT_15( .ZN(G67), .A(II158) );
  INV_X1 NOT_16( .ZN(G76), .A(G10) );
  INV_X1 NOT_17( .ZN(G82), .A(G11) );
  INV_X1 NOT_18( .ZN(G87), .A(G16) );
  INV_X1 NOT_19( .ZN(G91), .A(G12) );
  INV_X1 NOT_20( .ZN(G93), .A(G17) );
  INV_X1 NOT_21( .ZN(G96), .A(G14) );
  INV_X1 NOT_22( .ZN(G99), .A(G18) );
  INV_X1 NOT_23( .ZN(G103), .A(G13) );
  INV_X1 NOT_24( .ZN(G108), .A(G112) );
  INV_X1 NOT_25( .ZN(G114), .A(G21) );
  INV_X2 NOT_26( .ZN(II210), .A(G18) );
  INV_X2 NOT_27( .ZN(G117), .A(II210) );
  INV_X4 NOT_28( .ZN(II213), .A(G19) );
  INV_X8 NOT_29( .ZN(G118), .A(II213) );
  INV_X8 NOT_30( .ZN(G120), .A(G124) );
  INV_X16 NOT_31( .ZN(G121), .A(G22) );
  INV_X1 NOT_32( .ZN(II221), .A(G2) );
  INV_X1 NOT_33( .ZN(G124), .A(II221) );
  INV_X1 NOT_34( .ZN(G126), .A(G131) );
  INV_X1 NOT_35( .ZN(G127), .A(G23) );
  INV_X1 NOT_36( .ZN(II229), .A(G0) );
  INV_X1 NOT_37( .ZN(G130), .A(II229) );
  INV_X1 NOT_38( .ZN(II232), .A(G1) );
  INV_X1 NOT_39( .ZN(G131), .A(II232) );
  INV_X1 NOT_40( .ZN(II235), .A(G20) );
  INV_X2 NOT_41( .ZN(G132), .A(II235) );
  INV_X2 NOT_42( .ZN(II238), .A(G21) );
  INV_X2 NOT_43( .ZN(G133), .A(II238) );
  AND2_X1 AND2_0( .ZN(G26), .A1(G28), .A2(G50) );
  AND2_X1 AND2_1( .ZN(G27), .A1(G51), .A2(G28) );
  AND3_X1 AND3_0( .ZN(G31), .A1(G10), .A2(G45), .A3(G13) );
  AND2_X1 AND2_2( .ZN(G32), .A1(G10), .A2(G11) );
  AND2_X1 AND2_3( .ZN(G33), .A1(G38), .A2(G46) );
  AND3_X1 AND3_1( .ZN(G35), .A1(G10), .A2(G11), .A3(G12) );
  AND2_X1 AND2_4( .ZN(G36), .A1(G38), .A2(G45) );
  AND2_X1 AND2_5( .ZN(G37), .A1(G46), .A2(G45) );
  AND2_X1 AND2_6( .ZN(G42), .A1(G40), .A2(G41) );
  AND4_X1 AND4_0( .ZN(G48), .A1(G45), .A2(G46), .A3(G10), .A4(G47) );
  AND3_X1 AND3_2( .ZN(G49), .A1(G50), .A2(G51), .A3(G52) );
  AND4_X2 AND4_1( .ZN(G57), .A1(G59), .A2(G11), .A3(G60), .A4(G61) );
  AND2_X2 AND2_7( .ZN(G58), .A1(G64), .A2(G65) );
  AND4_X1 AND4_2( .ZN(G62), .A1(G59), .A2(G11), .A3(G60), .A4(G61) );
  AND2_X1 AND2_8( .ZN(G63), .A1(G64), .A2(G65) );
  AND3_X1 AND3_3( .ZN(G74), .A1(G12), .A2(G14), .A3(G19) );
  AND3_X1 AND3_4( .ZN(G75), .A1(G82), .A2(G91), .A3(G14) );
  AND2_X1 AND2_9( .ZN(G88), .A1(G14), .A2(G87) );
  AND2_X1 AND2_10( .ZN(G89), .A1(G103), .A2(G96) );
  AND2_X1 AND2_11( .ZN(G90), .A1(G91), .A2(G103) );
  AND2_X1 AND2_12( .ZN(G94), .A1(G93), .A2(G13) );
  AND2_X1 AND2_13( .ZN(G95), .A1(G96), .A2(G13) );
  AND3_X1 AND3_5( .ZN(G100), .A1(G99), .A2(G14), .A3(G12) );
  AND3_X2 AND3_6( .ZN(G105), .A1(G103), .A2(G108), .A3(G104) );
  AND2_X2 AND2_14( .ZN(G110), .A1(G108), .A2(G109) );
  AND2_X2 AND2_15( .ZN(G111), .A1(G10), .A2(G112) );
  AND2_X1 AND2_16( .ZN(G115), .A1(G114), .A2(G14) );
  AND2_X1 AND2_17( .ZN(G122), .A1(G120), .A2(G121) );
  AND2_X1 AND2_18( .ZN(G123), .A1(G124), .A2(G22) );
  AND2_X1 AND2_19( .ZN(G128), .A1(G126), .A2(G127) );
  AND2_X1 AND2_20( .ZN(G129), .A1(G131), .A2(G23) );
  OR4_X1 OR4_0( .ZN(G24), .A1(G38), .A2(G46), .A3(G45), .A4(G40) );
  OR3_X1 OR3_0( .ZN(G25), .A1(G38), .A2(G11), .A3(G12) );
  OR4_X1 OR4_1( .ZN(G68), .A1(G11), .A2(G12), .A3(G13), .A4(G96) );
  OR2_X1 OR2_0( .ZN(G69), .A1(G103), .A2(G18) );
  OR2_X1 OR2_1( .ZN(G70), .A1(G103), .A2(G14) );
  OR3_X2 OR3_1( .ZN(G71), .A1(G82), .A2(G12), .A3(G13) );
  OR2_X2 OR2_2( .ZN(G72), .A1(G91), .A2(G20) );
  OR2_X2 OR2_3( .ZN(G73), .A1(G103), .A2(G20) );
  OR4_X1 OR4_2( .ZN(G77), .A1(G112), .A2(G103), .A3(G96), .A4(G19) );
  OR2_X1 OR2_4( .ZN(G78), .A1(G108), .A2(G76) );
  OR2_X1 OR2_5( .ZN(G79), .A1(G103), .A2(G14) );
  OR2_X1 OR2_6( .ZN(G80), .A1(G11), .A2(G14) );
  OR2_X1 OR2_7( .ZN(G81), .A1(G12), .A2(G13) );
  OR4_X1 OR4_3( .ZN(G83), .A1(G11), .A2(G12), .A3(G13), .A4(G96) );
  OR3_X1 OR3_2( .ZN(G84), .A1(G82), .A2(G91), .A3(G14) );
  OR3_X1 OR3_3( .ZN(G85), .A1(G91), .A2(G96), .A3(G17) );
  NAND3_X1 NAND3_0( .ZN(G41), .A1(G12), .A2(G11), .A3(G10) );
  NAND3_X1 NAND3_1( .ZN(G43), .A1(G24), .A2(G25), .A3(G28) );
  NAND4_X1 NAND4_0( .ZN(G52), .A1(G13), .A2(G45), .A3(G46), .A4(G10) );
  NAND4_X2 NAND4_1( .ZN(G65), .A1(G59), .A2(G54), .A3(G22), .A4(G61) );
  NAND4_X1 NAND4_2( .ZN(G97), .A1(G83), .A2(G84), .A3(G85), .A4(G108) );
  NAND4_X1 NAND4_3( .ZN(G101), .A1(G68), .A2(G69), .A3(G70), .A4(G108) );
  NAND2_X1 NAND2_0( .ZN(G106), .A1(G77), .A2(G78) );
  NAND4_X2 NAND4_4( .ZN(G109), .A1(G71), .A2(G72), .A3(G73), .A4(G14) );
  NAND4_X1 NAND4_5( .ZN(G116), .A1(G79), .A2(G80), .A3(G81), .A4(G108) );
  NOR2_X1 NOR2_0( .ZN(G29), .A1(G10), .A2(G130) );
  NOR3_X1 NOR4_0_A( .ZN(extra0), .A1(G31), .A2(G32), .A3(G33) );
  NOR2_X1 NOR4_0( .ZN(G30), .A1(extra0), .A2(G130) );
  NOR3_X1 NOR4_1_A( .ZN(extra1), .A1(G35), .A2(G36), .A3(G37) );
  NOR2_X1 NOR4_1( .ZN(G34), .A1(extra1), .A2(G130) );
  NOR2_X2 NOR2_1( .ZN(G39), .A1(G42), .A2(G43) );
  NOR3_X1 NOR3_0( .ZN(G44), .A1(G48), .A2(G49), .A3(G53) );
  NOR2_X1 NOR2_2( .ZN(G47), .A1(G50), .A2(G40) );
  NOR2_X1 NOR2_3( .ZN(G53), .A1(G26), .A2(G27) );
  NOR3_X1 NOR3_1( .ZN(G56), .A1(G57), .A2(G58), .A3(G130) );
  NOR2_X1 NOR2_4( .ZN(G61), .A1(G14), .A2(G55) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(G88), .A2(G89), .A3(G90) );
  NOR2_X1 NOR4_2( .ZN(G86), .A1(extra2), .A2(G112) );
  NOR3_X1 NOR3_2( .ZN(G92), .A1(G94), .A2(G95), .A3(G97) );
  NOR2_X1 NOR2_5( .ZN(G98), .A1(G100), .A2(G101) );
  NOR2_X1 NOR2_6( .ZN(G102), .A1(G105), .A2(G106) );
  NOR2_X2 NOR2_7( .ZN(G104), .A1(G74), .A2(G75) );
  NOR2_X2 NOR2_8( .ZN(G107), .A1(G110), .A2(G111) );
  NOR2_X1 NOR2_9( .ZN(G112), .A1(G62), .A2(G63) );
  NOR2_X1 NOR2_10( .ZN(G113), .A1(G115), .A2(G116) );
  NOR3_X1 NOR3_3( .ZN(G119), .A1(G122), .A2(G123), .A3(G130) );
  NOR3_X2 NOR3_4( .ZN(G125), .A1(G128), .A2(G129), .A3(G130) );

endmodule
