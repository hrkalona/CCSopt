//# 3 inputs
//# 6 outputs
//# 21 D-type flipflops
//# 59 inverters
//# 99 gates (11 ANDs + 30 NANDs + 24 ORs + 34 NORs)

module s382(CK,CLR,FM,GRN1,GRN2,RED1,RED2,TEST,YLW1,YLW2);
input CK,FM,TEST,CLR;
output GRN1,GRN2,RED1,YLW2,RED2,YLW1;

  wire TESTL,TESTLVIINLATCHVCDAD,FML,FMLVIINLATCHVCDAD,OLATCH_Y2L,TCOMB_YA2,OLATCHVUC_6,Y1C,OLATCHVUC_5,R2C,OLATCH_R1L,TCOMB_RA1,OLATCH_G2L,TCOMB_GA2,OLATCH_G1L,TCOMB_GA1,
    OLATCH_FEL,TCOMB_FE_BF,C3_Q3,C3_Q3VD,C3_Q2,C3_Q2VD,C3_Q1,C3_Q1VD,C3_Q0,C3_Q0VD,UC_16,UC_16VD,UC_17,UC_17VD,UC_18,UC_18VD,
    UC_19,UC_19VD,UC_8,UC_8VD,UC_9,UC_9VD,UC_10,UC_10VD,UC_11,UC_11VD,TESTLVIINLATCHN,FMLVIINLATCHN,OLATCH_Y1L,OLATCH_R2L,UC_23,UC_24,
    UC_25,UC_26,UC_20,C2_QN2,UC_21,UC_22,UC_12,UC_13,UC_14,UC_15,FMBVIIR1,CLRBVIIR1,TCOMBVNFM,TESTBVIIR1,TCOMBVNQA,TCOMBVNQB,
    TCOMBVNQC,TCOMBVNQD,UC_11VUC_0,OUTBUFVBUFG1VIIR1,OUTBUFVBUFG2VIIR1,TCOMBVNFEL,OUTBUFVBUFR1VIIR1,OUTBUFVBUFY2VIIR1,FMB,CLRB,TESTB,UC_11VZ,C1VCO0,OUTBUFVBUFR2VIIR1,OUTBUFVBUFY1VIIR1,FMLVIINMUXVIIR1,
    TESTLVIINLATCHVCDN,FMLVIINLATCHVCDN,TCOMBVNCLR,TESTLVIINMUXVIIR1,C2VIINHN,CTST,UC_8VZ,UC_8VZVOR1NF,CO2,C2_CO,FMLVIINMUX,FMLVIINMUXVND1,TESTLVIINMUX,TESTLVIINMUXVND1,II84,TCOMB_FE,
    FEN,UC_16VZ,UC_16VZVOR1NF,C3VIINHN,C3_Q3VZ,C3_Q3VZVOR1NF,TCOMB_GA1VAD1NF,TCOMBVNODE6,TCOMB_GA2VAD4NF,TCOMB_GA2VAD3NF,TCOMB_GA2VAD2NF,TCOMB_GA2VAD1NF,R2CVAD1NF,Y1CVAD1NF,TCOMB_YA1,Y1CVAD2NF,
    R2CVAD2NF,TCOMB_RA2,TCOMB_RA1VOR2NF,TCOMBVNODE8VOR1NF,TCOMB_RA1VOR1NF,TCOMBVNODE8VOR2NF,FMLVIINMUXVOR1NF,TCOMB_RA2VOR3NF,TCOMB_RA2VOR1NF,TCOMBVNODE4VOR2NF,TCOMBVNODE4VOR1NF,TESTLVIINMUXVOR1NF,TCOMBVNODE16VOR1NF,TCOMBVNODE18,C1VCO2,UC_9VZVOR1NF,
    C1VCO1,UC_10VZVOR1NF,FMLVIINMUXVOR2NF,TESTLVIINMUXVOR2NF,C2VCO2,UC_17VZVOR1NF,C2VCO1,UC_18VZVOR1NF,C2VCO0,UC_19VZVOR1NF,C3VCO2,C3_Q2VZVOR1NF,C3VCO1,C3_Q1VZVOR1NF,C3VCO0,C3_Q0VZVOR1NF,
    UC_9VUC_0,UC_10VUC_0,TCOMBVNODE4,TCOMBVNODE14,TCOMBVNODE15,TCOMBVNODE12,TCOMBVNODE8,TCOMBVNODE16,TCOMBVNODE19,UC_9VZ,UC_10VZ,TCOMBVNODE3,UC_17VUC_0,UC_18VUC_0,UC_19VUC_0,UC_17VZ,
    UC_18VZ,UC_19VZ,C3_Q2VUC_0,C3_Q1VUC_0,C3_Q0VUC_0,C3_Q2VZ,C3_Q1VZ,C3_Q0VZ,C3VCIIA,C1VCIIA,C2VCIIA,C1_CO,UC_27,extra0,extra1,extra2,
    extra3;

  DFF_X1 DFF_0( .CK(CK), .Q(TESTL), .D(TESTLVIINLATCHVCDAD) );
  DFF_X1 DFF_1( .CK(CK), .Q(FML), .D(FMLVIINLATCHVCDAD) );
  DFF_X2 DFF_2( .CK(CK), .Q(OLATCH_Y2L), .D(TCOMB_YA2) );
  DFF_X2 DFF_3( .CK(CK), .Q(OLATCHVUC_6), .D(Y1C) );
  DFF_X2 DFF_4( .CK(CK), .Q(OLATCHVUC_5), .D(R2C) );
  DFF_X1 DFF_5( .CK(CK), .Q(OLATCH_R1L), .D(TCOMB_RA1) );
  DFF_X1 DFF_6( .CK(CK), .Q(OLATCH_G2L), .D(TCOMB_GA2) );
  DFF_X1 DFF_7( .CK(CK), .Q(OLATCH_G1L), .D(TCOMB_GA1) );
  DFF_X1 DFF_8( .CK(CK), .Q(OLATCH_FEL), .D(TCOMB_FE_BF) );
  DFF_X1 DFF_9( .CK(CK), .Q(C3_Q3), .D(C3_Q3VD) );
  DFF_X1 DFF_10( .CK(CK), .Q(C3_Q2), .D(C3_Q2VD) );
  DFF_X1 DFF_11( .CK(CK), .Q(C3_Q1), .D(C3_Q1VD) );
  DFF_X1 DFF_12( .CK(CK), .Q(C3_Q0), .D(C3_Q0VD) );
  DFF_X2 DFF_13( .CK(CK), .Q(UC_16), .D(UC_16VD) );
  DFF_X1 DFF_14( .CK(CK), .Q(UC_17), .D(UC_17VD) );
  DFF_X1 DFF_15( .CK(CK), .Q(UC_18), .D(UC_18VD) );
  DFF_X1 DFF_16( .CK(CK), .Q(UC_19), .D(UC_19VD) );
  DFF_X1 DFF_17( .CK(CK), .Q(UC_8), .D(UC_8VD) );
  DFF_X1 DFF_18( .CK(CK), .Q(UC_9), .D(UC_9VD) );
  DFF_X1 DFF_19( .CK(CK), .Q(UC_10), .D(UC_10VD) );
  DFF_X1 DFF_20( .CK(CK), .Q(UC_11), .D(UC_11VD) );
  INV_X1 NOT_0( .ZN(TESTLVIINLATCHN), .A(TESTL) );
  INV_X1 NOT_1( .ZN(FMLVIINLATCHN), .A(FML) );
  INV_X1 NOT_2( .ZN(OLATCH_Y1L), .A(OLATCHVUC_6) );
  INV_X1 NOT_3( .ZN(OLATCH_R2L), .A(OLATCHVUC_5) );
  INV_X1 NOT_4( .ZN(UC_23), .A(C3_Q3) );
  INV_X1 NOT_5( .ZN(UC_24), .A(C3_Q2) );
  INV_X1 NOT_6( .ZN(UC_25), .A(C3_Q1) );
  INV_X1 NOT_7( .ZN(UC_26), .A(C3_Q0) );
  INV_X1 NOT_8( .ZN(UC_20), .A(UC_16) );
  INV_X1 NOT_9( .ZN(C2_QN2), .A(UC_17) );
  INV_X1 NOT_10( .ZN(UC_21), .A(UC_18) );
  INV_X1 NOT_11( .ZN(UC_22), .A(UC_19) );
  INV_X1 NOT_12( .ZN(UC_12), .A(UC_8) );
  INV_X1 NOT_13( .ZN(UC_13), .A(UC_9) );
  INV_X1 NOT_14( .ZN(UC_14), .A(UC_10) );
  INV_X2 NOT_15( .ZN(UC_15), .A(UC_11) );
  INV_X2 NOT_16( .ZN(FMBVIIR1), .A(FM) );
  INV_X2 NOT_17( .ZN(CLRBVIIR1), .A(CLR) );
  INV_X2 NOT_18( .ZN(TCOMBVNFM), .A(FML) );
  INV_X2 NOT_19( .ZN(TESTBVIIR1), .A(TEST) );
  INV_X1 NOT_20( .ZN(TCOMBVNQA), .A(C3_Q0) );
  INV_X1 NOT_21( .ZN(TCOMBVNQB), .A(C3_Q1) );
  INV_X1 NOT_22( .ZN(TCOMBVNQC), .A(C3_Q2) );
  INV_X1 NOT_23( .ZN(TCOMBVNQD), .A(C3_Q3) );
  INV_X1 NOT_24( .ZN(UC_11VUC_0), .A(UC_11) );
  INV_X1 NOT_25( .ZN(OUTBUFVBUFG1VIIR1), .A(OLATCH_G1L) );
  INV_X1 NOT_26( .ZN(OUTBUFVBUFG2VIIR1), .A(OLATCH_G2L) );
  INV_X1 NOT_27( .ZN(TCOMBVNFEL), .A(OLATCH_FEL) );
  INV_X1 NOT_28( .ZN(OUTBUFVBUFR1VIIR1), .A(OLATCH_R1L) );
  INV_X1 NOT_29( .ZN(OUTBUFVBUFY2VIIR1), .A(OLATCH_Y2L) );
  INV_X1 NOT_30( .ZN(FMB), .A(FMBVIIR1) );
  INV_X1 NOT_31( .ZN(CLRB), .A(CLRBVIIR1) );
  INV_X1 NOT_32( .ZN(TESTB), .A(TESTBVIIR1) );
  INV_X1 NOT_33( .ZN(UC_11VZ), .A(UC_11VUC_0) );
  INV_X1 NOT_34( .ZN(C1VCO0), .A(UC_15) );
  INV_X1 NOT_35( .ZN(GRN1), .A(OUTBUFVBUFG1VIIR1) );
  INV_X1 NOT_36( .ZN(GRN2), .A(OUTBUFVBUFG2VIIR1) );
  INV_X1 NOT_37( .ZN(RED1), .A(OUTBUFVBUFR1VIIR1) );
  INV_X1 NOT_38( .ZN(YLW2), .A(OUTBUFVBUFY2VIIR1) );
  INV_X1 NOT_39( .ZN(OUTBUFVBUFR2VIIR1), .A(OLATCH_R2L) );
  INV_X1 NOT_40( .ZN(OUTBUFVBUFY1VIIR1), .A(OLATCH_Y1L) );
  INV_X1 NOT_41( .ZN(FMLVIINMUXVIIR1), .A(FMB) );
  INV_X1 NOT_42( .ZN(TESTLVIINLATCHVCDN), .A(CLRB) );
  INV_X1 NOT_43( .ZN(FMLVIINLATCHVCDN), .A(CLRB) );
  INV_X4 NOT_44( .ZN(TCOMBVNCLR), .A(CLRB) );
  INV_X4 NOT_45( .ZN(TESTLVIINMUXVIIR1), .A(TESTB) );
  INV_X4 NOT_46( .ZN(RED2), .A(OUTBUFVBUFR2VIIR1) );
  INV_X4 NOT_47( .ZN(YLW1), .A(OUTBUFVBUFY1VIIR1) );
  INV_X1 NOT_48( .ZN(C2VIINHN), .A(CTST) );
  INV_X1 NOT_49( .ZN(UC_8VZ), .A(UC_8VZVOR1NF) );
  INV_X1 NOT_50( .ZN(CO2), .A(C2_CO) );
  INV_X1 NOT_51( .ZN(FMLVIINMUX), .A(FMLVIINMUXVND1) );
  INV_X1 NOT_52( .ZN(TESTLVIINMUX), .A(TESTLVIINMUXVND1) );
  INV_X1 NOT_53( .ZN(II84), .A(TCOMB_FE) );
  INV_X1 NOT_54( .ZN(FEN), .A(TCOMB_FE) );
  INV_X1 NOT_55( .ZN(UC_16VZ), .A(UC_16VZVOR1NF) );
  INV_X1 NOT_56( .ZN(C3VIINHN), .A(CO2) );
  INV_X1 NOT_57( .ZN(TCOMB_FE_BF), .A(II84) );
  INV_X1 NOT_58( .ZN(C3_Q3VZ), .A(C3_Q3VZVOR1NF) );
  AND2_X1 AND2_0( .ZN(TCOMB_GA1VAD1NF), .A1(TCOMBVNODE6), .A2(OLATCH_FEL) );
  AND2_X1 AND2_1( .ZN(TCOMB_GA2VAD4NF), .A1(OLATCH_FEL), .A2(TCOMBVNCLR) );
  AND2_X1 AND2_2( .ZN(TCOMB_GA2VAD3NF), .A1(C3_Q2), .A2(TCOMBVNCLR) );
  AND3_X1 AND3_0( .ZN(TCOMB_GA2VAD2NF), .A1(C3_Q0), .A2(C3_Q1), .A3(TCOMBVNCLR) );
  AND3_X1 AND3_1( .ZN(TCOMB_GA2VAD1NF), .A1(TCOMBVNQA), .A2(C3_Q3), .A3(TCOMBVNCLR) );
  AND2_X1 AND2_3( .ZN(R2CVAD1NF), .A1(TCOMB_FE), .A2(C2_QN2) );
  AND2_X4 AND2_4( .ZN(FMLVIINLATCHVCDAD), .A1(FMLVIINLATCHVCDN), .A2(FMLVIINMUX) );
  AND2_X4 AND2_5( .ZN(Y1CVAD1NF), .A1(TCOMB_YA1), .A2(C2_QN2) );
  AND2_X2 AND2_6( .ZN(TESTLVIINLATCHVCDAD), .A1(TESTLVIINLATCHVCDN), .A2(TESTLVIINMUX) );
  AND2_X1 AND2_7( .ZN(Y1CVAD2NF), .A1(FEN), .A2(TCOMB_YA1) );
  AND2_X1 AND2_8( .ZN(R2CVAD2NF), .A1(FEN), .A2(TCOMB_RA2) );
  OR3_X1 OR3_0( .ZN(TCOMB_RA1VOR2NF), .A1(C3_Q2), .A2(C3_Q3), .A3(OLATCH_FEL) );
  OR3_X1 OR3_1( .ZN(TCOMBVNODE8VOR1NF), .A1(C3_Q0), .A2(C3_Q1), .A3(TCOMBVNFM) );
  OR4_X1 OR4_0( .ZN(TCOMB_RA1VOR1NF), .A1(TCOMBVNQA), .A2(C3_Q1), .A3(C3_Q2), .A4(OLATCH_FEL) );
  OR2_X1 OR2_0( .ZN(TCOMBVNODE8VOR2NF), .A1(TCOMBVNQD), .A2(TCOMBVNFM) );
  OR2_X1 OR2_1( .ZN(FMLVIINMUXVOR1NF), .A1(FMB), .A2(FML) );
  OR2_X1 OR2_2( .ZN(TCOMB_RA2VOR3NF), .A1(TCOMBVNQC), .A2(CLRB) );
  OR4_X1 OR4_1( .ZN(TCOMB_RA2VOR1NF), .A1(C3_Q0), .A2(C3_Q1), .A3(TCOMBVNQD), .A4(CLRB) );
  OR3_X1 OR3_2( .ZN(TCOMBVNODE4VOR2NF), .A1(C3_Q2), .A2(TCOMBVNQD), .A3(CLRB) );
  OR4_X1 OR4_2( .ZN(TCOMBVNODE4VOR1NF), .A1(TCOMBVNQC), .A2(C3_Q3), .A3(TCOMBVNFM), .A4(CLRB) );
  OR2_X1 OR2_3( .ZN(TESTLVIINMUXVOR1NF), .A1(TESTB), .A2(TESTL) );
  OR4_X1 OR4_3( .ZN(TCOMBVNODE16VOR1NF), .A1(TCOMBVNODE18), .A2(FML), .A3(C3_Q3), .A4(TCOMBVNQC) );
  OR2_X1 OR2_4( .ZN(UC_8VZVOR1NF), .A1(C1VCO2), .A2(UC_8) );
  OR2_X1 OR2_5( .ZN(UC_9VZVOR1NF), .A1(C1VCO1), .A2(UC_9) );
  OR2_X1 OR2_6( .ZN(UC_10VZVOR1NF), .A1(C1VCO0), .A2(UC_10) );
  OR2_X2 OR2_7( .ZN(FMLVIINMUXVOR2NF), .A1(FMLVIINMUXVIIR1), .A2(FMLVIINLATCHN) );
  OR2_X2 OR2_8( .ZN(TESTLVIINMUXVOR2NF), .A1(TESTLVIINMUXVIIR1), .A2(TESTLVIINLATCHN) );
  OR2_X2 OR2_9( .ZN(UC_16VZVOR1NF), .A1(C2VCO2), .A2(UC_16) );
  OR2_X2 OR2_10( .ZN(UC_17VZVOR1NF), .A1(C2VCO1), .A2(UC_17) );
  OR2_X1 OR2_11( .ZN(UC_18VZVOR1NF), .A1(C2VCO0), .A2(UC_18) );
  OR2_X1 OR2_12( .ZN(UC_19VZVOR1NF), .A1(C2VIINHN), .A2(UC_19) );
  OR2_X1 OR2_13( .ZN(C3_Q3VZVOR1NF), .A1(C3VCO2), .A2(C3_Q3) );
  OR2_X1 OR2_14( .ZN(C3_Q2VZVOR1NF), .A1(C3VCO1), .A2(C3_Q2) );
  OR2_X1 OR2_15( .ZN(C3_Q1VZVOR1NF), .A1(C3VCO0), .A2(C3_Q1) );
  OR2_X1 OR2_16( .ZN(C3_Q0VZVOR1NF), .A1(C3VIINHN), .A2(C3_Q0) );
  NAND2_X1 NAND2_0( .ZN(TCOMBVNODE18), .A1(TCOMBVNQB), .A2(C3_Q0) );
  NAND4_X1 NAND4_0( .ZN(TCOMBVNODE6), .A1(TCOMBVNFM), .A2(TCOMBVNQD), .A3(TCOMBVNQB), .A4(C3_Q0) );
  NAND2_X1 NAND2_1( .ZN(UC_9VUC_0), .A1(C1VCO1), .A2(UC_9) );
  NAND2_X1 NAND2_2( .ZN(UC_10VUC_0), .A1(C1VCO0), .A2(UC_10) );
  NAND2_X1 NAND2_3( .ZN(TCOMB_RA2), .A1(TCOMB_RA2VOR3NF), .A2(TCOMB_RA2VOR1NF) );
  NAND2_X1 NAND2_4( .ZN(TCOMBVNODE4), .A1(TCOMBVNODE4VOR2NF), .A2(TCOMBVNODE4VOR1NF) );
  NAND2_X1 NAND2_5( .ZN(TCOMBVNODE14), .A1(TCOMBVNODE15), .A2(TCOMBVNQA) );
  NAND4_X1 NAND4_1( .ZN(TCOMBVNODE12), .A1(TCOMBVNCLR), .A2(TCOMBVNFEL), .A3(TCOMBVNQC), .A4(C3_Q1) );
  NAND4_X1 NAND4_2( .ZN(TCOMBVNODE8), .A1(TCOMBVNCLR), .A2(C3_Q2), .A3(TCOMBVNODE8VOR2NF), .A4(TCOMBVNODE8VOR1NF) );
  NAND3_X1 NAND3_0( .ZN(TCOMB_RA1), .A1(TCOMBVNCLR), .A2(TCOMB_RA1VOR2NF), .A3(TCOMB_RA1VOR1NF) );
  NAND2_X1 NAND2_6( .ZN(TCOMBVNODE16), .A1(TCOMBVNODE19), .A2(TCOMBVNODE16VOR1NF) );
  NAND2_X1 NAND2_7( .ZN(UC_9VZ), .A1(UC_9VZVOR1NF), .A2(UC_9VUC_0) );
  NAND2_X1 NAND2_8( .ZN(UC_10VZ), .A1(UC_10VZVOR1NF), .A2(UC_10VUC_0) );
  NAND2_X1 NAND2_9( .ZN(FMLVIINMUXVND1), .A1(FMLVIINMUXVOR2NF), .A2(FMLVIINMUXVOR1NF) );
  NAND3_X1 NAND3_1( .ZN(TCOMBVNODE3), .A1(TCOMBVNODE4), .A2(TCOMBVNQB), .A3(TCOMBVNQA) );
  NAND2_X1 NAND2_10( .ZN(TESTLVIINMUXVND1), .A1(TESTLVIINMUXVOR2NF), .A2(TESTLVIINMUXVOR1NF) );
  NAND2_X1 NAND2_11( .ZN(TCOMB_FE), .A1(TCOMBVNODE16), .A2(TCOMBVNODE14) );
  NAND2_X1 NAND2_12( .ZN(UC_17VUC_0), .A1(C2VCO1), .A2(UC_17) );
  NAND2_X2 NAND2_13( .ZN(UC_18VUC_0), .A1(C2VCO0), .A2(UC_18) );
  NAND2_X2 NAND2_14( .ZN(UC_19VUC_0), .A1(C2VIINHN), .A2(UC_19) );
  NAND2_X2 NAND2_15( .ZN(TCOMB_YA1), .A1(TCOMBVNODE16), .A2(TCOMBVNODE3) );
  NAND2_X2 NAND2_16( .ZN(UC_17VZ), .A1(UC_17VZVOR1NF), .A2(UC_17VUC_0) );
  NAND2_X1 NAND2_17( .ZN(UC_18VZ), .A1(UC_18VZVOR1NF), .A2(UC_18VUC_0) );
  NAND2_X1 NAND2_18( .ZN(UC_19VZ), .A1(UC_19VZVOR1NF), .A2(UC_19VUC_0) );
  NAND2_X1 NAND2_19( .ZN(C3_Q2VUC_0), .A1(C3VCO1), .A2(C3_Q2) );
  NAND2_X1 NAND2_20( .ZN(C3_Q1VUC_0), .A1(C3VCO0), .A2(C3_Q1) );
  NAND2_X1 NAND2_21( .ZN(C3_Q0VUC_0), .A1(C3VIINHN), .A2(C3_Q0) );
  NAND2_X1 NAND2_22( .ZN(C3_Q2VZ), .A1(C3_Q2VZVOR1NF), .A2(C3_Q2VUC_0) );
  NAND2_X1 NAND2_23( .ZN(C3_Q1VZ), .A1(C3_Q1VZVOR1NF), .A2(C3_Q1VUC_0) );
  NAND2_X1 NAND2_24( .ZN(C3_Q0VZ), .A1(C3_Q0VZVOR1NF), .A2(C3_Q0VUC_0) );
  NOR3_X1 NOR3_0( .ZN(C3VCIIA), .A1(C3_Q2), .A2(C3_Q1), .A3(C3_Q0) );
  NOR3_X1 NOR3_1( .ZN(C1VCIIA), .A1(UC_9), .A2(UC_10), .A3(UC_11) );
  NOR3_X1 NOR3_2( .ZN(C2VCIIA), .A1(UC_17), .A2(UC_18), .A3(UC_19) );
  NOR2_X1 NOR2_0( .ZN(C1_CO), .A1(C1VCIIA), .A2(UC_12) );
  NOR3_X1 NOR3_3( .ZN(C1VCO2), .A1(UC_13), .A2(UC_14), .A3(UC_15) );
  NOR2_X1 NOR2_1( .ZN(C1VCO1), .A1(UC_14), .A2(UC_15) );
  NOR2_X1 NOR2_2( .ZN(TCOMBVNODE19), .A1(CLRB), .A2(TCOMBVNFEL) );
  NOR3_X1 NOR4_0_A( .ZN(extra0), .A1(CLRB), .A2(TCOMBVNFM), .A3(TCOMBVNQC) );
  NOR2_X1 NOR4_0( .ZN(TCOMBVNODE15), .A1(extra0), .A2(C3_Q1) );
  NOR2_X1 NOR2_3( .ZN(CTST), .A1(C1_CO), .A2(TESTL) );
  NOR3_X1 NOR3_4( .ZN(UC_11VD), .A1(CLRB), .A2(UC_11VZ), .A3(C1_CO) );
  NOR3_X1 NOR4_1_A( .ZN(extra1), .A1(CTST), .A2(C2_QN2), .A3(UC_21) );
  NOR2_X1 NOR4_1( .ZN(C2VCO2), .A1(extra1), .A2(UC_22) );
  NOR3_X1 NOR3_5( .ZN(C2VCO1), .A1(CTST), .A2(UC_21), .A3(UC_22) );
  NOR3_X1 NOR3_6( .ZN(C2_CO), .A1(C2VCIIA), .A2(CTST), .A3(UC_20) );
  NOR2_X1 NOR2_4( .ZN(C2VCO0), .A1(CTST), .A2(UC_22) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(TCOMB_GA2VAD4NF), .A2(TCOMB_GA2VAD3NF), .A3(TCOMB_GA2VAD2NF) );
  NOR2_X1 NOR4_2( .ZN(TCOMB_GA2), .A1(extra2), .A2(TCOMB_GA2VAD1NF) );
  NOR2_X1 NOR2_5( .ZN(TCOMB_YA2), .A1(TCOMBVNODE12), .A2(TCOMBVNQA) );
  NOR2_X1 NOR2_6( .ZN(TCOMB_GA1), .A1(TCOMBVNODE8), .A2(TCOMB_GA1VAD1NF) );
  NOR3_X2 NOR3_7( .ZN(UC_8VD), .A1(CLRB), .A2(UC_8VZ), .A3(C1_CO) );
  NOR3_X2 NOR3_8( .ZN(UC_9VD), .A1(CLRB), .A2(UC_9VZ), .A3(C1_CO) );
  NOR3_X2 NOR3_9( .ZN(UC_10VD), .A1(CLRB), .A2(UC_10VZ), .A3(C1_CO) );
  NOR3_X2 NOR4_3_A( .ZN(extra3), .A1(CO2), .A2(UC_24), .A3(UC_25) );
  NOR2_X2 NOR4_3( .ZN(C3VCO2), .A1(extra3), .A2(UC_26) );
  NOR3_X1 NOR3_10( .ZN(C3VCO1), .A1(CO2), .A2(UC_25), .A3(UC_26) );
  NOR3_X1 NOR3_11( .ZN(UC_27), .A1(C3VCIIA), .A2(CO2), .A3(UC_23) );
  NOR2_X1 NOR2_7( .ZN(C3VCO0), .A1(CO2), .A2(UC_26) );
  NOR3_X1 NOR3_12( .ZN(UC_16VD), .A1(CLRB), .A2(UC_16VZ), .A3(C2_CO) );
  NOR3_X1 NOR3_13( .ZN(UC_17VD), .A1(CLRB), .A2(UC_17VZ), .A3(C2_CO) );
  NOR3_X1 NOR3_14( .ZN(UC_18VD), .A1(CLRB), .A2(UC_18VZ), .A3(C2_CO) );
  NOR3_X1 NOR3_15( .ZN(UC_19VD), .A1(CLRB), .A2(UC_19VZ), .A3(C2_CO) );
  NOR2_X1 NOR2_8( .ZN(Y1C), .A1(Y1CVAD2NF), .A2(Y1CVAD1NF) );
  NOR2_X1 NOR2_9( .ZN(R2C), .A1(R2CVAD2NF), .A2(R2CVAD1NF) );
  NOR3_X1 NOR3_16( .ZN(C3_Q3VD), .A1(CLRB), .A2(C3_Q3VZ), .A3(UC_27) );
  NOR3_X1 NOR3_17( .ZN(C3_Q2VD), .A1(CLRB), .A2(C3_Q2VZ), .A3(UC_27) );
  NOR3_X1 NOR3_18( .ZN(C3_Q1VD), .A1(CLRB), .A2(C3_Q1VZ), .A3(UC_27) );
  NOR3_X4 NOR3_19( .ZN(C3_Q0VD), .A1(CLRB), .A2(C3_Q0VZ), .A3(UC_27) );

endmodule
