// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module c432(N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,
  N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115,
  N223,N329,N370,N421,N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
  N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115;
output N223,N329,N370,N421,N430,N431,N432;

  wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,N138,N139,N142,N143,N146,N147,
    N150,N151,N154,N157,N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,N184,N185,
    N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N203,N213,
    N224,N227,N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,N254,N255,N256,N257,
    N258,N259,N260,N263,N264,N267,N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
    N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N319,
    N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
    N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,N371,N372,N373,
    N374,N375,N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,N407,N411,N414,N415,
    N416,N417,N418,N419,N420,N422,N425,N428,N429,extra0,extra1,extra2,extra3,extra4,extra5,extra6,
    extra7;

  INV_X1 NOT1_1( .ZN(N118), .A(N1) );
  INV_X1 NOT1_2( .ZN(N119), .A(N4) );
  INV_X1 NOT1_3( .ZN(N122), .A(N11) );
  INV_X1 NOT1_4( .ZN(N123), .A(N17) );
  INV_X1 NOT1_5( .ZN(N126), .A(N24) );
  INV_X1 NOT1_6( .ZN(N127), .A(N30) );
  INV_X2 NOT1_7( .ZN(N130), .A(N37) );
  INV_X2 NOT1_8( .ZN(N131), .A(N43) );
  INV_X2 NOT1_9( .ZN(N134), .A(N50) );
  INV_X2 NOT1_10( .ZN(N135), .A(N56) );
  INV_X1 NOT1_11( .ZN(N138), .A(N63) );
  INV_X1 NOT1_12( .ZN(N139), .A(N69) );
  INV_X1 NOT1_13( .ZN(N142), .A(N76) );
  INV_X1 NOT1_14( .ZN(N143), .A(N82) );
  INV_X1 NOT1_15( .ZN(N146), .A(N89) );
  INV_X1 NOT1_16( .ZN(N147), .A(N95) );
  INV_X1 NOT1_17( .ZN(N150), .A(N102) );
  INV_X1 NOT1_18( .ZN(N151), .A(N108) );
  NAND2_X1 NAND2_19( .ZN(N154), .A1(N118), .A2(N4) );
  NOR2_X1 NOR2_20( .ZN(N157), .A1(N8), .A2(N119) );
  NOR2_X1 NOR2_21( .ZN(N158), .A1(N14), .A2(N119) );
  NAND2_X1 NAND2_22( .ZN(N159), .A1(N122), .A2(N17) );
  NAND2_X1 NAND2_23( .ZN(N162), .A1(N126), .A2(N30) );
  NAND2_X1 NAND2_24( .ZN(N165), .A1(N130), .A2(N43) );
  NAND2_X1 NAND2_25( .ZN(N168), .A1(N134), .A2(N56) );
  NAND2_X1 NAND2_26( .ZN(N171), .A1(N138), .A2(N69) );
  NAND2_X1 NAND2_27( .ZN(N174), .A1(N142), .A2(N82) );
  NAND2_X1 NAND2_28( .ZN(N177), .A1(N146), .A2(N95) );
  NAND2_X1 NAND2_29( .ZN(N180), .A1(N150), .A2(N108) );
  NOR2_X2 NOR2_30( .ZN(N183), .A1(N21), .A2(N123) );
  NOR2_X2 NOR2_31( .ZN(N184), .A1(N27), .A2(N123) );
  NOR2_X2 NOR2_32( .ZN(N185), .A1(N34), .A2(N127) );
  NOR2_X2 NOR2_33( .ZN(N186), .A1(N40), .A2(N127) );
  NOR2_X2 NOR2_34( .ZN(N187), .A1(N47), .A2(N131) );
  NOR2_X1 NOR2_35( .ZN(N188), .A1(N53), .A2(N131) );
  NOR2_X1 NOR2_36( .ZN(N189), .A1(N60), .A2(N135) );
  NOR2_X1 NOR2_37( .ZN(N190), .A1(N66), .A2(N135) );
  NOR2_X1 NOR2_38( .ZN(N191), .A1(N73), .A2(N139) );
  NOR2_X1 NOR2_39( .ZN(N192), .A1(N79), .A2(N139) );
  NOR2_X1 NOR2_40( .ZN(N193), .A1(N86), .A2(N143) );
  NOR2_X1 NOR2_41( .ZN(N194), .A1(N92), .A2(N143) );
  NOR2_X1 NOR2_42( .ZN(N195), .A1(N99), .A2(N147) );
  NOR2_X2 NOR2_43( .ZN(N196), .A1(N105), .A2(N147) );
  NOR2_X2 NOR2_44( .ZN(N197), .A1(N112), .A2(N151) );
  NOR2_X1 NOR2_45( .ZN(N198), .A1(N115), .A2(N151) );
  AND4_X1 AND9_46_A( .ZN(extra0), .A1(N154), .A2(N159), .A3(N162), .A4(N165) );
  AND4_X1 AND9_46_B( .ZN(extra1), .A1(extra0), .A2(N168), .A3(N171), .A4(N174) );
  AND3_X1 AND9_46( .ZN(N199), .A1(extra1), .A2(N177), .A3(N180) );
  INV_X1 NOT1_47( .ZN(N203), .A(N199) );
  INV_X1 NOT1_48( .ZN(N213), .A(N199) );
  INV_X1 NOT1_49( .ZN(N223), .A(N199) );
  XOR2_X1 XOR2_50( .Z(N224), .A(N203), .B(N154) );
  XOR2_X1 XOR2_51( .Z(N227), .A(N203), .B(N159) );
  XOR2_X1 XOR2_52( .Z(N230), .A(N203), .B(N162) );
  XOR2_X1 XOR2_53( .Z(N233), .A(N203), .B(N165) );
  XOR2_X1 XOR2_54( .Z(N236), .A(N203), .B(N168) );
  XOR2_X1 XOR2_55( .Z(N239), .A(N203), .B(N171) );
  NAND2_X1 NAND2_56( .ZN(N242), .A1(N1), .A2(N213) );
  XOR2_X1 XOR2_57( .Z(N243), .A(N203), .B(N174) );
  NAND2_X1 NAND2_58( .ZN(N246), .A1(N213), .A2(N11) );
  XOR2_X1 XOR2_59( .Z(N247), .A(N203), .B(N177) );
  NAND2_X1 NAND2_60( .ZN(N250), .A1(N213), .A2(N24) );
  XOR2_X1 XOR2_61( .Z(N251), .A(N203), .B(N180) );
  NAND2_X1 NAND2_62( .ZN(N254), .A1(N213), .A2(N37) );
  NAND2_X1 NAND2_63( .ZN(N255), .A1(N213), .A2(N50) );
  NAND2_X1 NAND2_64( .ZN(N256), .A1(N213), .A2(N63) );
  NAND2_X1 NAND2_65( .ZN(N257), .A1(N213), .A2(N76) );
  NAND2_X1 NAND2_66( .ZN(N258), .A1(N213), .A2(N89) );
  NAND2_X1 NAND2_67( .ZN(N259), .A1(N213), .A2(N102) );
  NAND2_X1 NAND2_68( .ZN(N260), .A1(N224), .A2(N157) );
  NAND2_X1 NAND2_69( .ZN(N263), .A1(N224), .A2(N158) );
  NAND2_X1 NAND2_70( .ZN(N264), .A1(N227), .A2(N183) );
  NAND2_X2 NAND2_71( .ZN(N267), .A1(N230), .A2(N185) );
  NAND2_X2 NAND2_72( .ZN(N270), .A1(N233), .A2(N187) );
  NAND2_X2 NAND2_73( .ZN(N273), .A1(N236), .A2(N189) );
  NAND2_X2 NAND2_74( .ZN(N276), .A1(N239), .A2(N191) );
  NAND2_X2 NAND2_75( .ZN(N279), .A1(N243), .A2(N193) );
  NAND2_X2 NAND2_76( .ZN(N282), .A1(N247), .A2(N195) );
  NAND2_X2 NAND2_77( .ZN(N285), .A1(N251), .A2(N197) );
  NAND2_X1 NAND2_78( .ZN(N288), .A1(N227), .A2(N184) );
  NAND2_X1 NAND2_79( .ZN(N289), .A1(N230), .A2(N186) );
  NAND2_X1 NAND2_80( .ZN(N290), .A1(N233), .A2(N188) );
  NAND2_X1 NAND2_81( .ZN(N291), .A1(N236), .A2(N190) );
  NAND2_X1 NAND2_82( .ZN(N292), .A1(N239), .A2(N192) );
  NAND2_X1 NAND2_83( .ZN(N293), .A1(N243), .A2(N194) );
  NAND2_X1 NAND2_84( .ZN(N294), .A1(N247), .A2(N196) );
  NAND2_X1 NAND2_85( .ZN(N295), .A1(N251), .A2(N198) );
  AND4_X1 AND9_86_A( .ZN(extra2), .A1(N260), .A2(N264), .A3(N267), .A4(N270) );
  AND4_X1 AND9_86_B( .ZN(extra3), .A1(extra2), .A2(N273), .A3(N276), .A4(N279) );
  AND3_X1 AND9_86( .ZN(N296), .A1(extra3), .A2(N282), .A3(N285) );
  INV_X1 NOT1_87( .ZN(N300), .A(N263) );
  INV_X1 NOT1_88( .ZN(N301), .A(N288) );
  INV_X1 NOT1_89( .ZN(N302), .A(N289) );
  INV_X2 NOT1_90( .ZN(N303), .A(N290) );
  INV_X2 NOT1_91( .ZN(N304), .A(N291) );
  INV_X2 NOT1_92( .ZN(N305), .A(N292) );
  INV_X1 NOT1_93( .ZN(N306), .A(N293) );
  INV_X1 NOT1_94( .ZN(N307), .A(N294) );
  INV_X1 NOT1_95( .ZN(N308), .A(N295) );
  INV_X1 NOT1_96( .ZN(N309), .A(N296) );
  INV_X1 NOT1_97( .ZN(N319), .A(N296) );
  INV_X1 NOT1_98( .ZN(N329), .A(N296) );
  XOR2_X1 XOR2_99( .Z(N330), .A(N309), .B(N260) );
  XOR2_X1 XOR2_100( .Z(N331), .A(N309), .B(N264) );
  XOR2_X1 XOR2_101( .Z(N332), .A(N309), .B(N267) );
  XOR2_X1 XOR2_102( .Z(N333), .A(N309), .B(N270) );
  NAND2_X1 NAND2_103( .ZN(N334), .A1(N8), .A2(N319) );
  XOR2_X1 XOR2_104( .Z(N335), .A(N309), .B(N273) );
  NAND2_X1 NAND2_105( .ZN(N336), .A1(N319), .A2(N21) );
  XOR2_X1 XOR2_106( .Z(N337), .A(N309), .B(N276) );
  NAND2_X1 NAND2_107( .ZN(N338), .A1(N319), .A2(N34) );
  XOR2_X1 XOR2_108( .Z(N339), .A(N309), .B(N279) );
  NAND2_X1 NAND2_109( .ZN(N340), .A1(N319), .A2(N47) );
  XOR2_X1 XOR2_110( .Z(N341), .A(N309), .B(N282) );
  NAND2_X1 NAND2_111( .ZN(N342), .A1(N319), .A2(N60) );
  XOR2_X1 XOR2_112( .Z(N343), .A(N309), .B(N285) );
  NAND2_X1 NAND2_113( .ZN(N344), .A1(N319), .A2(N73) );
  NAND2_X1 NAND2_114( .ZN(N345), .A1(N319), .A2(N86) );
  NAND2_X1 NAND2_115( .ZN(N346), .A1(N319), .A2(N99) );
  NAND2_X1 NAND2_116( .ZN(N347), .A1(N319), .A2(N112) );
  NAND2_X1 NAND2_117( .ZN(N348), .A1(N330), .A2(N300) );
  NAND2_X2 NAND2_118( .ZN(N349), .A1(N331), .A2(N301) );
  NAND2_X4 NAND2_119( .ZN(N350), .A1(N332), .A2(N302) );
  NAND2_X2 NAND2_120( .ZN(N351), .A1(N333), .A2(N303) );
  NAND2_X1 NAND2_121( .ZN(N352), .A1(N335), .A2(N304) );
  NAND2_X1 NAND2_122( .ZN(N353), .A1(N337), .A2(N305) );
  NAND2_X1 NAND2_123( .ZN(N354), .A1(N339), .A2(N306) );
  NAND2_X1 NAND2_124( .ZN(N355), .A1(N341), .A2(N307) );
  NAND2_X1 NAND2_125( .ZN(N356), .A1(N343), .A2(N308) );
  AND4_X1 AND9_126_A( .ZN(extra4), .A1(N348), .A2(N349), .A3(N350), .A4(N351) );
  AND4_X1 AND9_126_B( .ZN(extra5), .A1(extra4), .A2(N352), .A3(N353), .A4(N354) );
  AND3_X1 AND9_126( .ZN(N357), .A1(extra5), .A2(N355), .A3(N356) );
  INV_X1 NOT1_127( .ZN(N360), .A(N357) );
  INV_X1 NOT1_128( .ZN(N370), .A(N357) );
  NAND2_X1 NAND2_129( .ZN(N371), .A1(N14), .A2(N360) );
  NAND2_X1 NAND2_130( .ZN(N372), .A1(N360), .A2(N27) );
  NAND2_X1 NAND2_131( .ZN(N373), .A1(N360), .A2(N40) );
  NAND2_X2 NAND2_132( .ZN(N374), .A1(N360), .A2(N53) );
  NAND2_X1 NAND2_133( .ZN(N375), .A1(N360), .A2(N66) );
  NAND2_X1 NAND2_134( .ZN(N376), .A1(N360), .A2(N79) );
  NAND2_X2 NAND2_135( .ZN(N377), .A1(N360), .A2(N92) );
  NAND2_X2 NAND2_136( .ZN(N378), .A1(N360), .A2(N105) );
  NAND2_X2 NAND2_137( .ZN(N379), .A1(N360), .A2(N115) );
  NAND4_X1 NAND4_138( .ZN(N380), .A1(N4), .A2(N242), .A3(N334), .A4(N371) );
  NAND4_X1 NAND4_139( .ZN(N381), .A1(N246), .A2(N336), .A3(N372), .A4(N17) );
  NAND4_X1 NAND4_140( .ZN(N386), .A1(N250), .A2(N338), .A3(N373), .A4(N30) );
  NAND4_X1 NAND4_141( .ZN(N393), .A1(N254), .A2(N340), .A3(N374), .A4(N43) );
  NAND4_X1 NAND4_142( .ZN(N399), .A1(N255), .A2(N342), .A3(N375), .A4(N56) );
  NAND4_X1 NAND4_143( .ZN(N404), .A1(N256), .A2(N344), .A3(N376), .A4(N69) );
  NAND4_X1 NAND4_144( .ZN(N407), .A1(N257), .A2(N345), .A3(N377), .A4(N82) );
  NAND4_X1 NAND4_145( .ZN(N411), .A1(N258), .A2(N346), .A3(N378), .A4(N95) );
  NAND4_X1 NAND4_146( .ZN(N414), .A1(N259), .A2(N347), .A3(N379), .A4(N108) );
  INV_X1 NOT1_147( .ZN(N415), .A(N380) );
  AND4_X1 AND8_148_A( .ZN(extra6), .A1(N381), .A2(N386), .A3(N393), .A4(N399) );
  AND4_X2 AND8_148_B( .ZN(extra7), .A1(extra6), .A2(N404), .A3(N407), .A4(N411) );
  AND2_X4 AND8_148( .ZN(N416), .A1(extra7), .A2(N414) );
  INV_X1 NOT1_149( .ZN(N417), .A(N393) );
  INV_X1 NOT1_150( .ZN(N418), .A(N404) );
  INV_X1 NOT1_151( .ZN(N419), .A(N407) );
  INV_X1 NOT1_152( .ZN(N420), .A(N411) );
  NOR2_X2 NOR2_153( .ZN(N421), .A1(N415), .A2(N416) );
  NAND2_X1 NAND2_154( .ZN(N422), .A1(N386), .A2(N417) );
  NAND4_X1 NAND4_155( .ZN(N425), .A1(N386), .A2(N393), .A3(N418), .A4(N399) );
  NAND3_X1 NAND3_156( .ZN(N428), .A1(N399), .A2(N393), .A3(N419) );
  NAND4_X2 NAND4_157( .ZN(N429), .A1(N386), .A2(N393), .A3(N407), .A4(N420) );
  NAND4_X2 NAND4_158( .ZN(N430), .A1(N381), .A2(N386), .A3(N422), .A4(N399) );
  NAND4_X1 NAND4_159( .ZN(N431), .A1(N381), .A2(N386), .A3(N425), .A4(N428) );
  NAND4_X1 NAND4_160( .ZN(N432), .A1(N381), .A2(N422), .A3(N425), .A4(N429) );

endmodule
