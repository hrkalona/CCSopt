// Verilog
// c2670
// Ninputs 233
// Noutputs 140
// NtotalGates 1269
// BUFF1 272
// AND2 203
// NOT1 321
// AND4 11
// AND3 112
// NAND2 254
// OR2 51
// OR4 22
// NOR2 12
// AND5 7
// OR3 2
// OR5 2

module c2670(N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,
  N51,N52,N53,N54,N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N135,N136,
  N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,N237,N241,N246,N253,N256,N259,
  N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,N305,N309,N313,N316,
  N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,N146_I,N147_I,
  N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
  N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,
  N184_I,N185_I,N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,
  N202_I,N203_I,N204_I,N205_I,N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I,N398,
  N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,
  N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
  N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,
  N3546,N3671,N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,
  N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,
  N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,
  N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
  N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O);
input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
  N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
  N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
  N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
  N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
  N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
  N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
  N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
  N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,N216_I,N217_I,N218_I;
output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
  N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
  N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
  N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
  N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
  N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
  N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;

  wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,N506,N509,N521,N533,N537,N543,
    N544,N547,N550,N562,N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,N612,N613,
    N625,N637,N643,N650,N651,N655,N659,N663,N667,N671,N675,N679,N683,N687,N693,N699,
    N705,N711,N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,N744,N747,N750,N753,
    N756,N759,N762,N765,N768,N771,N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
    N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,N1053,N1064,N1065,N1066,N1067,N1068,
    N1069,N1070,N1075,N1086,N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,N1127,N1128,
    N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,
    N1173,N1178,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,N1210,N1211,N1212,N1213,
    N1214,N1215,N1216,N1219,N1222,N1225,N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
    N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,N1353,N1354,N1355,N1395,N1396,N1397,
    N1398,N1399,N1422,N1423,N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,N1453,N1454,
    N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,
    N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,
    N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
    N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,
    N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,
    N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
    N1575,N1576,N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,N1612,N1615,N1619,N1624,
    N1628,N1631,N1634,N1637,N1642,N1647,N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
    N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,N1808,N1809,N1810,N1811,N1813,N1814,
    N1815,N1822,N1823,N1824,N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,N1863,N1870,
    N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,
    N1917,N1918,N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1939,N1940,N1941,N1942,
    N1945,N1948,N1951,N1954,N1957,N1960,N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
    N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,N2067,N2070,N2073,N2076,N2079,N2095,
    N2098,N2101,N2104,N2107,N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,N2144,N2147,
    N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,
    N2188,N2191,N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,N2234,N2235,N2236,N2237,
    N2250,N2266,N2269,N2291,N2294,N2297,N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
    N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,
    N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,
    N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,
    N2377,N2382,N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,
    N2415,N2416,N2417,N2421,N2425,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
    N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,N2475,N2478,N2481,N2484,N2487,N2490,
    N2493,N2503,N2504,N2510,N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,N2547,N2548,
    N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,
    N2610,N2611,N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,N2630,N2631,N2632,N2633,
    N2634,N2635,N2636,N2638,N2645,N2646,N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
    N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2684,N2687,N2690,
    N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,N2709,N2710,
    N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,
    N2773,N2774,N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,N2791,N2792,N2793,N2796,
    N2800,N2803,N2806,N2809,N2810,N2811,N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
    N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,N2882,N2885,N2888,N2894,N2895,N2896,
    N2897,N2898,N2899,N2900,N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,N2938,N2939,
    N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,
    N3009,N3010,N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,N3037,N3039,N3044,N3045,
    N3046,N3047,N3048,N3049,N3050,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
    N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3088,N3091,N3110,N3113,N3137,
    N3140,N3143,N3146,N3149,N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,N3178,N3180,
    N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,
    N3219,N3220,N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,N3256,N3259,N3262,N3265,
    N3268,N3271,N3274,N3277,N3281,N3282,N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
    N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,N3321,N3324,N3327,N3330,N3333,N3334,
    N3335,N3336,N3337,N3340,N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,N3382,N3386,
    N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,
    N3420,N3422,N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,N3459,N3478,N3479,N3480,
    N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
    N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3515,
    N3517,N3522,N3525,N3528,N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
    N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,
    N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,N3622,N3629,N3630,N3631,
    N3632,N3633,N3634,N3635,N3640,N3644,N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
    N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3726,N3727,
    N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,N3744,N3745,
    N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,
    N3780,N3790,N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,N3814,N3815,N3816,N3817,
    N3818,N3819,N3820,N3821,N3822,N3823,N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
    N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877,extra0,extra1,extra2,extra3,extra4,extra5,extra6,
    extra7,extra8;

  BUF_X1 BUFF1_1( .Z(N398), .A(N219) );
  BUF_X2 BUFF1_2( .Z(N400), .A(N219) );
  BUF_X1 BUFF1_3( .Z(N401), .A(N219) );
  AND2_X1 AND2_4( .ZN(N405), .A1(N1), .A2(N3) );
  INV_X2 NOT1_5( .ZN(N408), .A(N230) );
  BUF_X1 BUFF1_6( .Z(N419), .A(N253) );
  BUF_X1 BUFF1_7( .Z(N420), .A(N253) );
  INV_X1 NOT1_8( .ZN(N425), .A(N262) );
  BUF_X1 BUFF1_9( .Z(N456), .A(N290) );
  BUF_X1 BUFF1_10( .Z(N457), .A(N290) );
  BUF_X1 BUFF1_11( .Z(N458), .A(N290) );
  AND4_X1 AND4_12( .ZN(N485), .A1(N309), .A2(N305), .A3(N301), .A4(N297) );
  INV_X1 NOT1_13( .ZN(N486), .A(N405) );
  INV_X1 NOT1_14( .ZN(N487), .A(N44) );
  INV_X1 NOT1_15( .ZN(N488), .A(N132) );
  INV_X1 NOT1_16( .ZN(N489), .A(N82) );
  INV_X1 NOT1_17( .ZN(N490), .A(N96) );
  INV_X1 NOT1_18( .ZN(N491), .A(N69) );
  INV_X1 NOT1_19( .ZN(N492), .A(N120) );
  INV_X1 NOT1_20( .ZN(N493), .A(N57) );
  INV_X1 NOT1_21( .ZN(N494), .A(N108) );
  AND3_X1 AND3_22( .ZN(N495), .A1(N2), .A2(N15), .A3(N237) );
  BUF_X1 BUFF1_23( .Z(N496), .A(N237) );
  AND2_X2 AND2_24( .ZN(N499), .A1(N37), .A2(N37) );
  BUF_X1 BUFF1_25( .Z(N500), .A(N219) );
  BUF_X1 BUFF1_26( .Z(N503), .A(N8) );
  BUF_X1 BUFF1_27( .Z(N506), .A(N8) );
  BUF_X1 BUFF1_28( .Z(N509), .A(N227) );
  BUF_X1 BUFF1_29( .Z(N521), .A(N234) );
  INV_X1 NOT1_30( .ZN(N533), .A(N241) );
  INV_X1 NOT1_31( .ZN(N537), .A(N246) );
  AND2_X1 AND2_32( .ZN(N543), .A1(N11), .A2(N246) );
  AND4_X1 AND4_33( .ZN(N544), .A1(N132), .A2(N82), .A3(N96), .A4(N44) );
  AND4_X1 AND4_34( .ZN(N547), .A1(N120), .A2(N57), .A3(N108), .A4(N69) );
  BUF_X1 BUFF1_35( .Z(N550), .A(N227) );
  BUF_X1 BUFF1_36( .Z(N562), .A(N234) );
  INV_X1 NOT1_37( .ZN(N574), .A(N256) );
  INV_X1 NOT1_38( .ZN(N578), .A(N259) );
  BUF_X1 BUFF1_39( .Z(N582), .A(N319) );
  BUF_X1 BUFF1_40( .Z(N594), .A(N322) );
  INV_X1 NOT1_41( .ZN(N606), .A(N328) );
  INV_X1 NOT1_42( .ZN(N607), .A(N331) );
  INV_X1 NOT1_43( .ZN(N608), .A(N334) );
  INV_X1 NOT1_44( .ZN(N609), .A(N337) );
  INV_X1 NOT1_45( .ZN(N610), .A(N340) );
  INV_X1 NOT1_46( .ZN(N611), .A(N343) );
  INV_X1 NOT1_47( .ZN(N612), .A(N352) );
  BUF_X1 BUFF1_48( .Z(N613), .A(N319) );
  BUF_X1 BUFF1_49( .Z(N625), .A(N322) );
  BUF_X1 BUFF1_50( .Z(N637), .A(N16) );
  BUF_X1 BUFF1_51( .Z(N643), .A(N16) );
  INV_X1 NOT1_52( .ZN(N650), .A(N355) );
  AND2_X1 AND2_53( .ZN(N651), .A1(N7), .A2(N237) );
  INV_X1 NOT1_54( .ZN(N655), .A(N263) );
  INV_X1 NOT1_55( .ZN(N659), .A(N266) );
  INV_X1 NOT1_56( .ZN(N663), .A(N269) );
  INV_X1 NOT1_57( .ZN(N667), .A(N272) );
  INV_X1 NOT1_58( .ZN(N671), .A(N275) );
  INV_X1 NOT1_59( .ZN(N675), .A(N278) );
  INV_X1 NOT1_60( .ZN(N679), .A(N281) );
  INV_X1 NOT1_61( .ZN(N683), .A(N284) );
  INV_X1 NOT1_62( .ZN(N687), .A(N287) );
  BUF_X1 BUFF1_63( .Z(N693), .A(N29) );
  BUF_X1 BUFF1_64( .Z(N699), .A(N29) );
  INV_X1 NOT1_65( .ZN(N705), .A(N294) );
  INV_X1 NOT1_66( .ZN(N711), .A(N297) );
  INV_X1 NOT1_67( .ZN(N715), .A(N301) );
  INV_X1 NOT1_68( .ZN(N719), .A(N305) );
  INV_X1 NOT1_69( .ZN(N723), .A(N309) );
  INV_X1 NOT1_70( .ZN(N727), .A(N313) );
  INV_X1 NOT1_71( .ZN(N730), .A(N316) );
  INV_X1 NOT1_72( .ZN(N733), .A(N346) );
  INV_X1 NOT1_73( .ZN(N734), .A(N349) );
  BUF_X1 BUFF1_74( .Z(N735), .A(N259) );
  BUF_X1 BUFF1_75( .Z(N738), .A(N256) );
  BUF_X1 BUFF1_76( .Z(N741), .A(N263) );
  BUF_X1 BUFF1_77( .Z(N744), .A(N269) );
  BUF_X1 BUFF1_78( .Z(N747), .A(N266) );
  BUF_X1 BUFF1_79( .Z(N750), .A(N275) );
  BUF_X1 BUFF1_80( .Z(N753), .A(N272) );
  BUF_X1 BUFF1_81( .Z(N756), .A(N281) );
  BUF_X1 BUFF1_82( .Z(N759), .A(N278) );
  BUF_X1 BUFF1_83( .Z(N762), .A(N287) );
  BUF_X1 BUFF1_84( .Z(N765), .A(N284) );
  BUF_X1 BUFF1_85( .Z(N768), .A(N294) );
  BUF_X1 BUFF1_86( .Z(N771), .A(N301) );
  BUF_X1 BUFF1_87( .Z(N774), .A(N297) );
  BUF_X1 BUFF1_88( .Z(N777), .A(N309) );
  BUF_X1 BUFF1_89( .Z(N780), .A(N305) );
  BUF_X1 BUFF1_90( .Z(N783), .A(N316) );
  BUF_X1 BUFF1_91( .Z(N786), .A(N313) );
  INV_X1 NOT1_92( .ZN(N792), .A(N485) );
  INV_X1 NOT1_93( .ZN(N799), .A(N495) );
  INV_X1 NOT1_94( .ZN(N800), .A(N499) );
  BUF_X1 BUFF1_95( .Z(N805), .A(N500) );
  NAND2_X2 NAND2_96( .ZN(N900), .A1(N331), .A2(N606) );
  NAND2_X1 NAND2_97( .ZN(N901), .A1(N328), .A2(N607) );
  NAND2_X1 NAND2_98( .ZN(N902), .A1(N337), .A2(N608) );
  NAND2_X1 NAND2_99( .ZN(N903), .A1(N334), .A2(N609) );
  NAND2_X1 NAND2_100( .ZN(N904), .A1(N343), .A2(N610) );
  NAND2_X1 NAND2_101( .ZN(N905), .A1(N340), .A2(N611) );
  NAND2_X1 NAND2_102( .ZN(N998), .A1(N349), .A2(N733) );
  NAND2_X1 NAND2_103( .ZN(N999), .A1(N346), .A2(N734) );
  AND2_X1 AND2_104( .ZN(N1026), .A1(N94), .A2(N500) );
  AND2_X1 AND2_105( .ZN(N1027), .A1(N325), .A2(N651) );
  INV_X1 NOT1_106( .ZN(N1028), .A(N651) );
  NAND2_X1 NAND2_107( .ZN(N1029), .A1(N231), .A2(N651) );
  INV_X1 NOT1_108( .ZN(N1032), .A(N544) );
  INV_X2 NOT1_109( .ZN(N1033), .A(N547) );
  AND2_X1 AND2_110( .ZN(N1034), .A1(N547), .A2(N544) );
  BUF_X2 BUFF1_111( .Z(N1037), .A(N503) );
  INV_X1 NOT1_112( .ZN(N1042), .A(N509) );
  INV_X1 NOT1_113( .ZN(N1053), .A(N521) );
  AND3_X1 AND3_114( .ZN(N1064), .A1(N80), .A2(N509), .A3(N521) );
  AND3_X1 AND3_115( .ZN(N1065), .A1(N68), .A2(N509), .A3(N521) );
  AND3_X1 AND3_116( .ZN(N1066), .A1(N79), .A2(N509), .A3(N521) );
  AND3_X1 AND3_117( .ZN(N1067), .A1(N78), .A2(N509), .A3(N521) );
  AND3_X1 AND3_118( .ZN(N1068), .A1(N77), .A2(N509), .A3(N521) );
  AND2_X1 AND2_119( .ZN(N1069), .A1(N11), .A2(N537) );
  BUF_X2 BUFF1_120( .Z(N1070), .A(N503) );
  INV_X1 NOT1_121( .ZN(N1075), .A(N550) );
  INV_X1 NOT1_122( .ZN(N1086), .A(N562) );
  AND3_X1 AND3_123( .ZN(N1097), .A1(N76), .A2(N550), .A3(N562) );
  AND3_X1 AND3_124( .ZN(N1098), .A1(N75), .A2(N550), .A3(N562) );
  AND3_X1 AND3_125( .ZN(N1099), .A1(N74), .A2(N550), .A3(N562) );
  AND3_X1 AND3_126( .ZN(N1100), .A1(N73), .A2(N550), .A3(N562) );
  AND3_X1 AND3_127( .ZN(N1101), .A1(N72), .A2(N550), .A3(N562) );
  INV_X1 NOT1_128( .ZN(N1102), .A(N582) );
  INV_X1 NOT1_129( .ZN(N1113), .A(N594) );
  AND3_X1 AND3_130( .ZN(N1124), .A1(N114), .A2(N582), .A3(N594) );
  AND3_X1 AND3_131( .ZN(N1125), .A1(N113), .A2(N582), .A3(N594) );
  AND3_X1 AND3_132( .ZN(N1126), .A1(N112), .A2(N582), .A3(N594) );
  AND3_X1 AND3_133( .ZN(N1127), .A1(N111), .A2(N582), .A3(N594) );
  AND2_X1 AND2_134( .ZN(N1128), .A1(N582), .A2(N594) );
  NAND2_X1 NAND2_135( .ZN(N1129), .A1(N900), .A2(N901) );
  NAND2_X1 NAND2_136( .ZN(N1133), .A1(N902), .A2(N903) );
  NAND2_X1 NAND2_137( .ZN(N1137), .A1(N904), .A2(N905) );
  INV_X1 NOT1_138( .ZN(N1140), .A(N741) );
  NAND2_X1 NAND2_139( .ZN(N1141), .A1(N741), .A2(N612) );
  INV_X1 NOT1_140( .ZN(N1142), .A(N744) );
  INV_X1 NOT1_141( .ZN(N1143), .A(N747) );
  INV_X1 NOT1_142( .ZN(N1144), .A(N750) );
  INV_X1 NOT1_143( .ZN(N1145), .A(N753) );
  INV_X1 NOT1_144( .ZN(N1146), .A(N613) );
  INV_X1 NOT1_145( .ZN(N1157), .A(N625) );
  AND3_X1 AND3_146( .ZN(N1168), .A1(N118), .A2(N613), .A3(N625) );
  AND3_X1 AND3_147( .ZN(N1169), .A1(N107), .A2(N613), .A3(N625) );
  AND3_X1 AND3_148( .ZN(N1170), .A1(N117), .A2(N613), .A3(N625) );
  AND3_X1 AND3_149( .ZN(N1171), .A1(N116), .A2(N613), .A3(N625) );
  AND3_X1 AND3_150( .ZN(N1172), .A1(N115), .A2(N613), .A3(N625) );
  INV_X1 NOT1_151( .ZN(N1173), .A(N637) );
  INV_X1 NOT1_152( .ZN(N1178), .A(N643) );
  INV_X1 NOT1_153( .ZN(N1184), .A(N768) );
  NAND2_X1 NAND2_154( .ZN(N1185), .A1(N768), .A2(N650) );
  INV_X1 NOT1_155( .ZN(N1186), .A(N771) );
  INV_X1 NOT1_156( .ZN(N1187), .A(N774) );
  INV_X1 NOT1_157( .ZN(N1188), .A(N777) );
  INV_X1 NOT1_158( .ZN(N1189), .A(N780) );
  BUF_X1 BUFF1_159( .Z(N1190), .A(N506) );
  BUF_X1 BUFF1_160( .Z(N1195), .A(N506) );
  INV_X1 NOT1_161( .ZN(N1200), .A(N693) );
  INV_X1 NOT1_162( .ZN(N1205), .A(N699) );
  INV_X1 NOT1_163( .ZN(N1210), .A(N735) );
  INV_X1 NOT1_164( .ZN(N1211), .A(N738) );
  INV_X1 NOT1_165( .ZN(N1212), .A(N756) );
  INV_X1 NOT1_166( .ZN(N1213), .A(N759) );
  INV_X1 NOT1_167( .ZN(N1214), .A(N762) );
  INV_X1 NOT1_168( .ZN(N1215), .A(N765) );
  NAND2_X1 NAND2_169( .ZN(N1216), .A1(N998), .A2(N999) );
  BUF_X1 BUFF1_170( .Z(N1219), .A(N574) );
  BUF_X1 BUFF1_171( .Z(N1222), .A(N578) );
  BUF_X1 BUFF1_172( .Z(N1225), .A(N655) );
  BUF_X1 BUFF1_173( .Z(N1228), .A(N659) );
  BUF_X1 BUFF1_174( .Z(N1231), .A(N663) );
  BUF_X1 BUFF1_175( .Z(N1234), .A(N667) );
  BUF_X1 BUFF1_176( .Z(N1237), .A(N671) );
  BUF_X1 BUFF1_177( .Z(N1240), .A(N675) );
  BUF_X1 BUFF1_178( .Z(N1243), .A(N679) );
  BUF_X1 BUFF1_179( .Z(N1246), .A(N683) );
  INV_X1 NOT1_180( .ZN(N1249), .A(N783) );
  INV_X1 NOT1_181( .ZN(N1250), .A(N786) );
  BUF_X1 BUFF1_182( .Z(N1251), .A(N687) );
  BUF_X1 BUFF1_183( .Z(N1254), .A(N705) );
  BUF_X1 BUFF1_184( .Z(N1257), .A(N711) );
  BUF_X1 BUFF1_185( .Z(N1260), .A(N715) );
  BUF_X1 BUFF1_186( .Z(N1263), .A(N719) );
  BUF_X1 BUFF1_187( .Z(N1266), .A(N723) );
  INV_X1 NOT1_188( .ZN(N1269), .A(N1027) );
  AND2_X2 AND2_189( .ZN(N1275), .A1(N325), .A2(N1032) );
  AND2_X1 AND2_190( .ZN(N1276), .A1(N231), .A2(N1033) );
  BUF_X1 BUFF1_191( .Z(N1277), .A(N1034) );
  OR2_X1 OR2_192( .ZN(N1302), .A1(N1069), .A2(N543) );
  NAND2_X1 NAND2_193( .ZN(N1351), .A1(N352), .A2(N1140) );
  NAND2_X2 NAND2_194( .ZN(N1352), .A1(N747), .A2(N1142) );
  NAND2_X2 NAND2_195( .ZN(N1353), .A1(N744), .A2(N1143) );
  NAND2_X2 NAND2_196( .ZN(N1354), .A1(N753), .A2(N1144) );
  NAND2_X2 NAND2_197( .ZN(N1355), .A1(N750), .A2(N1145) );
  NAND2_X2 NAND2_198( .ZN(N1395), .A1(N355), .A2(N1184) );
  NAND2_X2 NAND2_199( .ZN(N1396), .A1(N774), .A2(N1186) );
  NAND2_X1 NAND2_200( .ZN(N1397), .A1(N771), .A2(N1187) );
  NAND2_X1 NAND2_201( .ZN(N1398), .A1(N780), .A2(N1188) );
  NAND2_X1 NAND2_202( .ZN(N1399), .A1(N777), .A2(N1189) );
  NAND2_X1 NAND2_203( .ZN(N1422), .A1(N738), .A2(N1210) );
  NAND2_X1 NAND2_204( .ZN(N1423), .A1(N735), .A2(N1211) );
  NAND2_X1 NAND2_205( .ZN(N1424), .A1(N759), .A2(N1212) );
  NAND2_X1 NAND2_206( .ZN(N1425), .A1(N756), .A2(N1213) );
  NAND2_X1 NAND2_207( .ZN(N1426), .A1(N765), .A2(N1214) );
  NAND2_X1 NAND2_208( .ZN(N1427), .A1(N762), .A2(N1215) );
  NAND2_X1 NAND2_209( .ZN(N1440), .A1(N786), .A2(N1249) );
  NAND2_X1 NAND2_210( .ZN(N1441), .A1(N783), .A2(N1250) );
  INV_X2 NOT1_211( .ZN(N1448), .A(N1034) );
  INV_X2 NOT1_212( .ZN(N1449), .A(N1275) );
  INV_X1 NOT1_213( .ZN(N1450), .A(N1276) );
  AND3_X1 AND3_214( .ZN(N1451), .A1(N93), .A2(N1042), .A3(N1053) );
  AND3_X1 AND3_215( .ZN(N1452), .A1(N55), .A2(N509), .A3(N1053) );
  AND3_X1 AND3_216( .ZN(N1453), .A1(N67), .A2(N1042), .A3(N521) );
  AND3_X1 AND3_217( .ZN(N1454), .A1(N81), .A2(N1042), .A3(N1053) );
  AND3_X1 AND3_218( .ZN(N1455), .A1(N43), .A2(N509), .A3(N1053) );
  AND3_X1 AND3_219( .ZN(N1456), .A1(N56), .A2(N1042), .A3(N521) );
  AND3_X1 AND3_220( .ZN(N1457), .A1(N92), .A2(N1042), .A3(N1053) );
  AND3_X1 AND3_221( .ZN(N1458), .A1(N54), .A2(N509), .A3(N1053) );
  AND3_X1 AND3_222( .ZN(N1459), .A1(N66), .A2(N1042), .A3(N521) );
  AND3_X1 AND3_223( .ZN(N1460), .A1(N91), .A2(N1042), .A3(N1053) );
  AND3_X1 AND3_224( .ZN(N1461), .A1(N53), .A2(N509), .A3(N1053) );
  AND3_X1 AND3_225( .ZN(N1462), .A1(N65), .A2(N1042), .A3(N521) );
  AND3_X1 AND3_226( .ZN(N1463), .A1(N90), .A2(N1042), .A3(N1053) );
  AND3_X1 AND3_227( .ZN(N1464), .A1(N52), .A2(N509), .A3(N1053) );
  AND3_X1 AND3_228( .ZN(N1465), .A1(N64), .A2(N1042), .A3(N521) );
  AND3_X1 AND3_229( .ZN(N1466), .A1(N89), .A2(N1075), .A3(N1086) );
  AND3_X1 AND3_230( .ZN(N1467), .A1(N51), .A2(N550), .A3(N1086) );
  AND3_X1 AND3_231( .ZN(N1468), .A1(N63), .A2(N1075), .A3(N562) );
  AND3_X1 AND3_232( .ZN(N1469), .A1(N88), .A2(N1075), .A3(N1086) );
  AND3_X1 AND3_233( .ZN(N1470), .A1(N50), .A2(N550), .A3(N1086) );
  AND3_X1 AND3_234( .ZN(N1471), .A1(N62), .A2(N1075), .A3(N562) );
  AND3_X1 AND3_235( .ZN(N1472), .A1(N87), .A2(N1075), .A3(N1086) );
  AND3_X1 AND3_236( .ZN(N1473), .A1(N49), .A2(N550), .A3(N1086) );
  AND2_X1 AND2_237( .ZN(N1474), .A1(N1075), .A2(N562) );
  AND3_X1 AND3_238( .ZN(N1475), .A1(N86), .A2(N1075), .A3(N1086) );
  AND3_X1 AND3_239( .ZN(N1476), .A1(N48), .A2(N550), .A3(N1086) );
  AND3_X1 AND3_240( .ZN(N1477), .A1(N61), .A2(N1075), .A3(N562) );
  AND3_X1 AND3_241( .ZN(N1478), .A1(N85), .A2(N1075), .A3(N1086) );
  AND3_X1 AND3_242( .ZN(N1479), .A1(N47), .A2(N550), .A3(N1086) );
  AND3_X1 AND3_243( .ZN(N1480), .A1(N60), .A2(N1075), .A3(N562) );
  AND3_X1 AND3_244( .ZN(N1481), .A1(N138), .A2(N1102), .A3(N1113) );
  AND3_X1 AND3_245( .ZN(N1482), .A1(N102), .A2(N582), .A3(N1113) );
  AND3_X1 AND3_246( .ZN(N1483), .A1(N126), .A2(N1102), .A3(N594) );
  AND3_X1 AND3_247( .ZN(N1484), .A1(N137), .A2(N1102), .A3(N1113) );
  AND3_X1 AND3_248( .ZN(N1485), .A1(N101), .A2(N582), .A3(N1113) );
  AND3_X1 AND3_249( .ZN(N1486), .A1(N125), .A2(N1102), .A3(N594) );
  AND3_X1 AND3_250( .ZN(N1487), .A1(N136), .A2(N1102), .A3(N1113) );
  AND3_X1 AND3_251( .ZN(N1488), .A1(N100), .A2(N582), .A3(N1113) );
  AND3_X1 AND3_252( .ZN(N1489), .A1(N124), .A2(N1102), .A3(N594) );
  AND3_X1 AND3_253( .ZN(N1490), .A1(N135), .A2(N1102), .A3(N1113) );
  AND3_X1 AND3_254( .ZN(N1491), .A1(N99), .A2(N582), .A3(N1113) );
  AND3_X1 AND3_255( .ZN(N1492), .A1(N123), .A2(N1102), .A3(N594) );
  AND2_X1 AND2_256( .ZN(N1493), .A1(N1102), .A2(N1113) );
  AND2_X1 AND2_257( .ZN(N1494), .A1(N582), .A2(N1113) );
  AND2_X1 AND2_258( .ZN(N1495), .A1(N1102), .A2(N594) );
  INV_X1 NOT1_259( .ZN(N1496), .A(N1129) );
  INV_X1 NOT1_260( .ZN(N1499), .A(N1133) );
  NAND2_X1 NAND2_261( .ZN(N1502), .A1(N1351), .A2(N1141) );
  NAND2_X1 NAND2_262( .ZN(N1506), .A1(N1352), .A2(N1353) );
  NAND2_X1 NAND2_263( .ZN(N1510), .A1(N1354), .A2(N1355) );
  BUF_X2 BUFF1_264( .Z(N1513), .A(N1137) );
  BUF_X2 BUFF1_265( .Z(N1516), .A(N1137) );
  INV_X1 NOT1_266( .ZN(N1519), .A(N1219) );
  INV_X1 NOT1_267( .ZN(N1520), .A(N1222) );
  INV_X1 NOT1_268( .ZN(N1521), .A(N1225) );
  INV_X1 NOT1_269( .ZN(N1522), .A(N1228) );
  INV_X1 NOT1_270( .ZN(N1523), .A(N1231) );
  INV_X1 NOT1_271( .ZN(N1524), .A(N1234) );
  INV_X1 NOT1_272( .ZN(N1525), .A(N1237) );
  INV_X1 NOT1_273( .ZN(N1526), .A(N1240) );
  INV_X1 NOT1_274( .ZN(N1527), .A(N1243) );
  INV_X1 NOT1_275( .ZN(N1528), .A(N1246) );
  AND3_X1 AND3_276( .ZN(N1529), .A1(N142), .A2(N1146), .A3(N1157) );
  AND3_X1 AND3_277( .ZN(N1530), .A1(N106), .A2(N613), .A3(N1157) );
  AND3_X1 AND3_278( .ZN(N1531), .A1(N130), .A2(N1146), .A3(N625) );
  AND3_X1 AND3_279( .ZN(N1532), .A1(N131), .A2(N1146), .A3(N1157) );
  AND3_X1 AND3_280( .ZN(N1533), .A1(N95), .A2(N613), .A3(N1157) );
  AND3_X1 AND3_281( .ZN(N1534), .A1(N119), .A2(N1146), .A3(N625) );
  AND3_X1 AND3_282( .ZN(N1535), .A1(N141), .A2(N1146), .A3(N1157) );
  AND3_X1 AND3_283( .ZN(N1536), .A1(N105), .A2(N613), .A3(N1157) );
  AND3_X1 AND3_284( .ZN(N1537), .A1(N129), .A2(N1146), .A3(N625) );
  AND3_X1 AND3_285( .ZN(N1538), .A1(N140), .A2(N1146), .A3(N1157) );
  AND3_X1 AND3_286( .ZN(N1539), .A1(N104), .A2(N613), .A3(N1157) );
  AND3_X1 AND3_287( .ZN(N1540), .A1(N128), .A2(N1146), .A3(N625) );
  AND3_X1 AND3_288( .ZN(N1541), .A1(N139), .A2(N1146), .A3(N1157) );
  AND3_X1 AND3_289( .ZN(N1542), .A1(N103), .A2(N613), .A3(N1157) );
  AND3_X1 AND3_290( .ZN(N1543), .A1(N127), .A2(N1146), .A3(N625) );
  AND2_X1 AND2_291( .ZN(N1544), .A1(N19), .A2(N1173) );
  AND2_X1 AND2_292( .ZN(N1545), .A1(N4), .A2(N1173) );
  AND2_X1 AND2_293( .ZN(N1546), .A1(N20), .A2(N1173) );
  AND2_X1 AND2_294( .ZN(N1547), .A1(N5), .A2(N1173) );
  AND2_X1 AND2_295( .ZN(N1548), .A1(N21), .A2(N1178) );
  AND2_X1 AND2_296( .ZN(N1549), .A1(N22), .A2(N1178) );
  AND2_X1 AND2_297( .ZN(N1550), .A1(N23), .A2(N1178) );
  AND2_X1 AND2_298( .ZN(N1551), .A1(N6), .A2(N1178) );
  AND2_X1 AND2_299( .ZN(N1552), .A1(N24), .A2(N1178) );
  NAND2_X1 NAND2_300( .ZN(N1553), .A1(N1395), .A2(N1185) );
  NAND2_X1 NAND2_301( .ZN(N1557), .A1(N1396), .A2(N1397) );
  NAND2_X1 NAND2_302( .ZN(N1561), .A1(N1398), .A2(N1399) );
  AND2_X1 AND2_303( .ZN(N1564), .A1(N25), .A2(N1200) );
  AND2_X1 AND2_304( .ZN(N1565), .A1(N32), .A2(N1200) );
  AND2_X1 AND2_305( .ZN(N1566), .A1(N26), .A2(N1200) );
  AND2_X1 AND2_306( .ZN(N1567), .A1(N33), .A2(N1200) );
  AND2_X1 AND2_307( .ZN(N1568), .A1(N27), .A2(N1205) );
  AND2_X1 AND2_308( .ZN(N1569), .A1(N34), .A2(N1205) );
  AND2_X1 AND2_309( .ZN(N1570), .A1(N35), .A2(N1205) );
  AND2_X1 AND2_310( .ZN(N1571), .A1(N28), .A2(N1205) );
  INV_X2 NOT1_311( .ZN(N1572), .A(N1251) );
  INV_X2 NOT1_312( .ZN(N1573), .A(N1254) );
  INV_X2 NOT1_313( .ZN(N1574), .A(N1257) );
  INV_X1 NOT1_314( .ZN(N1575), .A(N1260) );
  INV_X1 NOT1_315( .ZN(N1576), .A(N1263) );
  INV_X1 NOT1_316( .ZN(N1577), .A(N1266) );
  NAND2_X1 NAND2_317( .ZN(N1578), .A1(N1422), .A2(N1423) );
  INV_X1 NOT1_318( .ZN(N1581), .A(N1216) );
  NAND2_X1 NAND2_319( .ZN(N1582), .A1(N1426), .A2(N1427) );
  NAND2_X1 NAND2_320( .ZN(N1585), .A1(N1424), .A2(N1425) );
  NAND2_X1 NAND2_321( .ZN(N1588), .A1(N1440), .A2(N1441) );
  AND2_X1 AND2_322( .ZN(N1591), .A1(N1449), .A2(N1450) );
  OR4_X1 OR4_323( .ZN(N1596), .A1(N1451), .A2(N1452), .A3(N1453), .A4(N1064) );
  OR4_X1 OR4_324( .ZN(N1600), .A1(N1454), .A2(N1455), .A3(N1456), .A4(N1065) );
  OR4_X1 OR4_325( .ZN(N1606), .A1(N1457), .A2(N1458), .A3(N1459), .A4(N1066) );
  OR4_X1 OR4_326( .ZN(N1612), .A1(N1460), .A2(N1461), .A3(N1462), .A4(N1067) );
  OR4_X1 OR4_327( .ZN(N1615), .A1(N1463), .A2(N1464), .A3(N1465), .A4(N1068) );
  OR4_X1 OR4_328( .ZN(N1619), .A1(N1466), .A2(N1467), .A3(N1468), .A4(N1097) );
  OR4_X1 OR4_329( .ZN(N1624), .A1(N1469), .A2(N1470), .A3(N1471), .A4(N1098) );
  OR4_X1 OR4_330( .ZN(N1628), .A1(N1472), .A2(N1473), .A3(N1474), .A4(N1099) );
  OR4_X1 OR4_331( .ZN(N1631), .A1(N1475), .A2(N1476), .A3(N1477), .A4(N1100) );
  OR4_X1 OR4_332( .ZN(N1634), .A1(N1478), .A2(N1479), .A3(N1480), .A4(N1101) );
  OR4_X1 OR4_333( .ZN(N1637), .A1(N1481), .A2(N1482), .A3(N1483), .A4(N1124) );
  OR4_X1 OR4_334( .ZN(N1642), .A1(N1484), .A2(N1485), .A3(N1486), .A4(N1125) );
  OR4_X1 OR4_335( .ZN(N1647), .A1(N1487), .A2(N1488), .A3(N1489), .A4(N1126) );
  OR4_X1 OR4_336( .ZN(N1651), .A1(N1490), .A2(N1491), .A3(N1492), .A4(N1127) );
  OR4_X1 OR4_337( .ZN(N1656), .A1(N1493), .A2(N1494), .A3(N1495), .A4(N1128) );
  OR4_X1 OR4_338( .ZN(N1676), .A1(N1532), .A2(N1533), .A3(N1534), .A4(N1169) );
  OR4_X1 OR4_339( .ZN(N1681), .A1(N1535), .A2(N1536), .A3(N1537), .A4(N1170) );
  OR4_X1 OR4_340( .ZN(N1686), .A1(N1538), .A2(N1539), .A3(N1540), .A4(N1171) );
  OR4_X1 OR4_341( .ZN(N1690), .A1(N1541), .A2(N1542), .A3(N1543), .A4(N1172) );
  OR4_X1 OR4_342( .ZN(N1708), .A1(N1529), .A2(N1530), .A3(N1531), .A4(N1168) );
  BUF_X1 BUFF1_343( .Z(N1726), .A(N1591) );
  INV_X1 NOT1_344( .ZN(N1770), .A(N1502) );
  INV_X1 NOT1_345( .ZN(N1773), .A(N1506) );
  INV_X1 NOT1_346( .ZN(N1776), .A(N1513) );
  INV_X1 NOT1_347( .ZN(N1777), .A(N1516) );
  BUF_X1 BUFF1_348( .Z(N1778), .A(N1510) );
  BUF_X1 BUFF1_349( .Z(N1781), .A(N1510) );
  AND3_X1 AND3_350( .ZN(N1784), .A1(N1133), .A2(N1129), .A3(N1513) );
  AND3_X1 AND3_351( .ZN(N1785), .A1(N1499), .A2(N1496), .A3(N1516) );
  INV_X1 NOT1_352( .ZN(N1795), .A(N1553) );
  INV_X1 NOT1_353( .ZN(N1798), .A(N1557) );
  BUF_X1 BUFF1_354( .Z(N1801), .A(N1561) );
  BUF_X1 BUFF1_355( .Z(N1804), .A(N1561) );
  INV_X1 NOT1_356( .ZN(N1807), .A(N1588) );
  INV_X1 NOT1_357( .ZN(N1808), .A(N1578) );
  NAND2_X2 NAND2_358( .ZN(N1809), .A1(N1578), .A2(N1581) );
  INV_X1 NOT1_359( .ZN(N1810), .A(N1582) );
  INV_X1 NOT1_360( .ZN(N1811), .A(N1585) );
  AND2_X2 AND2_361( .ZN(N1813), .A1(N1596), .A2(N241) );
  AND2_X2 AND2_362( .ZN(N1814), .A1(N1606), .A2(N241) );
  AND2_X1 AND2_363( .ZN(N1815), .A1(N1600), .A2(N241) );
  INV_X1 NOT1_364( .ZN(N1816), .A(N1642) );
  INV_X1 NOT1_365( .ZN(N1817), .A(N1647) );
  INV_X1 NOT1_366( .ZN(N1818), .A(N1637) );
  INV_X1 NOT1_367( .ZN(N1819), .A(N1624) );
  INV_X1 NOT1_368( .ZN(N1820), .A(N1619) );
  INV_X1 NOT1_369( .ZN(N1821), .A(N1615) );
  AND4_X1 AND4_370( .ZN(N1822), .A1(N496), .A2(N224), .A3(N36), .A4(N1591) );
  AND4_X1 AND4_371( .ZN(N1823), .A1(N496), .A2(N224), .A3(N1591), .A4(N486) );
  BUF_X1 BUFF1_372( .Z(N1824), .A(N1596) );
  INV_X1 NOT1_373( .ZN(N1827), .A(N1606) );
  AND2_X1 AND2_374( .ZN(N1830), .A1(N1600), .A2(N537) );
  AND2_X1 AND2_375( .ZN(N1831), .A1(N1606), .A2(N537) );
  AND2_X1 AND2_376( .ZN(N1832), .A1(N1619), .A2(N246) );
  INV_X1 NOT1_377( .ZN(N1833), .A(N1596) );
  INV_X1 NOT1_378( .ZN(N1836), .A(N1600) );
  INV_X1 NOT1_379( .ZN(N1841), .A(N1606) );
  BUF_X1 BUFF1_380( .Z(N1848), .A(N1612) );
  BUF_X1 BUFF1_381( .Z(N1852), .A(N1615) );
  BUF_X1 BUFF1_382( .Z(N1856), .A(N1619) );
  BUF_X1 BUFF1_383( .Z(N1863), .A(N1624) );
  BUF_X1 BUFF1_384( .Z(N1870), .A(N1628) );
  BUF_X1 BUFF1_385( .Z(N1875), .A(N1631) );
  BUF_X1 BUFF1_386( .Z(N1880), .A(N1634) );
  NAND2_X1 NAND2_387( .ZN(N1885), .A1(N727), .A2(N1651) );
  NAND2_X1 NAND2_388( .ZN(N1888), .A1(N730), .A2(N1656) );
  BUF_X1 BUFF1_389( .Z(N1891), .A(N1686) );
  AND2_X1 AND2_390( .ZN(N1894), .A1(N1637), .A2(N425) );
  INV_X1 NOT1_391( .ZN(N1897), .A(N1642) );
  AND3_X1 AND3_392( .ZN(N1908), .A1(N1496), .A2(N1133), .A3(N1776) );
  AND3_X1 AND3_393( .ZN(N1909), .A1(N1129), .A2(N1499), .A3(N1777) );
  AND2_X1 AND2_394( .ZN(N1910), .A1(N1600), .A2(N637) );
  AND2_X1 AND2_395( .ZN(N1911), .A1(N1606), .A2(N637) );
  AND2_X1 AND2_396( .ZN(N1912), .A1(N1612), .A2(N637) );
  AND2_X1 AND2_397( .ZN(N1913), .A1(N1615), .A2(N637) );
  AND2_X1 AND2_398( .ZN(N1914), .A1(N1619), .A2(N643) );
  AND2_X1 AND2_399( .ZN(N1915), .A1(N1624), .A2(N643) );
  AND2_X1 AND2_400( .ZN(N1916), .A1(N1628), .A2(N643) );
  AND2_X1 AND2_401( .ZN(N1917), .A1(N1631), .A2(N643) );
  AND2_X1 AND2_402( .ZN(N1918), .A1(N1634), .A2(N643) );
  INV_X1 NOT1_403( .ZN(N1919), .A(N1708) );
  AND2_X1 AND2_404( .ZN(N1928), .A1(N1676), .A2(N693) );
  AND2_X1 AND2_405( .ZN(N1929), .A1(N1681), .A2(N693) );
  AND2_X1 AND2_406( .ZN(N1930), .A1(N1686), .A2(N693) );
  AND2_X1 AND2_407( .ZN(N1931), .A1(N1690), .A2(N693) );
  AND2_X1 AND2_408( .ZN(N1932), .A1(N1637), .A2(N699) );
  AND2_X1 AND2_409( .ZN(N1933), .A1(N1642), .A2(N699) );
  AND2_X1 AND2_410( .ZN(N1934), .A1(N1647), .A2(N699) );
  AND2_X1 AND2_411( .ZN(N1935), .A1(N1651), .A2(N699) );
  BUF_X1 BUFF1_412( .Z(N1936), .A(N1600) );
  NAND2_X1 NAND2_413( .ZN(N1939), .A1(N1216), .A2(N1808) );
  NAND2_X1 NAND2_414( .ZN(N1940), .A1(N1585), .A2(N1810) );
  NAND2_X1 NAND2_415( .ZN(N1941), .A1(N1582), .A2(N1811) );
  BUF_X1 BUFF1_416( .Z(N1942), .A(N1676) );
  BUF_X1 BUFF1_417( .Z(N1945), .A(N1686) );
  BUF_X1 BUFF1_418( .Z(N1948), .A(N1681) );
  BUF_X1 BUFF1_419( .Z(N1951), .A(N1637) );
  BUF_X1 BUFF1_420( .Z(N1954), .A(N1690) );
  BUF_X1 BUFF1_421( .Z(N1957), .A(N1647) );
  BUF_X1 BUFF1_422( .Z(N1960), .A(N1642) );
  BUF_X1 BUFF1_423( .Z(N1963), .A(N1656) );
  BUF_X1 BUFF1_424( .Z(N1966), .A(N1651) );
  OR2_X1 OR2_425( .ZN(N1969), .A1(N533), .A2(N1815) );
  INV_X1 NOT1_426( .ZN(N1970), .A(N1822) );
  INV_X1 NOT1_427( .ZN(N1971), .A(N1823) );
  BUF_X1 BUFF1_428( .Z(N2010), .A(N1848) );
  BUF_X1 BUFF1_429( .Z(N2012), .A(N1852) );
  BUF_X1 BUFF1_430( .Z(N2014), .A(N1856) );
  BUF_X1 BUFF1_431( .Z(N2016), .A(N1863) );
  BUF_X1 BUFF1_432( .Z(N2018), .A(N1870) );
  BUF_X1 BUFF1_433( .Z(N2020), .A(N1875) );
  BUF_X1 BUFF1_434( .Z(N2022), .A(N1880) );
  INV_X1 NOT1_435( .ZN(N2028), .A(N1778) );
  INV_X1 NOT1_436( .ZN(N2029), .A(N1781) );
  NOR2_X1 NOR2_437( .ZN(N2030), .A1(N1908), .A2(N1784) );
  NOR2_X1 NOR2_438( .ZN(N2031), .A1(N1909), .A2(N1785) );
  AND3_X1 AND3_439( .ZN(N2032), .A1(N1506), .A2(N1502), .A3(N1778) );
  AND3_X1 AND3_440( .ZN(N2033), .A1(N1773), .A2(N1770), .A3(N1781) );
  OR2_X1 OR2_441( .ZN(N2034), .A1(N1571), .A2(N1935) );
  INV_X1 NOT1_442( .ZN(N2040), .A(N1801) );
  INV_X1 NOT1_443( .ZN(N2041), .A(N1804) );
  AND3_X1 AND3_444( .ZN(N2042), .A1(N1557), .A2(N1553), .A3(N1801) );
  AND3_X1 AND3_445( .ZN(N2043), .A1(N1798), .A2(N1795), .A3(N1804) );
  NAND2_X1 NAND2_446( .ZN(N2046), .A1(N1939), .A2(N1809) );
  NAND2_X1 NAND2_447( .ZN(N2049), .A1(N1940), .A2(N1941) );
  OR2_X1 OR2_448( .ZN(N2052), .A1(N1544), .A2(N1910) );
  OR2_X1 OR2_449( .ZN(N2055), .A1(N1545), .A2(N1911) );
  OR2_X1 OR2_450( .ZN(N2058), .A1(N1546), .A2(N1912) );
  OR2_X1 OR2_451( .ZN(N2061), .A1(N1547), .A2(N1913) );
  OR2_X1 OR2_452( .ZN(N2064), .A1(N1548), .A2(N1914) );
  OR2_X1 OR2_453( .ZN(N2067), .A1(N1549), .A2(N1915) );
  OR2_X1 OR2_454( .ZN(N2070), .A1(N1550), .A2(N1916) );
  OR2_X1 OR2_455( .ZN(N2073), .A1(N1551), .A2(N1917) );
  OR2_X1 OR2_456( .ZN(N2076), .A1(N1552), .A2(N1918) );
  OR2_X1 OR2_457( .ZN(N2079), .A1(N1564), .A2(N1928) );
  OR2_X1 OR2_458( .ZN(N2095), .A1(N1565), .A2(N1929) );
  OR2_X1 OR2_459( .ZN(N2098), .A1(N1566), .A2(N1930) );
  OR2_X1 OR2_460( .ZN(N2101), .A1(N1567), .A2(N1931) );
  OR2_X1 OR2_461( .ZN(N2104), .A1(N1568), .A2(N1932) );
  OR2_X1 OR2_462( .ZN(N2107), .A1(N1569), .A2(N1933) );
  OR2_X1 OR2_463( .ZN(N2110), .A1(N1570), .A2(N1934) );
  AND3_X1 AND3_464( .ZN(N2113), .A1(N1897), .A2(N1894), .A3(N40) );
  INV_X2 NOT1_465( .ZN(N2119), .A(N1894) );
  NAND2_X1 NAND2_466( .ZN(N2120), .A1(N408), .A2(N1827) );
  AND2_X1 AND2_467( .ZN(N2125), .A1(N1824), .A2(N537) );
  AND2_X1 AND2_468( .ZN(N2126), .A1(N1852), .A2(N246) );
  AND2_X1 AND2_469( .ZN(N2127), .A1(N1848), .A2(N537) );
  INV_X1 NOT1_470( .ZN(N2128), .A(N1848) );
  INV_X1 NOT1_471( .ZN(N2135), .A(N1852) );
  INV_X1 NOT1_472( .ZN(N2141), .A(N1863) );
  INV_X1 NOT1_473( .ZN(N2144), .A(N1870) );
  INV_X1 NOT1_474( .ZN(N2147), .A(N1875) );
  INV_X1 NOT1_475( .ZN(N2150), .A(N1880) );
  AND2_X1 AND2_476( .ZN(N2153), .A1(N727), .A2(N1885) );
  AND2_X1 AND2_477( .ZN(N2154), .A1(N1885), .A2(N1651) );
  AND2_X1 AND2_478( .ZN(N2155), .A1(N730), .A2(N1888) );
  AND2_X1 AND2_479( .ZN(N2156), .A1(N1888), .A2(N1656) );
  AND3_X1 AND3_480( .ZN(N2157), .A1(N1770), .A2(N1506), .A3(N2028) );
  AND3_X1 AND3_481( .ZN(N2158), .A1(N1502), .A2(N1773), .A3(N2029) );
  INV_X1 NOT1_482( .ZN(N2171), .A(N1942) );
  NAND2_X1 NAND2_483( .ZN(N2172), .A1(N1942), .A2(N1919) );
  INV_X1 NOT1_484( .ZN(N2173), .A(N1945) );
  INV_X1 NOT1_485( .ZN(N2174), .A(N1948) );
  INV_X1 NOT1_486( .ZN(N2175), .A(N1951) );
  INV_X1 NOT1_487( .ZN(N2176), .A(N1954) );
  AND3_X1 AND3_488( .ZN(N2177), .A1(N1795), .A2(N1557), .A3(N2040) );
  AND3_X1 AND3_489( .ZN(N2178), .A1(N1553), .A2(N1798), .A3(N2041) );
  BUF_X2 BUFF1_490( .Z(N2185), .A(N1836) );
  BUF_X2 BUFF1_491( .Z(N2188), .A(N1833) );
  BUF_X1 BUFF1_492( .Z(N2191), .A(N1841) );
  INV_X2 NOT1_493( .ZN(N2194), .A(N1856) );
  INV_X1 NOT1_494( .ZN(N2197), .A(N1827) );
  INV_X1 NOT1_495( .ZN(N2200), .A(N1936) );
  BUF_X1 BUFF1_496( .Z(N2201), .A(N1836) );
  BUF_X1 BUFF1_497( .Z(N2204), .A(N1833) );
  BUF_X1 BUFF1_498( .Z(N2207), .A(N1841) );
  BUF_X1 BUFF1_499( .Z(N2210), .A(N1824) );
  BUF_X1 BUFF1_500( .Z(N2213), .A(N1841) );
  BUF_X1 BUFF1_501( .Z(N2216), .A(N1841) );
  NAND2_X1 NAND2_502( .ZN(N2219), .A1(N2031), .A2(N2030) );
  INV_X1 NOT1_503( .ZN(N2234), .A(N1957) );
  INV_X1 NOT1_504( .ZN(N2235), .A(N1960) );
  INV_X1 NOT1_505( .ZN(N2236), .A(N1963) );
  INV_X1 NOT1_506( .ZN(N2237), .A(N1966) );
  AND3_X1 AND3_507( .ZN(N2250), .A1(N40), .A2(N1897), .A3(N2119) );
  OR2_X1 OR2_508( .ZN(N2266), .A1(N1831), .A2(N2126) );
  OR2_X1 OR2_509( .ZN(N2269), .A1(N2127), .A2(N1832) );
  OR2_X1 OR2_510( .ZN(N2291), .A1(N2153), .A2(N2154) );
  OR2_X1 OR2_511( .ZN(N2294), .A1(N2155), .A2(N2156) );
  NOR2_X1 NOR2_512( .ZN(N2297), .A1(N2157), .A2(N2032) );
  NOR2_X1 NOR2_513( .ZN(N2298), .A1(N2158), .A2(N2033) );
  INV_X1 NOT1_514( .ZN(N2300), .A(N2046) );
  INV_X1 NOT1_515( .ZN(N2301), .A(N2049) );
  NAND2_X1 NAND2_516( .ZN(N2302), .A1(N2052), .A2(N1519) );
  INV_X1 NOT1_517( .ZN(N2303), .A(N2052) );
  NAND2_X1 NAND2_518( .ZN(N2304), .A1(N2055), .A2(N1520) );
  INV_X1 NOT1_519( .ZN(N2305), .A(N2055) );
  NAND2_X1 NAND2_520( .ZN(N2306), .A1(N2058), .A2(N1521) );
  INV_X1 NOT1_521( .ZN(N2307), .A(N2058) );
  NAND2_X1 NAND2_522( .ZN(N2308), .A1(N2061), .A2(N1522) );
  INV_X1 NOT1_523( .ZN(N2309), .A(N2061) );
  NAND2_X1 NAND2_524( .ZN(N2310), .A1(N2064), .A2(N1523) );
  INV_X1 NOT1_525( .ZN(N2311), .A(N2064) );
  NAND2_X1 NAND2_526( .ZN(N2312), .A1(N2067), .A2(N1524) );
  INV_X1 NOT1_527( .ZN(N2313), .A(N2067) );
  NAND2_X1 NAND2_528( .ZN(N2314), .A1(N2070), .A2(N1525) );
  INV_X1 NOT1_529( .ZN(N2315), .A(N2070) );
  NAND2_X1 NAND2_530( .ZN(N2316), .A1(N2073), .A2(N1526) );
  INV_X1 NOT1_531( .ZN(N2317), .A(N2073) );
  NAND2_X1 NAND2_532( .ZN(N2318), .A1(N2076), .A2(N1527) );
  INV_X1 NOT1_533( .ZN(N2319), .A(N2076) );
  NAND2_X1 NAND2_534( .ZN(N2320), .A1(N2079), .A2(N1528) );
  INV_X1 NOT1_535( .ZN(N2321), .A(N2079) );
  NAND2_X1 NAND2_536( .ZN(N2322), .A1(N1708), .A2(N2171) );
  NAND2_X1 NAND2_537( .ZN(N2323), .A1(N1948), .A2(N2173) );
  NAND2_X1 NAND2_538( .ZN(N2324), .A1(N1945), .A2(N2174) );
  NAND2_X1 NAND2_539( .ZN(N2325), .A1(N1954), .A2(N2175) );
  NAND2_X1 NAND2_540( .ZN(N2326), .A1(N1951), .A2(N2176) );
  NOR2_X1 NOR2_541( .ZN(N2327), .A1(N2177), .A2(N2042) );
  NOR2_X1 NOR2_542( .ZN(N2328), .A1(N2178), .A2(N2043) );
  NAND2_X1 NAND2_543( .ZN(N2329), .A1(N2095), .A2(N1572) );
  INV_X4 NOT1_544( .ZN(N2330), .A(N2095) );
  NAND2_X1 NAND2_545( .ZN(N2331), .A1(N2098), .A2(N1573) );
  INV_X1 NOT1_546( .ZN(N2332), .A(N2098) );
  NAND2_X1 NAND2_547( .ZN(N2333), .A1(N2101), .A2(N1574) );
  INV_X1 NOT1_548( .ZN(N2334), .A(N2101) );
  NAND2_X1 NAND2_549( .ZN(N2335), .A1(N2104), .A2(N1575) );
  INV_X1 NOT1_550( .ZN(N2336), .A(N2104) );
  NAND2_X1 NAND2_551( .ZN(N2337), .A1(N2107), .A2(N1576) );
  INV_X1 NOT1_552( .ZN(N2338), .A(N2107) );
  NAND2_X2 NAND2_553( .ZN(N2339), .A1(N2110), .A2(N1577) );
  INV_X1 NOT1_554( .ZN(N2340), .A(N2110) );
  NAND2_X1 NAND2_555( .ZN(N2354), .A1(N1960), .A2(N2234) );
  NAND2_X1 NAND2_556( .ZN(N2355), .A1(N1957), .A2(N2235) );
  NAND2_X1 NAND2_557( .ZN(N2356), .A1(N1966), .A2(N2236) );
  NAND2_X1 NAND2_558( .ZN(N2357), .A1(N1963), .A2(N2237) );
  AND2_X2 AND2_559( .ZN(N2358), .A1(N2120), .A2(N533) );
  INV_X1 NOT1_560( .ZN(N2359), .A(N2113) );
  INV_X1 NOT1_561( .ZN(N2364), .A(N2185) );
  INV_X1 NOT1_562( .ZN(N2365), .A(N2188) );
  INV_X1 NOT1_563( .ZN(N2366), .A(N2191) );
  INV_X1 NOT1_564( .ZN(N2367), .A(N2194) );
  BUF_X1 BUFF1_565( .Z(N2368), .A(N2120) );
  INV_X1 NOT1_566( .ZN(N2372), .A(N2201) );
  INV_X1 NOT1_567( .ZN(N2373), .A(N2204) );
  INV_X1 NOT1_568( .ZN(N2374), .A(N2207) );
  INV_X1 NOT1_569( .ZN(N2375), .A(N2210) );
  INV_X1 NOT1_570( .ZN(N2376), .A(N2213) );
  INV_X1 NOT1_571( .ZN(N2377), .A(N2113) );
  BUF_X1 BUFF1_572( .Z(N2382), .A(N2113) );
  AND2_X1 AND2_573( .ZN(N2386), .A1(N2120), .A2(N246) );
  BUF_X1 BUFF1_574( .Z(N2387), .A(N2266) );
  BUF_X1 BUFF1_575( .Z(N2388), .A(N2266) );
  BUF_X1 BUFF1_576( .Z(N2389), .A(N2269) );
  BUF_X1 BUFF1_577( .Z(N2390), .A(N2269) );
  BUF_X1 BUFF1_578( .Z(N2391), .A(N2113) );
  INV_X1 NOT1_579( .ZN(N2395), .A(N2113) );
  NAND2_X1 NAND2_580( .ZN(N2400), .A1(N2219), .A2(N2300) );
  INV_X1 NOT1_581( .ZN(N2403), .A(N2216) );
  INV_X1 NOT1_582( .ZN(N2406), .A(N2219) );
  NAND2_X1 NAND2_583( .ZN(N2407), .A1(N1219), .A2(N2303) );
  NAND2_X1 NAND2_584( .ZN(N2408), .A1(N1222), .A2(N2305) );
  NAND2_X1 NAND2_585( .ZN(N2409), .A1(N1225), .A2(N2307) );
  NAND2_X1 NAND2_586( .ZN(N2410), .A1(N1228), .A2(N2309) );
  NAND2_X1 NAND2_587( .ZN(N2411), .A1(N1231), .A2(N2311) );
  NAND2_X1 NAND2_588( .ZN(N2412), .A1(N1234), .A2(N2313) );
  NAND2_X1 NAND2_589( .ZN(N2413), .A1(N1237), .A2(N2315) );
  NAND2_X1 NAND2_590( .ZN(N2414), .A1(N1240), .A2(N2317) );
  NAND2_X1 NAND2_591( .ZN(N2415), .A1(N1243), .A2(N2319) );
  NAND2_X1 NAND2_592( .ZN(N2416), .A1(N1246), .A2(N2321) );
  NAND2_X1 NAND2_593( .ZN(N2417), .A1(N2322), .A2(N2172) );
  NAND2_X1 NAND2_594( .ZN(N2421), .A1(N2323), .A2(N2324) );
  NAND2_X1 NAND2_595( .ZN(N2425), .A1(N2325), .A2(N2326) );
  NAND2_X1 NAND2_596( .ZN(N2428), .A1(N1251), .A2(N2330) );
  NAND2_X1 NAND2_597( .ZN(N2429), .A1(N1254), .A2(N2332) );
  NAND2_X1 NAND2_598( .ZN(N2430), .A1(N1257), .A2(N2334) );
  NAND2_X1 NAND2_599( .ZN(N2431), .A1(N1260), .A2(N2336) );
  NAND2_X1 NAND2_600( .ZN(N2432), .A1(N1263), .A2(N2338) );
  NAND2_X1 NAND2_601( .ZN(N2433), .A1(N1266), .A2(N2340) );
  BUF_X4 BUFF1_602( .Z(N2434), .A(N2128) );
  BUF_X4 BUFF1_603( .Z(N2437), .A(N2135) );
  BUF_X1 BUFF1_604( .Z(N2440), .A(N2144) );
  BUF_X1 BUFF1_605( .Z(N2443), .A(N2141) );
  BUF_X1 BUFF1_606( .Z(N2446), .A(N2150) );
  BUF_X1 BUFF1_607( .Z(N2449), .A(N2147) );
  INV_X1 NOT1_608( .ZN(N2452), .A(N2197) );
  NAND2_X1 NAND2_609( .ZN(N2453), .A1(N2197), .A2(N2200) );
  BUF_X1 BUFF1_610( .Z(N2454), .A(N2128) );
  BUF_X1 BUFF1_611( .Z(N2457), .A(N2144) );
  BUF_X1 BUFF1_612( .Z(N2460), .A(N2141) );
  BUF_X1 BUFF1_613( .Z(N2463), .A(N2150) );
  BUF_X1 BUFF1_614( .Z(N2466), .A(N2147) );
  INV_X1 NOT1_615( .ZN(N2469), .A(N2120) );
  BUF_X1 BUFF1_616( .Z(N2472), .A(N2128) );
  BUF_X1 BUFF1_617( .Z(N2475), .A(N2135) );
  BUF_X1 BUFF1_618( .Z(N2478), .A(N2128) );
  BUF_X1 BUFF1_619( .Z(N2481), .A(N2135) );
  NAND2_X1 NAND2_620( .ZN(N2484), .A1(N2298), .A2(N2297) );
  NAND2_X1 NAND2_621( .ZN(N2487), .A1(N2356), .A2(N2357) );
  NAND2_X1 NAND2_622( .ZN(N2490), .A1(N2354), .A2(N2355) );
  NAND2_X1 NAND2_623( .ZN(N2493), .A1(N2328), .A2(N2327) );
  OR2_X1 OR2_624( .ZN(N2496), .A1(N2358), .A2(N1814) );
  NAND2_X1 NAND2_625( .ZN(N2503), .A1(N2188), .A2(N2364) );
  NAND2_X1 NAND2_626( .ZN(N2504), .A1(N2185), .A2(N2365) );
  NAND2_X1 NAND2_627( .ZN(N2510), .A1(N2204), .A2(N2372) );
  NAND2_X1 NAND2_628( .ZN(N2511), .A1(N2201), .A2(N2373) );
  OR2_X1 OR2_629( .ZN(N2521), .A1(N1830), .A2(N2386) );
  NAND2_X1 NAND2_630( .ZN(N2528), .A1(N2046), .A2(N2406) );
  INV_X1 NOT1_631( .ZN(N2531), .A(N2291) );
  INV_X1 NOT1_632( .ZN(N2534), .A(N2294) );
  BUF_X1 BUFF1_633( .Z(N2537), .A(N2250) );
  BUF_X1 BUFF1_634( .Z(N2540), .A(N2250) );
  NAND2_X1 NAND2_635( .ZN(N2544), .A1(N2302), .A2(N2407) );
  NAND2_X1 NAND2_636( .ZN(N2545), .A1(N2304), .A2(N2408) );
  NAND2_X1 NAND2_637( .ZN(N2546), .A1(N2306), .A2(N2409) );
  NAND2_X1 NAND2_638( .ZN(N2547), .A1(N2308), .A2(N2410) );
  NAND2_X1 NAND2_639( .ZN(N2548), .A1(N2310), .A2(N2411) );
  NAND2_X1 NAND2_640( .ZN(N2549), .A1(N2312), .A2(N2412) );
  NAND2_X1 NAND2_641( .ZN(N2550), .A1(N2314), .A2(N2413) );
  NAND2_X1 NAND2_642( .ZN(N2551), .A1(N2316), .A2(N2414) );
  NAND2_X1 NAND2_643( .ZN(N2552), .A1(N2318), .A2(N2415) );
  NAND2_X1 NAND2_644( .ZN(N2553), .A1(N2320), .A2(N2416) );
  NAND2_X1 NAND2_645( .ZN(N2563), .A1(N2329), .A2(N2428) );
  NAND2_X1 NAND2_646( .ZN(N2564), .A1(N2331), .A2(N2429) );
  NAND2_X1 NAND2_647( .ZN(N2565), .A1(N2333), .A2(N2430) );
  NAND2_X1 NAND2_648( .ZN(N2566), .A1(N2335), .A2(N2431) );
  NAND2_X1 NAND2_649( .ZN(N2567), .A1(N2337), .A2(N2432) );
  NAND2_X1 NAND2_650( .ZN(N2568), .A1(N2339), .A2(N2433) );
  NAND2_X1 NAND2_651( .ZN(N2579), .A1(N1936), .A2(N2452) );
  BUF_X1 BUFF1_652( .Z(N2603), .A(N2359) );
  AND2_X2 AND2_653( .ZN(N2607), .A1(N1880), .A2(N2377) );
  AND2_X2 AND2_654( .ZN(N2608), .A1(N1676), .A2(N2377) );
  AND2_X1 AND2_655( .ZN(N2609), .A1(N1681), .A2(N2377) );
  AND2_X1 AND2_656( .ZN(N2610), .A1(N1891), .A2(N2377) );
  AND2_X1 AND2_657( .ZN(N2611), .A1(N1856), .A2(N2382) );
  AND2_X1 AND2_658( .ZN(N2612), .A1(N1863), .A2(N2382) );
  NAND2_X1 NAND2_659( .ZN(N2613), .A1(N2503), .A2(N2504) );
  INV_X4 NOT1_660( .ZN(N2617), .A(N2434) );
  NAND2_X1 NAND2_661( .ZN(N2618), .A1(N2434), .A2(N2366) );
  NAND2_X1 NAND2_662( .ZN(N2619), .A1(N2437), .A2(N2367) );
  INV_X1 NOT1_663( .ZN(N2620), .A(N2437) );
  INV_X1 NOT1_664( .ZN(N2621), .A(N2368) );
  NAND2_X1 NAND2_665( .ZN(N2624), .A1(N2510), .A2(N2511) );
  INV_X1 NOT1_666( .ZN(N2628), .A(N2454) );
  NAND2_X1 NAND2_667( .ZN(N2629), .A1(N2454), .A2(N2374) );
  INV_X1 NOT1_668( .ZN(N2630), .A(N2472) );
  AND2_X1 AND2_669( .ZN(N2631), .A1(N1856), .A2(N2391) );
  AND2_X1 AND2_670( .ZN(N2632), .A1(N1863), .A2(N2391) );
  AND2_X1 AND2_671( .ZN(N2633), .A1(N1880), .A2(N2395) );
  AND2_X1 AND2_672( .ZN(N2634), .A1(N1676), .A2(N2395) );
  AND2_X1 AND2_673( .ZN(N2635), .A1(N1681), .A2(N2395) );
  AND2_X1 AND2_674( .ZN(N2636), .A1(N1891), .A2(N2395) );
  INV_X1 NOT1_675( .ZN(N2638), .A(N2382) );
  BUF_X1 BUFF1_676( .Z(N2643), .A(N2521) );
  BUF_X1 BUFF1_677( .Z(N2644), .A(N2521) );
  INV_X1 NOT1_678( .ZN(N2645), .A(N2475) );
  INV_X1 NOT1_679( .ZN(N2646), .A(N2391) );
  NAND2_X1 NAND2_680( .ZN(N2652), .A1(N2528), .A2(N2400) );
  INV_X1 NOT1_681( .ZN(N2655), .A(N2478) );
  INV_X1 NOT1_682( .ZN(N2656), .A(N2481) );
  BUF_X1 BUFF1_683( .Z(N2659), .A(N2359) );
  INV_X1 NOT1_684( .ZN(N2663), .A(N2484) );
  NAND2_X1 NAND2_685( .ZN(N2664), .A1(N2484), .A2(N2301) );
  INV_X1 NOT1_686( .ZN(N2665), .A(N2553) );
  INV_X1 NOT1_687( .ZN(N2666), .A(N2552) );
  INV_X1 NOT1_688( .ZN(N2667), .A(N2551) );
  INV_X1 NOT1_689( .ZN(N2668), .A(N2550) );
  INV_X1 NOT1_690( .ZN(N2669), .A(N2549) );
  INV_X1 NOT1_691( .ZN(N2670), .A(N2548) );
  INV_X1 NOT1_692( .ZN(N2671), .A(N2547) );
  INV_X1 NOT1_693( .ZN(N2672), .A(N2546) );
  INV_X1 NOT1_694( .ZN(N2673), .A(N2545) );
  INV_X1 NOT1_695( .ZN(N2674), .A(N2544) );
  INV_X1 NOT1_696( .ZN(N2675), .A(N2568) );
  INV_X1 NOT1_697( .ZN(N2676), .A(N2567) );
  INV_X1 NOT1_698( .ZN(N2677), .A(N2566) );
  INV_X1 NOT1_699( .ZN(N2678), .A(N2565) );
  INV_X1 NOT1_700( .ZN(N2679), .A(N2564) );
  INV_X1 NOT1_701( .ZN(N2680), .A(N2563) );
  INV_X1 NOT1_702( .ZN(N2681), .A(N2417) );
  INV_X1 NOT1_703( .ZN(N2684), .A(N2421) );
  BUF_X8 BUFF1_704( .Z(N2687), .A(N2425) );
  BUF_X1 BUFF1_705( .Z(N2690), .A(N2425) );
  INV_X1 NOT1_706( .ZN(N2693), .A(N2493) );
  NAND2_X2 NAND2_707( .ZN(N2694), .A1(N2493), .A2(N1807) );
  INV_X1 NOT1_708( .ZN(N2695), .A(N2440) );
  INV_X1 NOT1_709( .ZN(N2696), .A(N2443) );
  INV_X1 NOT1_710( .ZN(N2697), .A(N2446) );
  INV_X1 NOT1_711( .ZN(N2698), .A(N2449) );
  INV_X1 NOT1_712( .ZN(N2699), .A(N2457) );
  INV_X1 NOT1_713( .ZN(N2700), .A(N2460) );
  INV_X1 NOT1_714( .ZN(N2701), .A(N2463) );
  INV_X1 NOT1_715( .ZN(N2702), .A(N2466) );
  NAND2_X1 NAND2_716( .ZN(N2703), .A1(N2579), .A2(N2453) );
  INV_X1 NOT1_717( .ZN(N2706), .A(N2469) );
  INV_X1 NOT1_718( .ZN(N2707), .A(N2487) );
  INV_X1 NOT1_719( .ZN(N2708), .A(N2490) );
  AND2_X1 AND2_720( .ZN(N2709), .A1(N2294), .A2(N2534) );
  AND2_X1 AND2_721( .ZN(N2710), .A1(N2291), .A2(N2531) );
  NAND2_X1 NAND2_722( .ZN(N2719), .A1(N2191), .A2(N2617) );
  NAND2_X1 NAND2_723( .ZN(N2720), .A1(N2194), .A2(N2620) );
  NAND2_X1 NAND2_724( .ZN(N2726), .A1(N2207), .A2(N2628) );
  BUF_X1 BUFF1_725( .Z(N2729), .A(N2537) );
  BUF_X1 BUFF1_726( .Z(N2738), .A(N2537) );
  INV_X1 NOT1_727( .ZN(N2743), .A(N2652) );
  NAND2_X1 NAND2_728( .ZN(N2747), .A1(N2049), .A2(N2663) );
  AND4_X1 AND5_729_A( .ZN(extra0), .A1(N2665), .A2(N2666), .A3(N2667), .A4(N2668) );
  AND2_X1 AND5_729( .ZN(N2748), .A1(extra0), .A2(N2669) );
  AND4_X1 AND5_730_A( .ZN(extra1), .A1(N2670), .A2(N2671), .A3(N2672), .A4(N2673) );
  AND2_X1 AND5_730( .ZN(N2749), .A1(extra1), .A2(N2674) );
  AND2_X1 AND2_731( .ZN(N2750), .A1(N2034), .A2(N2675) );
  AND4_X1 AND5_732_A( .ZN(extra2), .A1(N2676), .A2(N2677), .A3(N2678), .A4(N2679) );
  AND2_X1 AND5_732( .ZN(N2751), .A1(extra2), .A2(N2680) );
  NAND2_X1 NAND2_733( .ZN(N2760), .A1(N1588), .A2(N2693) );
  BUF_X1 BUFF1_734( .Z(N2761), .A(N2540) );
  BUF_X1 BUFF1_735( .Z(N2766), .A(N2540) );
  NAND2_X1 NAND2_736( .ZN(N2771), .A1(N2443), .A2(N2695) );
  NAND2_X1 NAND2_737( .ZN(N2772), .A1(N2440), .A2(N2696) );
  NAND2_X1 NAND2_738( .ZN(N2773), .A1(N2449), .A2(N2697) );
  NAND2_X1 NAND2_739( .ZN(N2774), .A1(N2446), .A2(N2698) );
  NAND2_X1 NAND2_740( .ZN(N2775), .A1(N2460), .A2(N2699) );
  NAND2_X1 NAND2_741( .ZN(N2776), .A1(N2457), .A2(N2700) );
  NAND2_X1 NAND2_742( .ZN(N2777), .A1(N2466), .A2(N2701) );
  NAND2_X1 NAND2_743( .ZN(N2778), .A1(N2463), .A2(N2702) );
  NAND2_X1 NAND2_744( .ZN(N2781), .A1(N2490), .A2(N2707) );
  NAND2_X1 NAND2_745( .ZN(N2782), .A1(N2487), .A2(N2708) );
  OR2_X1 OR2_746( .ZN(N2783), .A1(N2709), .A2(N2534) );
  OR2_X1 OR2_747( .ZN(N2784), .A1(N2710), .A2(N2531) );
  AND2_X2 AND2_748( .ZN(N2789), .A1(N1856), .A2(N2638) );
  AND2_X1 AND2_749( .ZN(N2790), .A1(N1863), .A2(N2638) );
  AND2_X1 AND2_750( .ZN(N2791), .A1(N1870), .A2(N2638) );
  AND2_X1 AND2_751( .ZN(N2792), .A1(N1875), .A2(N2638) );
  INV_X1 NOT1_752( .ZN(N2793), .A(N2613) );
  NAND2_X1 NAND2_753( .ZN(N2796), .A1(N2719), .A2(N2618) );
  NAND2_X1 NAND2_754( .ZN(N2800), .A1(N2619), .A2(N2720) );
  INV_X1 NOT1_755( .ZN(N2803), .A(N2624) );
  NAND2_X1 NAND2_756( .ZN(N2806), .A1(N2726), .A2(N2629) );
  AND2_X1 AND2_757( .ZN(N2809), .A1(N1856), .A2(N2646) );
  AND2_X1 AND2_758( .ZN(N2810), .A1(N1863), .A2(N2646) );
  AND2_X1 AND2_759( .ZN(N2811), .A1(N1870), .A2(N2646) );
  AND2_X1 AND2_760( .ZN(N2812), .A1(N1875), .A2(N2646) );
  AND2_X1 AND2_761( .ZN(N2817), .A1(N2743), .A2(N14) );
  BUF_X1 BUFF1_762( .Z(N2820), .A(N2603) );
  NAND2_X1 NAND2_763( .ZN(N2826), .A1(N2747), .A2(N2664) );
  AND2_X1 AND2_764( .ZN(N2829), .A1(N2748), .A2(N2749) );
  AND2_X1 AND2_765( .ZN(N2830), .A1(N2750), .A2(N2751) );
  BUF_X1 BUFF1_766( .Z(N2831), .A(N2659) );
  INV_X1 NOT1_767( .ZN(N2837), .A(N2687) );
  INV_X1 NOT1_768( .ZN(N2838), .A(N2690) );
  AND3_X1 AND3_769( .ZN(N2839), .A1(N2421), .A2(N2417), .A3(N2687) );
  AND3_X1 AND3_770( .ZN(N2840), .A1(N2684), .A2(N2681), .A3(N2690) );
  NAND2_X1 NAND2_771( .ZN(N2841), .A1(N2760), .A2(N2694) );
  BUF_X1 BUFF1_772( .Z(N2844), .A(N2603) );
  BUF_X1 BUFF1_773( .Z(N2854), .A(N2603) );
  BUF_X1 BUFF1_774( .Z(N2859), .A(N2659) );
  BUF_X1 BUFF1_775( .Z(N2869), .A(N2659) );
  NAND2_X1 NAND2_776( .ZN(N2874), .A1(N2773), .A2(N2774) );
  NAND2_X1 NAND2_777( .ZN(N2877), .A1(N2771), .A2(N2772) );
  INV_X1 NOT1_778( .ZN(N2880), .A(N2703) );
  NAND2_X1 NAND2_779( .ZN(N2881), .A1(N2703), .A2(N2706) );
  NAND2_X1 NAND2_780( .ZN(N2882), .A1(N2777), .A2(N2778) );
  NAND2_X1 NAND2_781( .ZN(N2885), .A1(N2775), .A2(N2776) );
  NAND2_X1 NAND2_782( .ZN(N2888), .A1(N2781), .A2(N2782) );
  NAND2_X1 NAND2_783( .ZN(N2891), .A1(N2783), .A2(N2784) );
  AND2_X1 AND2_784( .ZN(N2894), .A1(N2607), .A2(N2729) );
  AND2_X1 AND2_785( .ZN(N2895), .A1(N2608), .A2(N2729) );
  AND2_X1 AND2_786( .ZN(N2896), .A1(N2609), .A2(N2729) );
  AND2_X1 AND2_787( .ZN(N2897), .A1(N2610), .A2(N2729) );
  OR2_X1 OR2_788( .ZN(N2898), .A1(N2789), .A2(N2611) );
  OR2_X1 OR2_789( .ZN(N2899), .A1(N2790), .A2(N2612) );
  AND2_X1 AND2_790( .ZN(N2900), .A1(N2791), .A2(N1037) );
  AND2_X1 AND2_791( .ZN(N2901), .A1(N2792), .A2(N1037) );
  OR2_X1 OR2_792( .ZN(N2914), .A1(N2809), .A2(N2631) );
  OR2_X1 OR2_793( .ZN(N2915), .A1(N2810), .A2(N2632) );
  AND2_X1 AND2_794( .ZN(N2916), .A1(N2811), .A2(N1070) );
  AND2_X1 AND2_795( .ZN(N2917), .A1(N2812), .A2(N1070) );
  AND2_X1 AND2_796( .ZN(N2918), .A1(N2633), .A2(N2738) );
  AND2_X1 AND2_797( .ZN(N2919), .A1(N2634), .A2(N2738) );
  AND2_X1 AND2_798( .ZN(N2920), .A1(N2635), .A2(N2738) );
  AND2_X1 AND2_799( .ZN(N2921), .A1(N2636), .A2(N2738) );
  BUF_X8 BUFF1_800( .Z(N2925), .A(N2817) );
  AND3_X1 AND3_801( .ZN(N2931), .A1(N2829), .A2(N2830), .A3(N1302) );
  AND3_X1 AND3_802( .ZN(N2938), .A1(N2681), .A2(N2421), .A3(N2837) );
  AND3_X1 AND3_803( .ZN(N2939), .A1(N2417), .A2(N2684), .A3(N2838) );
  NAND2_X1 NAND2_804( .ZN(N2963), .A1(N2469), .A2(N2880) );
  INV_X4 NOT1_805( .ZN(N2970), .A(N2841) );
  INV_X4 NOT1_806( .ZN(N2971), .A(N2826) );
  INV_X1 NOT1_807( .ZN(N2972), .A(N2894) );
  INV_X1 NOT1_808( .ZN(N2975), .A(N2895) );
  INV_X1 NOT1_809( .ZN(N2978), .A(N2896) );
  INV_X1 NOT1_810( .ZN(N2981), .A(N2897) );
  AND2_X1 AND2_811( .ZN(N2984), .A1(N2898), .A2(N1037) );
  AND2_X1 AND2_812( .ZN(N2985), .A1(N2899), .A2(N1037) );
  INV_X1 NOT1_813( .ZN(N2986), .A(N2900) );
  INV_X1 NOT1_814( .ZN(N2989), .A(N2901) );
  INV_X1 NOT1_815( .ZN(N2992), .A(N2796) );
  BUF_X8 BUFF1_816( .Z(N2995), .A(N2800) );
  BUF_X1 BUFF1_817( .Z(N2998), .A(N2800) );
  BUF_X1 BUFF1_818( .Z(N3001), .A(N2806) );
  BUF_X1 BUFF1_819( .Z(N3004), .A(N2806) );
  AND2_X1 AND2_820( .ZN(N3007), .A1(N574), .A2(N2820) );
  AND2_X1 AND2_821( .ZN(N3008), .A1(N2914), .A2(N1070) );
  AND2_X1 AND2_822( .ZN(N3009), .A1(N2915), .A2(N1070) );
  INV_X1 NOT1_823( .ZN(N3010), .A(N2916) );
  INV_X1 NOT1_824( .ZN(N3013), .A(N2917) );
  INV_X1 NOT1_825( .ZN(N3016), .A(N2918) );
  INV_X1 NOT1_826( .ZN(N3019), .A(N2919) );
  INV_X1 NOT1_827( .ZN(N3022), .A(N2920) );
  INV_X1 NOT1_828( .ZN(N3025), .A(N2921) );
  INV_X1 NOT1_829( .ZN(N3028), .A(N2817) );
  AND2_X1 AND2_830( .ZN(N3029), .A1(N574), .A2(N2831) );
  INV_X1 NOT1_831( .ZN(N3030), .A(N2820) );
  AND2_X1 AND2_832( .ZN(N3035), .A1(N578), .A2(N2820) );
  AND2_X1 AND2_833( .ZN(N3036), .A1(N655), .A2(N2820) );
  AND2_X1 AND2_834( .ZN(N3037), .A1(N659), .A2(N2820) );
  BUF_X1 BUFF1_835( .Z(N3038), .A(N2931) );
  INV_X1 NOT1_836( .ZN(N3039), .A(N2831) );
  AND2_X1 AND2_837( .ZN(N3044), .A1(N578), .A2(N2831) );
  AND2_X1 AND2_838( .ZN(N3045), .A1(N655), .A2(N2831) );
  AND2_X1 AND2_839( .ZN(N3046), .A1(N659), .A2(N2831) );
  NOR2_X1 NOR2_840( .ZN(N3047), .A1(N2938), .A2(N2839) );
  NOR2_X1 NOR2_841( .ZN(N3048), .A1(N2939), .A2(N2840) );
  INV_X1 NOT1_842( .ZN(N3049), .A(N2888) );
  INV_X1 NOT1_843( .ZN(N3050), .A(N2844) );
  AND2_X2 AND2_844( .ZN(N3053), .A1(N663), .A2(N2844) );
  AND2_X2 AND2_845( .ZN(N3054), .A1(N667), .A2(N2844) );
  AND2_X2 AND2_846( .ZN(N3055), .A1(N671), .A2(N2844) );
  AND2_X1 AND2_847( .ZN(N3056), .A1(N675), .A2(N2844) );
  AND2_X1 AND2_848( .ZN(N3057), .A1(N679), .A2(N2854) );
  AND2_X1 AND2_849( .ZN(N3058), .A1(N683), .A2(N2854) );
  AND2_X1 AND2_850( .ZN(N3059), .A1(N687), .A2(N2854) );
  AND2_X1 AND2_851( .ZN(N3060), .A1(N705), .A2(N2854) );
  INV_X1 NOT1_852( .ZN(N3061), .A(N2859) );
  AND2_X1 AND2_853( .ZN(N3064), .A1(N663), .A2(N2859) );
  AND2_X1 AND2_854( .ZN(N3065), .A1(N667), .A2(N2859) );
  AND2_X1 AND2_855( .ZN(N3066), .A1(N671), .A2(N2859) );
  AND2_X1 AND2_856( .ZN(N3067), .A1(N675), .A2(N2859) );
  AND2_X1 AND2_857( .ZN(N3068), .A1(N679), .A2(N2869) );
  AND2_X1 AND2_858( .ZN(N3069), .A1(N683), .A2(N2869) );
  AND2_X1 AND2_859( .ZN(N3070), .A1(N687), .A2(N2869) );
  AND2_X1 AND2_860( .ZN(N3071), .A1(N705), .A2(N2869) );
  INV_X1 NOT1_861( .ZN(N3072), .A(N2874) );
  INV_X1 NOT1_862( .ZN(N3073), .A(N2877) );
  INV_X1 NOT1_863( .ZN(N3074), .A(N2882) );
  INV_X1 NOT1_864( .ZN(N3075), .A(N2885) );
  NAND2_X1 NAND2_865( .ZN(N3076), .A1(N2881), .A2(N2963) );
  INV_X1 NOT1_866( .ZN(N3079), .A(N2931) );
  INV_X1 NOT1_867( .ZN(N3088), .A(N2984) );
  INV_X1 NOT1_868( .ZN(N3091), .A(N2985) );
  INV_X1 NOT1_869( .ZN(N3110), .A(N3008) );
  INV_X1 NOT1_870( .ZN(N3113), .A(N3009) );
  AND2_X1 AND2_871( .ZN(N3137), .A1(N3055), .A2(N1190) );
  AND2_X1 AND2_872( .ZN(N3140), .A1(N3056), .A2(N1190) );
  AND2_X1 AND2_873( .ZN(N3143), .A1(N3057), .A2(N2761) );
  AND2_X1 AND2_874( .ZN(N3146), .A1(N3058), .A2(N2761) );
  AND2_X1 AND2_875( .ZN(N3149), .A1(N3059), .A2(N2761) );
  AND2_X1 AND2_876( .ZN(N3152), .A1(N3060), .A2(N2761) );
  AND2_X1 AND2_877( .ZN(N3157), .A1(N3066), .A2(N1195) );
  AND2_X1 AND2_878( .ZN(N3160), .A1(N3067), .A2(N1195) );
  AND2_X1 AND2_879( .ZN(N3163), .A1(N3068), .A2(N2766) );
  AND2_X1 AND2_880( .ZN(N3166), .A1(N3069), .A2(N2766) );
  AND2_X1 AND2_881( .ZN(N3169), .A1(N3070), .A2(N2766) );
  AND2_X1 AND2_882( .ZN(N3172), .A1(N3071), .A2(N2766) );
  NAND2_X2 NAND2_883( .ZN(N3175), .A1(N2877), .A2(N3072) );
  NAND2_X2 NAND2_884( .ZN(N3176), .A1(N2874), .A2(N3073) );
  NAND2_X2 NAND2_885( .ZN(N3177), .A1(N2885), .A2(N3074) );
  NAND2_X1 NAND2_886( .ZN(N3178), .A1(N2882), .A2(N3075) );
  NAND2_X1 NAND2_887( .ZN(N3180), .A1(N3048), .A2(N3047) );
  INV_X1 NOT1_888( .ZN(N3187), .A(N2995) );
  INV_X1 NOT1_889( .ZN(N3188), .A(N2998) );
  INV_X1 NOT1_890( .ZN(N3189), .A(N3001) );
  INV_X1 NOT1_891( .ZN(N3190), .A(N3004) );
  AND3_X1 AND3_892( .ZN(N3191), .A1(N2796), .A2(N2613), .A3(N2995) );
  AND3_X1 AND3_893( .ZN(N3192), .A1(N2992), .A2(N2793), .A3(N2998) );
  AND3_X1 AND3_894( .ZN(N3193), .A1(N2624), .A2(N2368), .A3(N3001) );
  AND3_X1 AND3_895( .ZN(N3194), .A1(N2803), .A2(N2621), .A3(N3004) );
  NAND2_X1 NAND2_896( .ZN(N3195), .A1(N3076), .A2(N2375) );
  INV_X1 NOT1_897( .ZN(N3196), .A(N3076) );
  AND2_X1 AND2_898( .ZN(N3197), .A1(N687), .A2(N3030) );
  AND2_X1 AND2_899( .ZN(N3208), .A1(N687), .A2(N3039) );
  AND2_X1 AND2_900( .ZN(N3215), .A1(N705), .A2(N3030) );
  AND2_X1 AND2_901( .ZN(N3216), .A1(N711), .A2(N3030) );
  AND2_X1 AND2_902( .ZN(N3217), .A1(N715), .A2(N3030) );
  AND2_X1 AND2_903( .ZN(N3218), .A1(N705), .A2(N3039) );
  AND2_X1 AND2_904( .ZN(N3219), .A1(N711), .A2(N3039) );
  AND2_X1 AND2_905( .ZN(N3220), .A1(N715), .A2(N3039) );
  AND2_X1 AND2_906( .ZN(N3222), .A1(N719), .A2(N3050) );
  AND2_X1 AND2_907( .ZN(N3223), .A1(N723), .A2(N3050) );
  AND2_X1 AND2_908( .ZN(N3230), .A1(N719), .A2(N3061) );
  AND2_X1 AND2_909( .ZN(N3231), .A1(N723), .A2(N3061) );
  NAND2_X1 NAND2_910( .ZN(N3238), .A1(N3175), .A2(N3176) );
  NAND2_X1 NAND2_911( .ZN(N3241), .A1(N3177), .A2(N3178) );
  BUF_X1 BUFF1_912( .Z(N3244), .A(N2981) );
  BUF_X1 BUFF1_913( .Z(N3247), .A(N2978) );
  BUF_X1 BUFF1_914( .Z(N3250), .A(N2975) );
  BUF_X1 BUFF1_915( .Z(N3253), .A(N2972) );
  BUF_X1 BUFF1_916( .Z(N3256), .A(N2989) );
  BUF_X1 BUFF1_917( .Z(N3259), .A(N2986) );
  BUF_X1 BUFF1_918( .Z(N3262), .A(N3025) );
  BUF_X1 BUFF1_919( .Z(N3265), .A(N3022) );
  BUF_X1 BUFF1_920( .Z(N3268), .A(N3019) );
  BUF_X1 BUFF1_921( .Z(N3271), .A(N3016) );
  BUF_X1 BUFF1_922( .Z(N3274), .A(N3013) );
  BUF_X1 BUFF1_923( .Z(N3277), .A(N3010) );
  AND3_X1 AND3_924( .ZN(N3281), .A1(N2793), .A2(N2796), .A3(N3187) );
  AND3_X1 AND3_925( .ZN(N3282), .A1(N2613), .A2(N2992), .A3(N3188) );
  AND3_X1 AND3_926( .ZN(N3283), .A1(N2621), .A2(N2624), .A3(N3189) );
  AND3_X1 AND3_927( .ZN(N3284), .A1(N2368), .A2(N2803), .A3(N3190) );
  NAND2_X1 NAND2_928( .ZN(N3286), .A1(N2210), .A2(N3196) );
  OR2_X1 OR2_929( .ZN(N3288), .A1(N3197), .A2(N3007) );
  NAND2_X1 NAND2_930( .ZN(N3289), .A1(N3180), .A2(N3049) );
  AND2_X1 AND2_931( .ZN(N3291), .A1(N3152), .A2(N2981) );
  AND2_X1 AND2_932( .ZN(N3293), .A1(N3149), .A2(N2978) );
  AND2_X1 AND2_933( .ZN(N3295), .A1(N3146), .A2(N2975) );
  AND2_X1 AND2_934( .ZN(N3296), .A1(N2972), .A2(N3143) );
  AND2_X2 AND2_935( .ZN(N3299), .A1(N3140), .A2(N2989) );
  AND2_X2 AND2_936( .ZN(N3301), .A1(N3137), .A2(N2986) );
  OR2_X1 OR2_937( .ZN(N3302), .A1(N3208), .A2(N3029) );
  AND2_X1 AND2_938( .ZN(N3304), .A1(N3172), .A2(N3025) );
  AND2_X1 AND2_939( .ZN(N3306), .A1(N3169), .A2(N3022) );
  AND2_X1 AND2_940( .ZN(N3308), .A1(N3166), .A2(N3019) );
  AND2_X1 AND2_941( .ZN(N3309), .A1(N3016), .A2(N3163) );
  AND2_X1 AND2_942( .ZN(N3312), .A1(N3160), .A2(N3013) );
  AND2_X1 AND2_943( .ZN(N3314), .A1(N3157), .A2(N3010) );
  OR2_X1 OR2_944( .ZN(N3315), .A1(N3215), .A2(N3035) );
  OR2_X2 OR2_945( .ZN(N3318), .A1(N3216), .A2(N3036) );
  OR2_X4 OR2_946( .ZN(N3321), .A1(N3217), .A2(N3037) );
  OR2_X1 OR2_947( .ZN(N3324), .A1(N3218), .A2(N3044) );
  OR2_X1 OR2_948( .ZN(N3327), .A1(N3219), .A2(N3045) );
  OR2_X1 OR2_949( .ZN(N3330), .A1(N3220), .A2(N3046) );
  INV_X4 NOT1_950( .ZN(N3333), .A(N3180) );
  OR2_X1 OR2_951( .ZN(N3334), .A1(N3222), .A2(N3053) );
  OR2_X1 OR2_952( .ZN(N3335), .A1(N3223), .A2(N3054) );
  OR2_X2 OR2_953( .ZN(N3336), .A1(N3230), .A2(N3064) );
  OR2_X1 OR2_954( .ZN(N3337), .A1(N3231), .A2(N3065) );
  BUF_X1 BUFF1_955( .Z(N3340), .A(N3152) );
  BUF_X1 BUFF1_956( .Z(N3344), .A(N3149) );
  BUF_X1 BUFF1_957( .Z(N3348), .A(N3146) );
  BUF_X1 BUFF1_958( .Z(N3352), .A(N3143) );
  BUF_X2 BUFF1_959( .Z(N3356), .A(N3140) );
  BUF_X2 BUFF1_960( .Z(N3360), .A(N3137) );
  BUF_X2 BUFF1_961( .Z(N3364), .A(N3091) );
  BUF_X1 BUFF1_962( .Z(N3367), .A(N3088) );
  BUF_X1 BUFF1_963( .Z(N3370), .A(N3172) );
  BUF_X1 BUFF1_964( .Z(N3374), .A(N3169) );
  BUF_X1 BUFF1_965( .Z(N3378), .A(N3166) );
  BUF_X1 BUFF1_966( .Z(N3382), .A(N3163) );
  BUF_X1 BUFF1_967( .Z(N3386), .A(N3160) );
  BUF_X1 BUFF1_968( .Z(N3390), .A(N3157) );
  BUF_X1 BUFF1_969( .Z(N3394), .A(N3113) );
  BUF_X1 BUFF1_970( .Z(N3397), .A(N3110) );
  NAND2_X1 NAND2_971( .ZN(N3400), .A1(N3195), .A2(N3286) );
  NOR2_X1 NOR2_972( .ZN(N3401), .A1(N3281), .A2(N3191) );
  NOR2_X1 NOR2_973( .ZN(N3402), .A1(N3282), .A2(N3192) );
  NOR2_X1 NOR2_974( .ZN(N3403), .A1(N3283), .A2(N3193) );
  NOR2_X1 NOR2_975( .ZN(N3404), .A1(N3284), .A2(N3194) );
  INV_X1 NOT1_976( .ZN(N3405), .A(N3238) );
  INV_X1 NOT1_977( .ZN(N3406), .A(N3241) );
  AND2_X1 AND2_978( .ZN(N3409), .A1(N3288), .A2(N1836) );
  NAND2_X1 NAND2_979( .ZN(N3410), .A1(N2888), .A2(N3333) );
  INV_X1 NOT1_980( .ZN(N3412), .A(N3244) );
  INV_X1 NOT1_981( .ZN(N3414), .A(N3247) );
  INV_X1 NOT1_982( .ZN(N3416), .A(N3250) );
  INV_X1 NOT1_983( .ZN(N3418), .A(N3253) );
  INV_X1 NOT1_984( .ZN(N3420), .A(N3256) );
  INV_X1 NOT1_985( .ZN(N3422), .A(N3259) );
  AND2_X1 AND2_986( .ZN(N3428), .A1(N3302), .A2(N1836) );
  INV_X1 NOT1_987( .ZN(N3430), .A(N3262) );
  INV_X1 NOT1_988( .ZN(N3432), .A(N3265) );
  INV_X1 NOT1_989( .ZN(N3434), .A(N3268) );
  INV_X1 NOT1_990( .ZN(N3436), .A(N3271) );
  INV_X1 NOT1_991( .ZN(N3438), .A(N3274) );
  INV_X1 NOT1_992( .ZN(N3440), .A(N3277) );
  AND2_X1 AND2_993( .ZN(N3450), .A1(N3334), .A2(N1190) );
  AND2_X1 AND2_994( .ZN(N3453), .A1(N3335), .A2(N1190) );
  AND2_X1 AND2_995( .ZN(N3456), .A1(N3336), .A2(N1195) );
  AND2_X1 AND2_996( .ZN(N3459), .A1(N3337), .A2(N1195) );
  AND2_X1 AND2_997( .ZN(N3478), .A1(N3400), .A2(N533) );
  AND2_X1 AND2_998( .ZN(N3479), .A1(N3318), .A2(N2128) );
  AND2_X1 AND2_999( .ZN(N3480), .A1(N3315), .A2(N1841) );
  NAND2_X1 NAND2_1000( .ZN(N3481), .A1(N3410), .A2(N3289) );
  INV_X1 NOT1_1001( .ZN(N3482), .A(N3340) );
  NAND2_X1 NAND2_1002( .ZN(N3483), .A1(N3340), .A2(N3412) );
  INV_X1 NOT1_1003( .ZN(N3484), .A(N3344) );
  NAND2_X1 NAND2_1004( .ZN(N3485), .A1(N3344), .A2(N3414) );
  INV_X1 NOT1_1005( .ZN(N3486), .A(N3348) );
  NAND2_X1 NAND2_1006( .ZN(N3487), .A1(N3348), .A2(N3416) );
  INV_X1 NOT1_1007( .ZN(N3488), .A(N3352) );
  NAND2_X1 NAND2_1008( .ZN(N3489), .A1(N3352), .A2(N3418) );
  INV_X1 NOT1_1009( .ZN(N3490), .A(N3356) );
  NAND2_X1 NAND2_1010( .ZN(N3491), .A1(N3356), .A2(N3420) );
  INV_X1 NOT1_1011( .ZN(N3492), .A(N3360) );
  NAND2_X1 NAND2_1012( .ZN(N3493), .A1(N3360), .A2(N3422) );
  INV_X1 NOT1_1013( .ZN(N3494), .A(N3364) );
  INV_X1 NOT1_1014( .ZN(N3496), .A(N3367) );
  AND2_X1 AND2_1015( .ZN(N3498), .A1(N3321), .A2(N2135) );
  AND2_X1 AND2_1016( .ZN(N3499), .A1(N3327), .A2(N2128) );
  AND2_X1 AND2_1017( .ZN(N3500), .A1(N3324), .A2(N1841) );
  INV_X1 NOT1_1018( .ZN(N3501), .A(N3370) );
  NAND2_X1 NAND2_1019( .ZN(N3502), .A1(N3370), .A2(N3430) );
  INV_X1 NOT1_1020( .ZN(N3503), .A(N3374) );
  NAND2_X1 NAND2_1021( .ZN(N3504), .A1(N3374), .A2(N3432) );
  INV_X1 NOT1_1022( .ZN(N3505), .A(N3378) );
  NAND2_X1 NAND2_1023( .ZN(N3506), .A1(N3378), .A2(N3434) );
  INV_X1 NOT1_1024( .ZN(N3507), .A(N3382) );
  NAND2_X2 NAND2_1025( .ZN(N3508), .A1(N3382), .A2(N3436) );
  INV_X1 NOT1_1026( .ZN(N3509), .A(N3386) );
  NAND2_X1 NAND2_1027( .ZN(N3510), .A1(N3386), .A2(N3438) );
  INV_X1 NOT1_1028( .ZN(N3511), .A(N3390) );
  NAND2_X1 NAND2_1029( .ZN(N3512), .A1(N3390), .A2(N3440) );
  INV_X1 NOT1_1030( .ZN(N3513), .A(N3394) );
  INV_X1 NOT1_1031( .ZN(N3515), .A(N3397) );
  AND2_X2 AND2_1032( .ZN(N3517), .A1(N3330), .A2(N2135) );
  NAND2_X1 NAND2_1033( .ZN(N3522), .A1(N3402), .A2(N3401) );
  NAND2_X1 NAND2_1034( .ZN(N3525), .A1(N3404), .A2(N3403) );
  BUF_X1 BUFF1_1035( .Z(N3528), .A(N3318) );
  BUF_X1 BUFF1_1036( .Z(N3531), .A(N3315) );
  BUF_X1 BUFF1_1037( .Z(N3534), .A(N3321) );
  BUF_X1 BUFF1_1038( .Z(N3537), .A(N3327) );
  BUF_X1 BUFF1_1039( .Z(N3540), .A(N3324) );
  BUF_X1 BUFF1_1040( .Z(N3543), .A(N3330) );
  OR2_X1 OR2_1041( .ZN(N3546), .A1(N3478), .A2(N1813) );
  INV_X1 NOT1_1042( .ZN(N3551), .A(N3481) );
  NAND2_X1 NAND2_1043( .ZN(N3552), .A1(N3244), .A2(N3482) );
  NAND2_X1 NAND2_1044( .ZN(N3553), .A1(N3247), .A2(N3484) );
  NAND2_X1 NAND2_1045( .ZN(N3554), .A1(N3250), .A2(N3486) );
  NAND2_X1 NAND2_1046( .ZN(N3555), .A1(N3253), .A2(N3488) );
  NAND2_X1 NAND2_1047( .ZN(N3556), .A1(N3256), .A2(N3490) );
  NAND2_X1 NAND2_1048( .ZN(N3557), .A1(N3259), .A2(N3492) );
  AND2_X1 AND2_1049( .ZN(N3558), .A1(N3453), .A2(N3091) );
  AND2_X1 AND2_1050( .ZN(N3559), .A1(N3450), .A2(N3088) );
  NAND2_X1 NAND2_1051( .ZN(N3563), .A1(N3262), .A2(N3501) );
  NAND2_X1 NAND2_1052( .ZN(N3564), .A1(N3265), .A2(N3503) );
  NAND2_X1 NAND2_1053( .ZN(N3565), .A1(N3268), .A2(N3505) );
  NAND2_X1 NAND2_1054( .ZN(N3566), .A1(N3271), .A2(N3507) );
  NAND2_X1 NAND2_1055( .ZN(N3567), .A1(N3274), .A2(N3509) );
  NAND2_X1 NAND2_1056( .ZN(N3568), .A1(N3277), .A2(N3511) );
  AND2_X1 AND2_1057( .ZN(N3569), .A1(N3459), .A2(N3113) );
  AND2_X1 AND2_1058( .ZN(N3570), .A1(N3456), .A2(N3110) );
  BUF_X1 BUFF1_1059( .Z(N3576), .A(N3453) );
  BUF_X1 BUFF1_1060( .Z(N3579), .A(N3450) );
  BUF_X1 BUFF1_1061( .Z(N3585), .A(N3459) );
  BUF_X1 BUFF1_1062( .Z(N3588), .A(N3456) );
  INV_X4 NOT1_1063( .ZN(N3592), .A(N3522) );
  NAND2_X1 NAND2_1064( .ZN(N3593), .A1(N3522), .A2(N3405) );
  INV_X1 NOT1_1065( .ZN(N3594), .A(N3525) );
  NAND2_X1 NAND2_1066( .ZN(N3595), .A1(N3525), .A2(N3406) );
  INV_X1 NOT1_1067( .ZN(N3596), .A(N3528) );
  NAND2_X1 NAND2_1068( .ZN(N3597), .A1(N3528), .A2(N2630) );
  NAND2_X1 NAND2_1069( .ZN(N3598), .A1(N3531), .A2(N2376) );
  INV_X1 NOT1_1070( .ZN(N3599), .A(N3531) );
  AND2_X1 AND2_1071( .ZN(N3600), .A1(N3551), .A2(N800) );
  NAND2_X1 NAND2_1072( .ZN(N3603), .A1(N3552), .A2(N3483) );
  NAND2_X1 NAND2_1073( .ZN(N3608), .A1(N3553), .A2(N3485) );
  NAND2_X1 NAND2_1074( .ZN(N3612), .A1(N3554), .A2(N3487) );
  NAND2_X1 NAND2_1075( .ZN(N3615), .A1(N3555), .A2(N3489) );
  NAND2_X1 NAND2_1076( .ZN(N3616), .A1(N3556), .A2(N3491) );
  NAND2_X1 NAND2_1077( .ZN(N3622), .A1(N3557), .A2(N3493) );
  INV_X1 NOT1_1078( .ZN(N3629), .A(N3534) );
  NAND2_X1 NAND2_1079( .ZN(N3630), .A1(N3534), .A2(N2645) );
  INV_X1 NOT1_1080( .ZN(N3631), .A(N3537) );
  NAND2_X1 NAND2_1081( .ZN(N3632), .A1(N3537), .A2(N2655) );
  NAND2_X1 NAND2_1082( .ZN(N3633), .A1(N3540), .A2(N2403) );
  INV_X1 NOT1_1083( .ZN(N3634), .A(N3540) );
  NAND2_X1 NAND2_1084( .ZN(N3635), .A1(N3563), .A2(N3502) );
  NAND2_X1 NAND2_1085( .ZN(N3640), .A1(N3564), .A2(N3504) );
  NAND2_X1 NAND2_1086( .ZN(N3644), .A1(N3565), .A2(N3506) );
  NAND2_X1 NAND2_1087( .ZN(N3647), .A1(N3566), .A2(N3508) );
  NAND2_X1 NAND2_1088( .ZN(N3648), .A1(N3567), .A2(N3510) );
  NAND2_X1 NAND2_1089( .ZN(N3654), .A1(N3568), .A2(N3512) );
  INV_X1 NOT1_1090( .ZN(N3661), .A(N3543) );
  NAND2_X1 NAND2_1091( .ZN(N3662), .A1(N3543), .A2(N2656) );
  NAND2_X1 NAND2_1092( .ZN(N3667), .A1(N3238), .A2(N3592) );
  NAND2_X1 NAND2_1093( .ZN(N3668), .A1(N3241), .A2(N3594) );
  NAND2_X1 NAND2_1094( .ZN(N3669), .A1(N2472), .A2(N3596) );
  NAND2_X1 NAND2_1095( .ZN(N3670), .A1(N2213), .A2(N3599) );
  BUF_X1 BUFF1_1096( .Z(N3671), .A(N3600) );
  INV_X1 NOT1_1097( .ZN(N3691), .A(N3576) );
  NAND2_X1 NAND2_1098( .ZN(N3692), .A1(N3576), .A2(N3494) );
  INV_X1 NOT1_1099( .ZN(N3693), .A(N3579) );
  NAND2_X1 NAND2_1100( .ZN(N3694), .A1(N3579), .A2(N3496) );
  NAND2_X1 NAND2_1101( .ZN(N3695), .A1(N2475), .A2(N3629) );
  NAND2_X1 NAND2_1102( .ZN(N3696), .A1(N2478), .A2(N3631) );
  NAND2_X1 NAND2_1103( .ZN(N3697), .A1(N2216), .A2(N3634) );
  INV_X1 NOT1_1104( .ZN(N3716), .A(N3585) );
  NAND2_X1 NAND2_1105( .ZN(N3717), .A1(N3585), .A2(N3513) );
  INV_X1 NOT1_1106( .ZN(N3718), .A(N3588) );
  NAND2_X1 NAND2_1107( .ZN(N3719), .A1(N3588), .A2(N3515) );
  NAND2_X1 NAND2_1108( .ZN(N3720), .A1(N2481), .A2(N3661) );
  NAND2_X1 NAND2_1109( .ZN(N3721), .A1(N3667), .A2(N3593) );
  NAND2_X1 NAND2_1110( .ZN(N3722), .A1(N3668), .A2(N3595) );
  NAND2_X1 NAND2_1111( .ZN(N3723), .A1(N3669), .A2(N3597) );
  NAND2_X1 NAND2_1112( .ZN(N3726), .A1(N3670), .A2(N3598) );
  INV_X1 NOT1_1113( .ZN(N3727), .A(N3600) );
  NAND2_X1 NAND2_1114( .ZN(N3728), .A1(N3364), .A2(N3691) );
  NAND2_X1 NAND2_1115( .ZN(N3729), .A1(N3367), .A2(N3693) );
  NAND2_X1 NAND2_1116( .ZN(N3730), .A1(N3695), .A2(N3630) );
  AND4_X1 AND4_1117( .ZN(N3731), .A1(N3608), .A2(N3615), .A3(N3612), .A4(N3603) );
  AND2_X1 AND2_1118( .ZN(N3732), .A1(N3603), .A2(N3293) );
  AND3_X1 AND3_1119( .ZN(N3733), .A1(N3608), .A2(N3603), .A3(N3295) );
  AND4_X1 AND4_1120( .ZN(N3734), .A1(N3612), .A2(N3603), .A3(N3296), .A4(N3608) );
  AND2_X1 AND2_1121( .ZN(N3735), .A1(N3616), .A2(N3301) );
  AND3_X1 AND3_1122( .ZN(N3736), .A1(N3622), .A2(N3616), .A3(N3558) );
  NAND2_X2 NAND2_1123( .ZN(N3737), .A1(N3696), .A2(N3632) );
  NAND2_X2 NAND2_1124( .ZN(N3740), .A1(N3697), .A2(N3633) );
  NAND2_X1 NAND2_1125( .ZN(N3741), .A1(N3394), .A2(N3716) );
  NAND2_X1 NAND2_1126( .ZN(N3742), .A1(N3397), .A2(N3718) );
  NAND2_X1 NAND2_1127( .ZN(N3743), .A1(N3720), .A2(N3662) );
  AND4_X1 AND4_1128( .ZN(N3744), .A1(N3640), .A2(N3647), .A3(N3644), .A4(N3635) );
  AND2_X1 AND2_1129( .ZN(N3745), .A1(N3635), .A2(N3306) );
  AND3_X1 AND3_1130( .ZN(N3746), .A1(N3640), .A2(N3635), .A3(N3308) );
  AND4_X1 AND4_1131( .ZN(N3747), .A1(N3644), .A2(N3635), .A3(N3309), .A4(N3640) );
  AND2_X1 AND2_1132( .ZN(N3748), .A1(N3648), .A2(N3314) );
  AND3_X1 AND3_1133( .ZN(N3749), .A1(N3654), .A2(N3648), .A3(N3569) );
  INV_X1 NOT1_1134( .ZN(N3750), .A(N3721) );
  AND2_X1 AND2_1135( .ZN(N3753), .A1(N3722), .A2(N246) );
  NAND2_X1 NAND2_1136( .ZN(N3754), .A1(N3728), .A2(N3692) );
  NAND2_X1 NAND2_1137( .ZN(N3758), .A1(N3729), .A2(N3694) );
  INV_X4 NOT1_1138( .ZN(N3761), .A(N3731) );
  OR4_X1 OR4_1139( .ZN(N3762), .A1(N3291), .A2(N3732), .A3(N3733), .A4(N3734) );
  NAND2_X1 NAND2_1140( .ZN(N3767), .A1(N3741), .A2(N3717) );
  NAND2_X1 NAND2_1141( .ZN(N3771), .A1(N3742), .A2(N3719) );
  INV_X1 NOT1_1142( .ZN(N3774), .A(N3744) );
  OR4_X1 OR4_1143( .ZN(N3775), .A1(N3304), .A2(N3745), .A3(N3746), .A4(N3747) );
  AND2_X1 AND2_1144( .ZN(N3778), .A1(N3723), .A2(N3480) );
  AND3_X1 AND3_1145( .ZN(N3779), .A1(N3726), .A2(N3723), .A3(N3409) );
  OR2_X1 OR2_1146( .ZN(N3780), .A1(N2125), .A2(N3753) );
  AND2_X1 AND2_1147( .ZN(N3790), .A1(N3750), .A2(N800) );
  AND2_X1 AND2_1148( .ZN(N3793), .A1(N3737), .A2(N3500) );
  AND3_X1 AND3_1149( .ZN(N3794), .A1(N3740), .A2(N3737), .A3(N3428) );
  OR3_X1 OR3_1150( .ZN(N3802), .A1(N3479), .A2(N3778), .A3(N3779) );
  BUF_X2 BUFF1_1151( .Z(N3803), .A(N3780) );
  BUF_X2 BUFF1_1152( .Z(N3804), .A(N3780) );
  INV_X1 NOT1_1153( .ZN(N3805), .A(N3762) );
  AND4_X1 AND5_1154_A( .ZN(extra3), .A1(N3622), .A2(N3730), .A3(N3754), .A4(N3616) );
  AND2_X1 AND5_1154( .ZN(N3806), .A1(extra3), .A2(N3758) );
  AND4_X1 AND4_1155( .ZN(N3807), .A1(N3754), .A2(N3616), .A3(N3559), .A4(N3622) );
  AND4_X1 AND5_1156_A( .ZN(extra4), .A1(N3758), .A2(N3754), .A3(N3616), .A4(N3498) );
  AND2_X1 AND5_1156( .ZN(N3808), .A1(extra4), .A2(N3622) );
  BUF_X1 BUFF1_1157( .Z(N3809), .A(N3790) );
  OR3_X1 OR3_1158( .ZN(N3811), .A1(N3499), .A2(N3793), .A3(N3794) );
  INV_X1 NOT1_1159( .ZN(N3812), .A(N3775) );
  AND4_X1 AND5_1160_A( .ZN(extra5), .A1(N3654), .A2(N3743), .A3(N3767), .A4(N3648) );
  AND2_X1 AND5_1160( .ZN(N3813), .A1(extra5), .A2(N3771) );
  AND4_X1 AND4_1161( .ZN(N3814), .A1(N3767), .A2(N3648), .A3(N3570), .A4(N3654) );
  AND4_X1 AND5_1162_A( .ZN(extra6), .A1(N3771), .A2(N3767), .A3(N3648), .A4(N3517) );
  AND2_X1 AND5_1162( .ZN(N3815), .A1(extra6), .A2(N3654) );
  OR4_X1 OR5_1163_A( .ZN(extra7), .A1(N3299), .A2(N3735), .A3(N3736), .A4(N3807) );
  OR2_X1 OR5_1163( .ZN(N3816), .A1(extra7), .A2(N3808) );
  AND2_X1 AND2_1164( .ZN(N3817), .A1(N3806), .A2(N3802) );
  NAND2_X1 NAND2_1165( .ZN(N3818), .A1(N3805), .A2(N3761) );
  INV_X1 NOT1_1166( .ZN(N3819), .A(N3790) );
  OR4_X1 OR5_1167_A( .ZN(extra8), .A1(N3312), .A2(N3748), .A3(N3749), .A4(N3814) );
  OR2_X1 OR5_1167( .ZN(N3820), .A1(extra8), .A2(N3815) );
  AND2_X1 AND2_1168( .ZN(N3821), .A1(N3813), .A2(N3811) );
  NAND2_X1 NAND2_1169( .ZN(N3822), .A1(N3812), .A2(N3774) );
  OR2_X1 OR2_1170( .ZN(N3823), .A1(N3816), .A2(N3817) );
  AND3_X1 AND3_1171( .ZN(N3826), .A1(N3727), .A2(N3819), .A3(N2841) );
  OR2_X1 OR2_1172( .ZN(N3827), .A1(N3820), .A2(N3821) );
  INV_X1 NOT1_1173( .ZN(N3834), .A(N3823) );
  AND2_X2 AND2_1174( .ZN(N3835), .A1(N3818), .A2(N3823) );
  INV_X1 NOT1_1175( .ZN(N3836), .A(N3827) );
  AND2_X1 AND2_1176( .ZN(N3837), .A1(N3822), .A2(N3827) );
  AND2_X1 AND2_1177( .ZN(N3838), .A1(N3762), .A2(N3834) );
  AND2_X1 AND2_1178( .ZN(N3839), .A1(N3775), .A2(N3836) );
  OR2_X1 OR2_1179( .ZN(N3840), .A1(N3838), .A2(N3835) );
  OR2_X2 OR2_1180( .ZN(N3843), .A1(N3839), .A2(N3837) );
  BUF_X1 BUFF1_1181( .Z(N3851), .A(N3843) );
  NAND2_X1 NAND2_1182( .ZN(N3852), .A1(N3843), .A2(N3840) );
  AND2_X1 AND2_1183( .ZN(N3857), .A1(N3843), .A2(N3852) );
  AND2_X1 AND2_1184( .ZN(N3858), .A1(N3852), .A2(N3840) );
  OR2_X1 OR2_1185( .ZN(N3859), .A1(N3857), .A2(N3858) );
  INV_X1 NOT1_1186( .ZN(N3864), .A(N3859) );
  AND2_X1 AND2_1187( .ZN(N3869), .A1(N3859), .A2(N3864) );
  OR2_X1 OR2_1188( .ZN(N3870), .A1(N3869), .A2(N3864) );
  INV_X1 NOT1_1189( .ZN(N3875), .A(N3870) );
  AND3_X1 AND3_1190( .ZN(N3876), .A1(N2826), .A2(N3028), .A3(N3870) );
  AND3_X1 AND3_1191( .ZN(N3877), .A1(N3826), .A2(N3876), .A3(N1591) );
  BUF_X1 BUFF1_1192( .Z(N3881), .A(N3877) );
  INV_X1 NOT1_1193( .ZN(N3882), .A(N3877) );
  BUF_X1 BUFF1_1194( .Z(N143_O), .A(N143_I) );
  BUF_X1 BUFF1_1195( .Z(N144_O), .A(N144_I) );
  BUF_X1 BUFF1_1196( .Z(N145_O), .A(N145_I) );
  BUF_X1 BUFF1_1197( .Z(N146_O), .A(N146_I) );
  BUF_X1 BUFF1_1198( .Z(N147_O), .A(N147_I) );
  BUF_X1 BUFF1_1199( .Z(N148_O), .A(N148_I) );
  BUF_X1 BUFF1_1200( .Z(N149_O), .A(N149_I) );
  BUF_X1 BUFF1_1201( .Z(N150_O), .A(N150_I) );
  BUF_X1 BUFF1_1202( .Z(N151_O), .A(N151_I) );
  BUF_X1 BUFF1_1203( .Z(N152_O), .A(N152_I) );
  BUF_X1 BUFF1_1204( .Z(N153_O), .A(N153_I) );
  BUF_X1 BUFF1_1205( .Z(N154_O), .A(N154_I) );
  BUF_X1 BUFF1_1206( .Z(N155_O), .A(N155_I) );
  BUF_X1 BUFF1_1207( .Z(N156_O), .A(N156_I) );
  BUF_X1 BUFF1_1208( .Z(N157_O), .A(N157_I) );
  BUF_X1 BUFF1_1209( .Z(N158_O), .A(N158_I) );
  BUF_X1 BUFF1_1210( .Z(N159_O), .A(N159_I) );
  BUF_X1 BUFF1_1211( .Z(N160_O), .A(N160_I) );
  BUF_X1 BUFF1_1212( .Z(N161_O), .A(N161_I) );
  BUF_X1 BUFF1_1213( .Z(N162_O), .A(N162_I) );
  BUF_X1 BUFF1_1214( .Z(N163_O), .A(N163_I) );
  BUF_X1 BUFF1_1215( .Z(N164_O), .A(N164_I) );
  BUF_X1 BUFF1_1216( .Z(N165_O), .A(N165_I) );
  BUF_X1 BUFF1_1217( .Z(N166_O), .A(N166_I) );
  BUF_X1 BUFF1_1218( .Z(N167_O), .A(N167_I) );
  BUF_X1 BUFF1_1219( .Z(N168_O), .A(N168_I) );
  BUF_X1 BUFF1_1220( .Z(N169_O), .A(N169_I) );
  BUF_X1 BUFF1_1221( .Z(N170_O), .A(N170_I) );
  BUF_X1 BUFF1_1222( .Z(N171_O), .A(N171_I) );
  BUF_X1 BUFF1_1223( .Z(N172_O), .A(N172_I) );
  BUF_X1 BUFF1_1224( .Z(N173_O), .A(N173_I) );
  BUF_X1 BUFF1_1225( .Z(N174_O), .A(N174_I) );
  BUF_X1 BUFF1_1226( .Z(N175_O), .A(N175_I) );
  BUF_X1 BUFF1_1227( .Z(N176_O), .A(N176_I) );
  BUF_X1 BUFF1_1228( .Z(N177_O), .A(N177_I) );
  BUF_X1 BUFF1_1229( .Z(N178_O), .A(N178_I) );
  BUF_X1 BUFF1_1230( .Z(N179_O), .A(N179_I) );
  BUF_X1 BUFF1_1231( .Z(N180_O), .A(N180_I) );
  BUF_X1 BUFF1_1232( .Z(N181_O), .A(N181_I) );
  BUF_X1 BUFF1_1233( .Z(N182_O), .A(N182_I) );
  BUF_X1 BUFF1_1234( .Z(N183_O), .A(N183_I) );
  BUF_X1 BUFF1_1235( .Z(N184_O), .A(N184_I) );
  BUF_X1 BUFF1_1236( .Z(N185_O), .A(N185_I) );
  BUF_X2 BUFF1_1237( .Z(N186_O), .A(N186_I) );
  BUF_X2 BUFF1_1238( .Z(N187_O), .A(N187_I) );
  BUF_X2 BUFF1_1239( .Z(N188_O), .A(N188_I) );
  BUF_X1 BUFF1_1240( .Z(N189_O), .A(N189_I) );
  BUF_X1 BUFF1_1241( .Z(N190_O), .A(N190_I) );
  BUF_X1 BUFF1_1242( .Z(N191_O), .A(N191_I) );
  BUF_X1 BUFF1_1243( .Z(N192_O), .A(N192_I) );
  BUF_X1 BUFF1_1244( .Z(N193_O), .A(N193_I) );
  BUF_X1 BUFF1_1245( .Z(N194_O), .A(N194_I) );
  BUF_X2 BUFF1_1246( .Z(N195_O), .A(N195_I) );
  BUF_X2 BUFF1_1247( .Z(N196_O), .A(N196_I) );
  BUF_X1 BUFF1_1248( .Z(N197_O), .A(N197_I) );
  BUF_X1 BUFF1_1249( .Z(N198_O), .A(N198_I) );
  BUF_X1 BUFF1_1250( .Z(N199_O), .A(N199_I) );
  BUF_X1 BUFF1_1251( .Z(N200_O), .A(N200_I) );
  BUF_X2 BUFF1_1252( .Z(N201_O), .A(N201_I) );
  BUF_X2 BUFF1_1253( .Z(N202_O), .A(N202_I) );
  BUF_X2 BUFF1_1254( .Z(N203_O), .A(N203_I) );
  BUF_X1 BUFF1_1255( .Z(N204_O), .A(N204_I) );
  BUF_X1 BUFF1_1256( .Z(N205_O), .A(N205_I) );
  BUF_X1 BUFF1_1257( .Z(N206_O), .A(N206_I) );
  BUF_X1 BUFF1_1258( .Z(N207_O), .A(N207_I) );
  BUF_X1 BUFF1_1259( .Z(N208_O), .A(N208_I) );
  BUF_X1 BUFF1_1260( .Z(N209_O), .A(N209_I) );
  BUF_X1 BUFF1_1261( .Z(N210_O), .A(N210_I) );
  BUF_X1 BUFF1_1262( .Z(N211_O), .A(N211_I) );
  BUF_X1 BUFF1_1263( .Z(N212_O), .A(N212_I) );
  BUF_X1 BUFF1_1264( .Z(N213_O), .A(N213_I) );
  BUF_X1 BUFF1_1265( .Z(N214_O), .A(N214_I) );
  BUF_X1 BUFF1_1266( .Z(N215_O), .A(N215_I) );
  BUF_X1 BUFF1_1267( .Z(N216_O), .A(N216_I) );
  BUF_X1 BUFF1_1268( .Z(N217_O), .A(N217_I) );
  BUF_X1 BUFF1_1269( .Z(N218_O), .A(N218_I) );

endmodule
