//# 28 inputs
//# 106 outputs
//# 1636 D-type flipflops
//# 13470 inverters
//# 8709 gates (4154 ANDs + 2050 NANDs + 226 ORs + 2279 NORs)

module s38417(CK,g1249,g16297,g16355,g16399,g16437,g16496,g1943,g24734,g25420,g25435,g25442,g25489,g26104,g26135,g26149,
  g2637,g27380,g3212,g3213,g3214,g3215,g3216,g3217,g3218,g3219,g3220,g3221,g3222,g3223,g3224,g3225,g3226,g3227,
  g3228,g3229,g3230,g3231,g3232,g3233,g3234,g3993,g4088,g4090,g4200,g4321,g4323,g4450,g4590,g51,g5388,g5437,
  g5472,g5511,g5549,g5555,g5595,g5612,g5629,g563,g5637,g5648,g5657,g5686,g5695,g5738,g5747,g5796,g6225,g6231,
  g6313,g6368,g6442,g6447,g6485,g6518,g6573,g6642,g6677,g6712,g6750,g6782,g6837,g6895,g6911,g6944,g6979,g7014,
  g7052,g7084,g7161,g7194,g7229,g7264,g7302,g7334,g7357,g7390,g7425,g7487,g7519,g7909,g7956,g7961,g8007,g8012,
  g8021,g8023,g8030,g8082,g8087,g8096,g8106,g8167,g8175,g8249,g8251,g8258,g8259,g8260,g8261,g8262,g8263,g8264,
  g8265,g8266,g8267,g8268,g8269,g8270,g8271,g8272,g8273,g8274,g8275);
input CK,g51,g563,g1249,g1943,g2637,g3212,g3213,g3214,g3215,g3216,g3217,g3218,g3219,g3220,g3221,g3222,g3223,
  g3224,g3225,g3226,g3227,g3228,g3229,g3230,g3231,g3232,g3233,g3234;
output g3993,g4088,g4090,g4200,g4321,g4323,g4450,g4590,g5388,g5437,g5472,g5511,g5549,g5555,g5595,g5612,g5629,g5637,g5648,g5657,
  g5686,g5695,g5738,g5747,g5796,g6225,g6231,g6313,g6368,g6442,g6447,g6485,g6518,g6573,g6642,g6677,g6712,g6750,g6782,g6837,
  g6895,g6911,g6944,g6979,g7014,g7052,g7084,g7161,g7194,g7229,g7264,g7302,g7334,g7357,g7390,g7425,g7487,g7519,g7909,g7956,
  g7961,g8007,g8012,g8021,g8023,g8030,g8082,g8087,g8096,g8106,g8167,g8175,g8249,g8251,g8258,g8259,g8260,g8261,g8262,g8263,
  g8264,g8265,g8266,g8267,g8268,g8269,g8270,g8271,g8272,g8273,g8274,g8275,g16297,g16355,g16399,g16437,g16496,g24734,g25420,g25435,
  g25442,g25489,g26104,g26135,g26149,g27380;

  wire g2814,g16475,g2817,g20571,g2933,g20588,g2950,g21951,g2883,g23315,g2888,g24423,g2896,g25175,g2892,g26019,
    g2903,g26747,g2900,g27237,g2908,g27715,g2912,g24424,g2917,g25174,g2924,g26020,g2920,g26746,g2984,g19061,
    g2985,g19060,g2930,g19062,g2929,g2879,g16494,g2934,g16476,g2935,g16477,g2938,g16478,g2941,g16479,g2944,
    g16480,g2947,g16481,g2953,g16482,g2956,g16483,g2959,g16484,g2962,g16485,g2963,g16486,g2966,g16487,g2969,
    g16488,g2972,g16489,g2975,g16490,g2978,g16491,g2981,g16492,g2874,g16493,g1506,g20572,g1501,g20573,g1496,
    g20574,g1491,g20575,g1486,g20576,g1481,g20577,g1476,g20578,g1471,g20579,g2877,g23313,g2861,g21960,g813,
    g2864,g21961,g809,g2867,g21962,g805,g2870,g21963,g801,g2818,g21947,g797,g2821,g21948,g793,g2824,
    g21949,g789,g2827,g21950,g785,g2830,g23312,g2873,g2833,g21952,g125,g2836,g21953,g121,g2839,g21954,
    g117,g2842,g21955,g113,g2845,g21956,g109,g2848,g21957,g105,g2851,g21958,g101,g2854,g21959,g97,
    g2858,g23316,g2857,g2200,g20587,g2195,g20585,g2190,g20586,g2185,g20584,g2180,g20583,g2175,g20582,g2170,
    g20581,g2165,g20580,g2878,g23314,g3129,g13475,g3117,g3109,g3210,g20630,g3211,g20631,g3084,g20632,g3085,
    g20609,g3086,g20610,g3087,g20611,g3091,g20612,g3092,g20613,g3093,g20614,g3094,g20615,g3095,g20616,g3096,
    g20617,g3097,g26751,g3098,g26752,g3099,g26753,g3100,g29163,g3101,g29164,g3102,g29165,g3103,g30120,g3104,
    g30121,g3105,g30122,g3106,g30941,g3107,g30942,g3108,g30943,g3155,g20618,g3158,g20619,g3161,g20620,g3164,
    g20621,g3167,g20622,g3170,g20623,g3173,g20624,g3176,g20625,g3179,g20626,g3182,g20627,g3185,g20628,g3088,
    g20629,g3191,g27717,g3194,g28316,g3197,g28317,g3198,g28318,g3201,g28704,g3204,g28705,g3207,g28706,g3188,
    g29463,g3133,g29656,g3132,g28698,g3128,g29166,g3127,g28697,g3126,g28315,g3125,g28696,g3124,g28314,g3123,
    g28313,g3120,g28695,g3114,g28694,g3113,g28693,g3112,g28312,g3110,g28311,g3111,g28310,g3139,g29461,g3136,
    g28701,g3134,g28700,g3135,g28699,g3151,g29462,g3142,g28703,g3147,g28702,g185,g29657,g138,g13405,g135,
    g165,g130,g24259,g131,g24260,g129,g24261,g133,g24262,g134,g24263,g132,g24264,g142,g24265,g143,
    g24266,g141,g24267,g145,g24268,g146,g24269,g144,g24270,g148,g24271,g149,g24272,g147,g24273,g151,
    g24274,g152,g24275,g150,g24276,g154,g24277,g155,g24278,g153,g24279,g157,g24280,g158,g24281,g156,
    g24282,g160,g24283,g161,g24284,g159,g24285,g163,g24286,g164,g24287,g162,g24288,g169,g26679,g170,
    g26680,g168,g26681,g172,g26682,g173,g26683,g171,g26684,g175,g26685,g176,g26686,g174,g26687,g178,
    g26688,g179,g26689,g177,g26690,g186,g30506,g189,g30507,g192,g30508,g231,g30842,g234,g30843,g237,
    g30844,g195,g30836,g198,g30837,g201,g30838,g240,g30845,g243,g30846,g246,g30847,g204,g30509,g207,
    g30510,g210,g30511,g249,g30515,g252,g30516,g255,g30517,g213,g30512,g216,g30513,g219,g30514,g258,
    g30518,g261,g30519,g264,g30520,g222,g30839,g225,g30840,g228,g30841,g267,g30848,g270,g30849,g273,
    g30850,g92,g25983,g88,g26678,g83,g27189,g79,g27683,g74,g28206,g70,g28673,g65,g29131,g61,
    g29413,g56,g29627,g52,g29794,g180,g20555,g182,g181,g276,g13406,g405,g401,g309,g11496,g354,
    g28207,g343,g28208,g346,g28209,g369,g28210,g358,g28211,g361,g28212,g384,g28213,g373,g28214,g376,
    g28215,g398,g28216,g388,g28217,g391,g28218,g408,g29414,g411,g29415,g414,g29416,g417,g29631,g420,
    g29632,g423,g29633,g427,g29417,g428,g29418,g426,g29419,g429,g27684,g432,g27685,g435,g27686,g438,
    g27687,g441,g27688,g444,g27689,g448,g28674,g449,g28675,g447,g28676,g312,g29795,g313,g29796,g314,
    g29797,g315,g30851,g316,g30852,g317,g30853,g318,g30710,g319,g30711,g320,g30712,g322,g29628,g323,
    g29629,g321,g29630,g403,g27191,g404,g27192,g402,g27193,g450,g11509,g451,g452,g11510,g453,g454,
    g11511,g279,g280,g11491,g281,g282,g11492,g283,g284,g11493,g285,g286,g11494,g287,g288,g11495,
    g289,g290,g13407,g291,g299,g19012,g305,g23148,g308,g23149,g297,g23150,g296,g23151,g295,g23152,
    g294,g23153,g304,g19016,g303,g19015,g302,g19014,g301,g19013,g300,g25130,g298,g27190,g342,g11497,
    g349,g350,g11498,g351,g352,g11499,g353,g357,g11500,g364,g365,g11501,g366,g367,g11502,g368,
    g372,g11503,g379,g380,g11504,g381,g382,g11505,g383,g387,g11506,g394,g395,g11507,g396,g397,
    g11508,g324,g325,g13408,g331,g337,g545,g13419,g551,g550,g554,g23160,g557,g20556,g510,g20557,
    g513,g16467,g523,g524,g564,g11512,g569,g570,g11515,g571,g572,g11516,g573,g574,g11517,g565,
    g566,g11513,g567,g568,g11514,g489,g474,g13409,g481,g485,g486,g24292,g487,g24293,g488,g24294,
    g455,g25139,g458,g25131,g461,g25132,g477,g25136,g478,g25137,g479,g25138,g480,g24289,g484,g24290,
    g464,g24291,g465,g25133,g468,g25134,g471,g25135,g528,g16468,g535,g542,g543,g19021,g544,g548,
    g23159,g549,g19022,g499,g558,g19023,g559,g576,g28219,g577,g28220,g575,g28221,g579,g28222,g580,
    g28223,g578,g28224,g582,g28225,g583,g28226,g581,g28227,g585,g28228,g586,g28229,g584,g28230,g587,
    g25985,g590,g25986,g593,g25987,g596,g25988,g599,g25989,g602,g25990,g614,g29135,g617,g29136,g620,
    g29137,g605,g29132,g608,g29133,g611,g29134,g490,g27194,g493,g27195,g496,g27196,g506,g8284,g507,
    g24295,g508,g19017,g509,g19018,g514,g19019,g515,g19020,g516,g23158,g517,g23157,g518,g23156,g519,
    g23155,g520,g23154,g525,g529,g13410,g530,g13411,g531,g13412,g532,g13413,g533,g13414,g534,g13415,
    g536,g13416,g537,g13417,g538,g25984,g541,g13418,g623,g13420,g626,g629,g630,g20558,g659,g21943,
    g640,g23161,g633,g24296,g653,g25140,g646,g25991,g660,g26691,g672,g27197,g666,g27690,g679,g28231,
    g686,g28677,g692,g29138,g699,g23162,g700,g23163,g698,g23164,g702,g23165,g703,g23166,g701,g23167,
    g705,g23168,g706,g23169,g704,g23170,g708,g23171,g709,g23172,g707,g23173,g711,g23174,g712,g23175,
    g710,g23176,g714,g23177,g715,g23178,g713,g23179,g717,g23180,g718,g23181,g716,g23182,g720,g23183,
    g721,g23184,g719,g23185,g723,g23186,g724,g23187,g722,g23188,g726,g23189,g727,g23190,g725,g23191,
    g729,g23192,g730,g23193,g728,g23194,g732,g23195,g733,g23196,g731,g23197,g735,g26692,g736,g26693,
    g734,g26694,g738,g24297,g739,g24298,g737,g24299,g826,g13421,g823,g853,g818,g24300,g819,g24301,
    g817,g24302,g821,g24303,g822,g24304,g820,g24305,g830,g24306,g831,g24307,g829,g24308,g833,g24309,
    g834,g24310,g832,g24311,g836,g24312,g837,g24313,g835,g24314,g839,g24315,g840,g24316,g838,g24317,
    g842,g24318,g843,g24319,g841,g24320,g845,g24321,g846,g24322,g844,g24323,g848,g24324,g849,g24325,
    g847,g24326,g851,g24327,g852,g24328,g850,g24329,g857,g26696,g858,g26697,g856,g26698,g860,g26699,
    g861,g26700,g859,g26701,g863,g26702,g864,g26703,g862,g26704,g866,g26705,g867,g26706,g865,g26707,
    g873,g30521,g876,g30522,g879,g30523,g918,g30860,g921,g30861,g924,g30862,g882,g30854,g885,g30855,
    g888,g30856,g927,g30863,g930,g30864,g933,g30865,g891,g30524,g894,g30525,g897,g30526,g936,g30530,
    g939,g30531,g942,g30532,g900,g30527,g903,g30528,g906,g30529,g945,g30533,g948,g30534,g951,g30535,
    g909,g30857,g912,g30858,g915,g30859,g954,g30866,g957,g30867,g960,g30868,g780,g25992,g776,g26695,
    g771,g27198,g767,g27691,g762,g28232,g758,g28678,g753,g29139,g749,g29420,g744,g29634,g740,g29798,
    g868,g20559,g870,g869,g963,g13422,g1092,g1088,g996,g11523,g1041,g28233,g1030,g28234,g1033,g28235,
    g1056,g28236,g1045,g28237,g1048,g28238,g1071,g28239,g1060,g28240,g1063,g28241,g1085,g28242,g1075,g28243,
    g1078,g28244,g1095,g29421,g1098,g29422,g1101,g29423,g1104,g29638,g1107,g29639,g1110,g29640,g1114,g29424,
    g1115,g29425,g1113,g29426,g1116,g27692,g1119,g27693,g1122,g27694,g1125,g27695,g1128,g27696,g1131,g27697,
    g1135,g28679,g1136,g28680,g1134,g28681,g999,g29799,g1000,g29800,g1001,g29801,g1002,g30869,g1003,g30870,
    g1004,g30871,g1005,g30713,g1006,g30714,g1007,g30715,g1009,g29635,g1010,g29636,g1008,g29637,g1090,g27206,
    g1091,g27207,g1089,g27208,g1137,g11536,g1138,g1139,g11537,g1140,g1141,g11538,g966,g967,g11518,g968,
    g969,g11519,g970,g971,g11520,g972,g973,g11521,g974,g975,g11522,g976,g977,g13423,g978,g986,
    g19024,g992,g27200,g995,g27201,g984,g27202,g983,g27203,g982,g27204,g981,g27205,g991,g19028,g990,
    g19027,g989,g19026,g988,g19025,g987,g25141,g985,g27199,g1029,g11524,g1036,g1037,g11525,g1038,g1039,
    g11526,g1040,g1044,g11527,g1051,g1052,g11528,g1053,g1054,g11529,g1055,g1059,g11530,g1066,g1067,g11531,
    g1068,g1069,g11532,g1070,g1074,g11533,g1081,g1082,g11534,g1083,g1084,g11535,g1011,g1012,g13424,g1018,
    g1024,g1231,g13435,g1237,g1236,g1240,g23198,g1243,g20560,g1196,g20561,g1199,g16469,g1209,g1210,g1250,
    g11539,g1255,g1256,g11542,g1257,g1258,g11543,g1259,g1260,g11544,g1251,g1252,g11540,g1253,g1254,g11541,
    g1176,g1161,g13425,g1168,g1172,g1173,g24333,g1174,g24334,g1175,g24335,g1142,g25150,g1145,g25142,g1148,
    g25143,g1164,g25147,g1165,g25148,g1166,g25149,g1167,g24330,g1171,g24331,g1151,g24332,g1152,g25144,g1155,
    g25145,g1158,g25146,g1214,g16470,g1221,g1228,g1229,g19033,g1230,g1234,g27217,g1235,g19034,g1186,g1244,
    g19035,g1245,g1262,g28245,g1263,g28246,g1261,g28247,g1265,g28248,g1266,g28249,g1264,g28250,g1268,g28251,
    g1269,g28252,g1267,g28253,g1271,g28254,g1272,g28255,g1270,g28256,g1273,g25994,g1276,g25995,g1279,g25996,
    g1282,g25997,g1285,g25998,g1288,g25999,g1300,g29143,g1303,g29144,g1306,g29145,g1291,g29140,g1294,g29141,
    g1297,g29142,g1177,g27209,g1180,g27210,g1183,g27211,g1192,g8293,g1193,g24336,g1194,g19029,g1195,g19030,
    g1200,g19031,g1201,g19032,g1202,g27216,g1203,g27215,g1204,g27214,g1205,g27213,g1206,g27212,g1211,g1215,
    g13426,g1216,g13427,g1217,g13428,g1218,g13429,g1219,g13430,g1220,g13431,g1222,g13432,g1223,g13433,g1224,
    g25993,g1227,g13434,g1309,g13436,g1312,g1315,g1316,g20562,g1345,g21944,g1326,g23199,g1319,g24337,g1339,
    g25151,g1332,g26000,g1346,g26708,g1358,g27218,g1352,g27698,g1365,g28257,g1372,g28682,g1378,g29146,g1385,
    g23200,g1386,g23201,g1384,g23202,g1388,g23203,g1389,g23204,g1387,g23205,g1391,g23206,g1392,g23207,g1390,
    g23208,g1394,g23209,g1395,g23210,g1393,g23211,g1397,g23212,g1398,g23213,g1396,g23214,g1400,g23215,g1401,
    g23216,g1399,g23217,g1403,g23218,g1404,g23219,g1402,g23220,g1406,g23221,g1407,g23222,g1405,g23223,g1409,
    g23224,g1410,g23225,g1408,g23226,g1412,g23227,g1413,g23228,g1411,g23229,g1415,g23230,g1416,g23231,g1414,
    g23232,g1418,g23233,g1419,g23234,g1417,g23235,g1421,g26709,g1422,g26710,g1420,g26711,g1424,g24338,g1425,
    g24339,g1423,g24340,g1520,g13437,g1517,g1547,g1512,g24341,g1513,g24342,g1511,g24343,g1515,g24344,g1516,
    g24345,g1514,g24346,g1524,g24347,g1525,g24348,g1523,g24349,g1527,g24350,g1528,g24351,g1526,g24352,g1530,
    g24353,g1531,g24354,g1529,g24355,g1533,g24356,g1534,g24357,g1532,g24358,g1536,g24359,g1537,g24360,g1535,
    g24361,g1539,g24362,g1540,g24363,g1538,g24364,g1542,g24365,g1543,g24366,g1541,g24367,g1545,g24368,g1546,
    g24369,g1544,g24370,g1551,g26713,g1552,g26714,g1550,g26715,g1554,g26716,g1555,g26717,g1553,g26718,g1557,
    g26719,g1558,g26720,g1556,g26721,g1560,g26722,g1561,g26723,g1559,g26724,g1567,g30536,g1570,g30537,g1573,
    g30538,g1612,g30878,g1615,g30879,g1618,g30880,g1576,g30872,g1579,g30873,g1582,g30874,g1621,g30881,g1624,
    g30882,g1627,g30883,g1585,g30539,g1588,g30540,g1591,g30541,g1630,g30545,g1633,g30546,g1636,g30547,g1594,
    g30542,g1597,g30543,g1600,g30544,g1639,g30548,g1642,g30549,g1645,g30550,g1603,g30875,g1606,g30876,g1609,
    g30877,g1648,g30884,g1651,g30885,g1654,g30886,g1466,g26001,g1462,g26712,g1457,g27219,g1453,g27699,g1448,
    g28258,g1444,g28683,g1439,g29147,g1435,g29427,g1430,g29641,g1426,g29802,g1562,g20563,g1564,g1563,g1657,
    g13438,g1786,g1782,g1690,g11550,g1735,g28259,g1724,g28260,g1727,g28261,g1750,g28262,g1739,g28263,g1742,
    g28264,g1765,g28265,g1754,g28266,g1757,g28267,g1779,g28268,g1769,g28269,g1772,g28270,g1789,g29434,g1792,
    g29435,g1795,g29436,g1798,g29645,g1801,g29646,g1804,g29647,g1808,g29437,g1809,g29438,g1807,g29439,g1810,
    g27700,g1813,g27701,g1816,g27702,g1819,g27703,g1822,g27704,g1825,g27705,g1829,g28684,g1830,g28685,g1828,
    g28686,g1693,g29803,g1694,g29804,g1695,g29805,g1696,g30887,g1697,g30888,g1698,g30889,g1699,g30716,g1700,
    g30717,g1701,g30718,g1703,g29642,g1704,g29643,g1702,g29644,g1784,g27221,g1785,g27222,g1783,g27223,g1831,
    g11563,g1832,g1833,g11564,g1834,g1835,g11565,g1660,g1661,g11545,g1662,g1663,g11546,g1664,g1665,g11547,
    g1666,g1667,g11548,g1668,g1669,g11549,g1670,g1671,g13439,g1672,g1680,g19036,g1686,g29428,g1689,g29429,
    g1678,g29430,g1677,g29431,g1676,g29432,g1675,g29433,g1685,g19040,g1684,g19039,g1683,g19038,g1682,g19037,
    g1681,g25152,g1679,g27220,g1723,g11551,g1730,g1731,g11552,g1732,g1733,g11553,g1734,g1738,g11554,g1745,
    g1746,g11555,g1747,g1748,g11556,g1749,g1753,g11557,g1760,g1761,g11558,g1762,g1763,g11559,g1764,g1768,
    g11560,g1775,g1776,g11561,g1777,g1778,g11562,g1705,g1706,g13440,g1712,g1718,g1925,g13451,g1931,g1930,
    g1934,g23236,g1937,g20564,g1890,g20565,g1893,g16471,g1903,g1904,g1944,g11566,g1949,g1950,g11569,g1951,
    g1952,g11570,g1953,g1954,g11571,g1945,g1946,g11567,g1947,g1948,g11568,g1870,g1855,g13441,g1862,g1866,
    g1867,g24374,g1868,g24375,g1869,g24376,g1836,g25161,g1839,g25153,g1842,g25154,g1858,g25158,g1859,g25159,
    g1860,g25160,g1861,g24371,g1865,g24372,g1845,g24373,g1846,g25155,g1849,g25156,g1852,g25157,g1908,g16472,
    g1915,g1922,g1923,g19045,g1924,g1928,g29445,g1929,g19046,g1880,g1938,g19047,g1939,g1956,g28271,g1957,
    g28272,g1955,g28273,g1959,g28274,g1960,g28275,g1958,g28276,g1962,g28277,g1963,g28278,g1961,g28279,g1965,
    g28280,g1966,g28281,g1964,g28282,g1967,g26003,g1970,g26004,g1973,g26005,g1976,g26006,g1979,g26007,g1982,
    g26008,g1994,g29151,g1997,g29152,g2000,g29153,g1985,g29148,g1988,g29149,g1991,g29150,g1871,g27224,g1874,
    g27225,g1877,g27226,g1886,g8302,g1887,g24377,g1888,g19041,g1889,g19042,g1894,g19043,g1895,g19044,g1896,
    g29444,g1897,g29443,g1898,g29442,g1899,g29441,g1900,g29440,g1905,g1909,g13442,g1910,g13443,g1911,g13444,
    g1912,g13445,g1913,g13446,g1914,g13447,g1916,g13448,g1917,g13449,g1918,g26002,g1921,g13450,g2003,g13452,
    g2006,g2009,g2010,g20566,g2039,g21945,g2020,g23237,g2013,g24378,g2033,g25162,g2026,g26009,g2040,g26725,
    g2052,g27227,g2046,g27706,g2059,g28283,g2066,g28687,g2072,g29154,g2079,g23238,g2080,g23239,g2078,g23240,
    g2082,g23241,g2083,g23242,g2081,g23243,g2085,g23244,g2086,g23245,g2084,g23246,g2088,g23247,g2089,g23248,
    g2087,g23249,g2091,g23250,g2092,g23251,g2090,g23252,g2094,g23253,g2095,g23254,g2093,g23255,g2097,g23256,
    g2098,g23257,g2096,g23258,g2100,g23259,g2101,g23260,g2099,g23261,g2103,g23262,g2104,g23263,g2102,g23264,
    g2106,g23265,g2107,g23266,g2105,g23267,g2109,g23268,g2110,g23269,g2108,g23270,g2112,g23271,g2113,g23272,
    g2111,g23273,g2115,g26726,g2116,g26727,g2114,g26728,g2118,g24379,g2119,g24380,g2117,g24381,g2214,g13453,
    g2211,g2241,g2206,g24382,g2207,g24383,g2205,g24384,g2209,g24385,g2210,g24386,g2208,g24387,g2218,g24388,
    g2219,g24389,g2217,g24390,g2221,g24391,g2222,g24392,g2220,g24393,g2224,g24394,g2225,g24395,g2223,g24396,
    g2227,g24397,g2228,g24398,g2226,g24399,g2230,g24400,g2231,g24401,g2229,g24402,g2233,g24403,g2234,g24404,
    g2232,g24405,g2236,g24406,g2237,g24407,g2235,g24408,g2239,g24409,g2240,g24410,g2238,g24411,g2245,g26730,
    g2246,g26731,g2244,g26732,g2248,g26733,g2249,g26734,g2247,g26735,g2251,g26736,g2252,g26737,g2250,g26738,
    g2254,g26739,g2255,g26740,g2253,g26741,g2261,g30551,g2264,g30552,g2267,g30553,g2306,g30896,g2309,g30897,
    g2312,g30898,g2270,g30890,g2273,g30891,g2276,g30892,g2315,g30899,g2318,g30900,g2321,g30901,g2279,g30554,
    g2282,g30555,g2285,g30556,g2324,g30560,g2327,g30561,g2330,g30562,g2288,g30557,g2291,g30558,g2294,g30559,
    g2333,g30563,g2336,g30564,g2339,g30565,g2297,g30893,g2300,g30894,g2303,g30895,g2342,g30902,g2345,g30903,
    g2348,g30904,g2160,g26010,g2156,g26729,g2151,g27228,g2147,g27707,g2142,g28284,g2138,g28688,g2133,g29155,
    g2129,g29446,g2124,g29648,g2120,g29806,g2256,g20567,g2258,g2257,g2351,g13454,g2480,g2476,g2384,g11577,
    g2429,g28285,g2418,g28286,g2421,g28287,g2444,g28288,g2433,g28289,g2436,g28290,g2459,g28291,g2448,g28292,
    g2451,g28293,g2473,g28294,g2463,g28295,g2466,g28296,g2483,g29447,g2486,g29448,g2489,g29449,g2492,g29652,
    g2495,g29653,g2498,g29654,g2502,g29450,g2503,g29451,g2501,g29452,g2504,g27708,g2507,g27709,g2510,g27710,
    g2513,g27711,g2516,g27712,g2519,g27713,g2523,g28689,g2524,g28690,g2522,g28691,g2387,g29807,g2388,g29808,
    g2389,g29809,g2390,g30905,g2391,g30906,g2392,g30907,g2393,g30719,g2394,g30720,g2395,g30721,g2397,g29649,
    g2398,g29650,g2396,g29651,g2478,g27230,g2479,g27231,g2477,g27232,g2525,g11590,g2526,g2527,g11591,g2528,
    g2529,g11592,g2354,g2355,g11572,g2356,g2357,g11573,g2358,g2359,g11574,g2360,g2361,g11575,g2362,g2363,
    g11576,g2364,g2365,g13455,g2366,g2374,g19048,g2380,g30314,g2383,g30315,g2372,g30316,g2371,g30317,g2370,
    g30318,g2369,g30319,g2379,g19052,g2378,g19051,g2377,g19050,g2376,g19049,g2375,g25163,g2373,g27229,g2417,
    g11578,g2424,g2425,g11579,g2426,g2427,g11580,g2428,g2432,g11581,g2439,g2440,g11582,g2441,g2442,g11583,
    g2443,g2447,g11584,g2454,g2455,g11585,g2456,g2457,g11586,g2458,g2462,g11587,g2469,g2470,g11588,g2471,
    g2472,g11589,g2399,g2400,g13456,g2406,g2412,g2619,g13467,g2625,g2624,g2628,g23274,g2631,g20568,g2584,
    g20569,g2587,g16473,g2597,g2598,g2638,g11593,g2643,g2644,g11596,g2645,g2646,g11597,g2647,g2648,g11598,
    g2639,g2640,g11594,g2641,g2642,g11595,g2564,g2549,g13457,g2556,g2560,g2561,g24415,g2562,g24416,g2563,
    g24417,g2530,g25172,g2533,g25164,g2536,g25165,g2552,g25169,g2553,g25170,g2554,g25171,g2555,g24412,g2559,
    g24413,g2539,g24414,g2540,g25166,g2543,g25167,g2546,g25168,g2602,g16474,g2609,g2616,g2617,g19057,g2618,
    g2622,g30325,g2623,g19058,g2574,g2632,g19059,g2633,g2650,g28297,g2651,g28298,g2649,g28299,g2653,g28300,
    g2654,g28301,g2652,g28302,g2656,g28303,g2657,g28304,g2655,g28305,g2659,g28306,g2660,g28307,g2658,g28308,
    g2661,g26012,g2664,g26013,g2667,g26014,g2670,g26015,g2673,g26016,g2676,g26017,g2688,g29159,g2691,g29160,
    g2694,g29161,g2679,g29156,g2682,g29157,g2685,g29158,g2565,g27233,g2568,g27234,g2571,g27235,g2580,g8311,
    g2581,g24418,g2582,g19053,g2583,g19054,g2588,g19055,g2589,g19056,g2590,g30324,g2591,g30323,g2592,g30322,
    g2593,g30321,g2594,g30320,g2599,g2603,g13458,g2604,g13459,g2605,g13460,g2606,g13461,g2607,g13462,g2608,
    g13463,g2610,g13464,g2611,g13465,g2612,g26011,g2615,g13466,g2697,g13468,g2700,g2703,g2704,g20570,g2733,
    g21946,g2714,g23275,g2707,g24419,g2727,g25173,g2720,g26018,g2734,g26742,g2746,g27236,g2740,g27714,g2753,
    g28309,g2760,g28692,g2766,g29162,g2773,g23276,g2774,g23277,g2772,g23278,g2776,g23279,g2777,g23280,g2775,
    g23281,g2779,g23282,g2780,g23283,g2778,g23284,g2782,g23285,g2783,g23286,g2781,g23287,g2785,g23288,g2786,
    g23289,g2784,g23290,g2788,g23291,g2789,g23292,g2787,g23293,g2791,g23294,g2792,g23295,g2790,g23296,g2794,
    g23297,g2795,g23298,g2793,g23299,g2797,g23300,g2798,g23301,g2796,g23302,g2800,g23303,g2801,g23304,g2799,
    g23305,g2803,g23306,g2804,g23307,g2802,g23308,g2806,g23309,g2807,g23310,g2805,g23311,g2809,g26743,g2810,
    g26744,g2808,g26745,g2812,g24420,g2813,g24421,g2811,g24422,g3054,g23317,g3079,g23318,g3080,g21965,g3043,
    g29453,g3044,g29454,g3045,g29455,g3046,g29456,g3047,g29457,g3048,g29458,g3049,g29459,g3050,g29460,g3051,
    g29655,g3052,g29972,g3053,g29973,g3055,g29974,g3056,g29975,g3057,g29976,g3058,g29977,g3059,g29978,g3060,
    g29979,g3061,g30119,g3062,g30908,g3063,g30909,g3064,g30910,g3065,g30911,g3066,g30912,g3067,g30913,g3068,
    g30914,g3069,g30915,g3070,g30940,g3071,g30980,g3072,g30981,g3073,g30982,g3074,g30983,g3075,g30984,g3076,
    g30985,g3077,g30986,g3078,g30987,g2997,g30989,g2993,g26748,g2998,g27238,g3006,g25177,g3002,g26021,g3013,
    g26750,g3010,g27239,g3024,g27716,g3018,g24425,g3028,g25176,g3036,g26022,g3032,g26749,g3040,g16497,g2986,
    g2987,g16495,g48,g20595,g45,g20596,g42,g20597,g39,g20598,g27,g20599,g30,g20600,g33,g20601,
    g36,g20602,g3083,g20603,g26,g20604,g2992,g21966,g23,g20605,g20,g20606,g17,g20607,g11,g20608,
    g14,g20589,g5,g20590,g8,g20591,g2,g20592,g2990,g20593,g2991,g21964,g1,g20594,II13089,g562,
    II13092,g1248,II13095,g1942,II13098,g2636,II13101,g3235,II13104,g3236,II13107,g3237,II13110,g3238,II13113,g3239,
    II13116,g3240,II13119,g3241,II13122,g3242,II13125,g3243,II13128,g3244,II13131,g3245,II13134,g3246,II13137,g3247,
    II13140,g3248,II13143,g3249,II13146,g3250,II13149,g3251,II13152,g3252,II13155,g3253,II13158,g3254,II13161,g3304,
    g3305,II13165,g3306,g3337,II13169,g3338,g3365,II13173,g3366,II13176,g3398,II13179,g3410,II13182,g3460,g3461,
    II13186,g3462,g3493,II13190,g3494,g3521,II13194,g3522,II13197,g3554,II13200,g3566,II13203,g3616,g3617,II13207,
    g3618,g3649,II13211,g3650,g3677,II13215,g3678,II13218,g3710,II13221,g3722,II13224,g3772,g3773,II13228,g3774,
    g3805,II13232,g3806,g3833,II13236,g3834,II13239,g3866,II13242,g3878,g3897,II13246,g3900,g3919,g3922,g3925,
    g3928,g3931,g3934,g3937,g3940,g3941,g3942,g3945,g3948,g3951,g3954,g3957,g3960,g3963,g3966,g3969,
    g3972,g3975,g3978,g3981,g3984,g3987,g3990,II13275,g3994,g3995,g3996,g3997,g3998,g3999,g4000,g4003,
    g4006,g4009,g4012,g4015,g4016,g4017,g4020,g4023,g4026,g4029,g4032,g4035,g4038,g4041,g4044,g4047,
    g4048,g4049,g4052,g4055,g4058,g4061,g4064,g4067,g4070,g4073,g4076,g4079,g4082,g4085,II13316,g4089,
    II13320,g4091,g4092,g4093,g4094,g4095,g4098,g4101,g4104,g4107,g4110,g4111,g4112,g4115,g4118,g4121,
    g4124,g4127,g4130,g4133,g4136,g4139,g4142,g4143,g4144,g4147,g4150,g4153,g4156,g4159,g4162,g4165,
    g4168,g4171,g4174,g4175,g4176,g4179,g4182,g4185,g4188,g4191,g4194,g4197,II13366,g4201,g4202,g4203,
    g4204,g4205,g4208,g4211,g4214,g4217,g4220,g4221,g4224,g4225,g4228,g4231,g4234,g4237,g4240,g4243,
    g4246,g4249,g4250,g4251,g4254,g4257,g4260,g4263,g4266,g4269,g4272,g4275,g4278,g4281,g4282,g4283,
    g4286,g4289,g4292,g4295,g4298,g4301,g4304,g4307,g4310,g4313,g4314,g4315,g4318,II13417,g4322,II13421,
    g4324,g4325,g4326,g4329,g4332,g4335,II13430,g4338,II13433,g4339,g4340,g4343,g4346,g4347,g4348,g4351,
    g4354,g4357,g4360,g4363,g4366,g4369,g4372,g4375,g4376,g4379,g4380,g4383,g4386,g4389,g4392,g4395,
    g4398,g4401,g4404,g4405,g4406,g4409,g4412,g4415,g4418,g4421,g4424,g4427,g4430,g4433,g4436,g4437,
    g4438,g4441,g4444,g4447,II13478,g4451,g4452,g4453,g4456,g4465,g4468,g4471,g4474,g4475,g4476,g4479,
    g4480,g4483,g4486,g4489,g4492,g4495,g4498,g4501,g4504,II13501,g4507,II13504,g4508,g4509,g4512,g4515,
    g4516,g4517,g4520,g4523,g4526,g4529,g4532,g4535,g4538,g4541,g4544,g4545,g4548,g4549,g4552,g4555,
    g4558,g4561,g4564,g4567,g4570,g4573,g4574,g4575,g4578,g4581,g4584,g4587,II13538,g4591,g4592,g4595,
    g4598,g4601,g4602,g4603,g4606,g4609,g4610,g4611,g4614,g4617,g4620,g4623,g4626,g4629,g4632,g4641,
    g4644,g4647,g4650,g4651,g4652,g4655,g4656,g4659,g4662,g4665,g4668,g4671,g4674,g4677,g4680,II13575,
    g4683,II13578,g4684,g4685,g4688,g4691,g4692,g4693,g4696,g4699,g4702,g4705,g4708,g4711,g4714,g4717,
    g4720,g4721,g4724,g4725,g4728,g4731,g4734,II13601,g4735,II13604,g4736,g4737,g4740,g4743,g4746,g4749,
    g4752,g4753,g4754,g4757,g4760,g4763,g4766,g4769,g4772,g4775,g4778,g4779,g4780,g4783,g4786,g4787,
    g4788,g4791,g4794,g4797,g4800,g4803,g4806,g4809,g4818,g4821,g4824,g4827,g4828,g4829,g4832,g4833,
    g4836,g4839,g4842,g4845,g4848,g4851,g4854,g4857,II13652,g4860,II13655,g4861,g4862,g4865,g4868,g4869,
    g4870,g4873,g4876,g4879,g4882,g4885,g4888,g4891,g4894,g4897,g4898,g4899,g4902,g4905,g4908,II13677,
    g4911,II13680,g4912,g4913,g4916,g4919,g4922,g4925,g4928,g4929,g4930,g4933,g4936,g4939,g4942,g4945,
    g4948,g4951,g4954,g4955,g4956,g4959,g4962,g4963,g4964,g4967,g4970,g4973,g4976,g4979,g4982,g4985,
    g4994,g4997,g5000,g5003,g5004,g5005,g5008,g5009,g5012,g5015,g5018,g5021,g5024,g5027,g5030,g5033,
    g5034,g5035,g5038,g5041,g5044,g5047,g5050,g5053,g5056,g5057,g5058,g5061,g5064,g5067,II13742,g5070,
    II13745,g5071,g5072,g5075,g5078,g5081,g5084,g5087,g5088,g5089,g5092,g5095,g5098,g5101,g5104,g5107,
    g5110,g5113,g5114,g5115,g5118,g5121,g5122,g5123,g5126,g5129,g5132,g5135,g5138,II13775,g5141,g5142,
    g5145,g5148,g5149,g5150,g5153,g5156,g5159,g5162,g5163,g5164,g5167,g5170,g5173,g5176,g5179,g5182,
    g5185,g5186,g5187,g5190,g5193,g5196,II13801,g5199,II13804,g5200,g5201,g5204,g5207,g5210,g5213,g5216,
    g5217,g5218,g5221,g5224,g5227,g5230,g5233,II13820,g5234,g5235,g5238,g5241,g5242,g5243,g5246,g5249,
    g5252,g5255,g5256,g5257,g5260,g5263,g5266,g5269,g5272,g5275,g5278,g5279,g5280,g5283,g5286,g5289,
    g5292,g5293,g5296,II13849,g5297,g5298,g5301,g5304,g5305,g5306,g5309,g5312,g5315,g5318,g5319,g5320,
    g5323,g5326,g5327,g5330,g5333,II13868,g5334,g5335,g5338,g5341,g5342,g5343,g5346,g5349,g5352,g5355,
    g5358,g5361,g5362,g5363,g5366,g5369,g5372,g5375,g5378,g5379,g5382,g5385,II13892,g5389,II13896,g5390,
    g5391,g5394,II13901,g5395,II13904,g5396,II13907,g5397,II13910,g5398,II13913,g5399,II13916,g5400,II13919,g5401,
    II13922,g5402,II13925,g5403,II13928,g5404,II13931,g5405,II13934,g5406,II13937,g5407,II13940,g5408,II13943,g5409,
    g5410,II13947,g5411,II13950,g5412,II13953,g5413,II13956,g5414,II13959,g5415,II13962,g5416,II13965,g5417,II13968,
    g5418,II13971,g5419,II13974,g5420,II13977,g5421,II13980,g5422,g5423,II13984,g5424,II13987,g5425,II13990,g5426,
    II13993,g5427,g5428,g5431,g5434,II13999,II14002,g5438,g5469,II14006,II14009,g5473,g5504,g5507,II14014,g5508,
    II14017,II14020,g5512,g5543,g5546,g5547,g5548,II14027,II14030,g5550,g5551,II14034,g5552,II14037,II14040,g5556,
    g5587,g5590,g5591,g5592,g5593,g5594,II14049,II14052,g5596,g5597,II14056,g5598,g5601,g5604,g5605,g5606,
    g5609,g5610,g5611,II14066,II14069,g5613,g5614,II14073,g5615,g5618,g5621,g5622,g5623,g5626,g5627,g5628,
    II14083,g5631,g5634,g5635,g5636,II14091,II14094,g5638,g5639,g5640,g5641,g5642,g5645,g5646,g5647,II14104,
    g5651,g5654,g5655,g5656,II14113,g5659,g5662,g5663,g5664,g5665,g5666,g5667,g5668,g5675,g5679,g5680,
    g5683,g5684,g5685,II14134,g5689,g5692,g5693,g5694,II14143,g5697,g5700,II14149,g5701,g5702,g5703,g5704,
    g5705,g5706,g5707,g5708,g5712,II14163,g5713,g5714,g5715,g5716,g5717,g5718,g5719,g5720,g5727,g5731,
    g5732,g5735,g5736,g5737,II14182,g5741,g5744,g5745,g5746,II14191,II14195,g5749,g5750,g5751,g5752,g5753,
    g5754,g5755,g5756,g5759,g5760,g5761,g5762,g5763,g5764,g5765,g5766,g5770,II14219,g5771,g5772,g5773,
    g5774,g5775,g5776,g5777,g5778,g5785,g5789,g5790,g5793,g5794,g5795,II14238,II14243,g5799,II14246,g5800,
    II14249,g5801,g5802,g5803,g5804,g5805,g5806,g5808,g5809,g5810,g5811,g5812,g5813,g5814,g5815,g5818,
    g5819,g5820,g5821,g5822,g5823,g5824,g5825,g5829,II14280,g5830,g5831,g5832,g5833,g5834,g5835,g5836,
    g5837,g5844,g5848,II14295,g5849,II14298,g5850,g5851,g5852,g5853,g5854,g5855,II14306,g5856,g5857,g5858,
    g5859,g5860,g5861,g5862,g5864,g5865,g5866,g5867,g5868,g5869,g5870,g5871,g5874,g5875,g5876,g5877,
    g5878,g5879,g5880,g5881,g5885,II14338,g5886,g5887,g5888,II14343,g5889,g5890,g5893,g5894,g5895,g5896,
    g5897,g5898,g5899,g5900,g5901,g5902,II14357,g5903,g5904,g5905,g5906,g5907,g5908,g5909,g5911,g5912,
    g5913,g5914,g5915,g5916,g5917,g5918,g5921,II14378,g5922,II14381,g5923,II14384,g5924,g5925,g5926,g5927,
    g5928,g5929,g5932,g5933,g5934,g5935,g5936,g5937,g5938,g5939,g5940,g5941,II14402,g5942,g5943,g5944,
    g5945,g5946,g5947,g5948,g5950,II14413,g5951,II14416,g5952,g5953,g5954,g5955,g5956,g5957,II14424,g5958,
    g5959,g5960,g5961,g5962,g5963,g5966,g5967,g5968,g5969,g5970,g5971,g5972,g5973,g5974,g5975,II14442,
    g5976,g5977,II14446,g5978,II14449,g5979,g5980,g5981,g5982,g5983,g5984,g5985,g5986,II14459,g5987,g5988,
    g5989,g5990,g5991,g5992,g5995,g5996,g5997,g5998,g5999,II14472,g6000,II14475,g6014,II14478,g6015,g6016,
    g6017,g6018,g6019,g6020,g6021,g6022,g6023,II14489,g6024,g6025,g6026,g6027,g6028,II14496,g6029,II14499,
    g6030,II14502,g6031,g6032,g6033,g6034,g6035,g6036,g6037,g6038,g6039,II14513,g6040,II14516,g6041,II14519,
    g6042,g6043,g6044,g6045,II14525,g6046,g6047,II14529,g6048,II14532,g6051,II14535,g6052,II14538,g6053,II14541,
    g6054,II14544,g6055,II14547,g6056,II14550,g6057,II14553,g6058,II14556,g6059,II14559,g6060,II14562,g6061,II14565,
    g6062,II14568,g6063,II14571,g6064,II14574,g6065,II14577,g6066,II14580,g6067,g6068,II14584,g6079,II14587,g6080,
    II14590,g6081,II14593,g6082,II14596,g6083,II14599,g6084,II14602,g6085,II14605,g6086,g6087,II14609,g6098,II14612,
    g6099,II14615,g6100,II14618,g6101,II14621,g6102,II14624,g6103,g6104,II14628,g6115,II14631,g6116,II14634,g6117,
    II14637,g6118,g6119,II14641,g6130,II14644,g6131,II14647,g6134,II14650,g6135,g6136,II14654,g6139,g6140,g6141,
    g6142,II14660,g6145,g6146,g6149,II14665,g6153,II14668,g6156,g6157,g6161,g6162,g6163,II14675,g6166,g6167,
    g6170,g6173,g6177,g6180,g6183,g6184,g6188,g6189,g6190,II14688,g6193,g6194,g6197,g6200,g6201,g6204,
    g6205,g6209,g6212,g6215,g6216,g6220,g6221,g6222,II14704,g6226,g6227,II14709,g6230,II14712,II14715,g6232,
    g6281,g6284,g6288,g6289,g6290,g6293,g6294,g6298,g6301,g6304,g6305,g6309,g6310,II14731,II14734,g6314,
    g6363,g6367,II14739,II14742,g6369,g6418,g6421,g6425,g6426,g6427,g6430,g6431,g6435,g6438,g6441,II14755,
    g6443,g6444,II14760,II14763,g6448,II14766,II14769,g6486,g6512,g6513,g6517,II14775,II14778,g6519,g6568,g6572,
    II14783,II14786,g6574,g6623,g6626,g6630,g6631,g6632,g6635,g6636,g6637,g6638,g6641,II14799,II14802,g6643,
    g6672,g6675,g6676,II14808,II14811,g6678,g6707,g6711,II14816,II14819,g6713,II14822,II14825,g6751,g6776,g6777,
    g6781,II14831,II14834,g6783,g6832,g6836,II14839,II14842,g6838,g6887,g6890,g6894,II14848,g6896,g6897,g6898,
    g6901,g6905,g6908,II14857,II14860,g6912,g6942,g6943,II14865,II14868,g6945,g6974,g6977,g6978,II14874,II14877,
    g6980,g7009,g7013,II14882,II14885,g7015,II14888,II14891,g7053,g7078,g7079,g7083,II14897,II14900,g7085,g7134,
    g7138,g7139,g7140,g7141,g7142,g7143,g7146,g7149,g7152,g7153,g7156,g7157,g7158,II14917,II14920,g7162,
    g7192,g7193,II14925,II14928,g7195,g7224,g7227,g7228,II14934,II14937,g7230,g7259,g7263,II14942,II14945,g7265,
    II14948,II14951,g7303,g7328,g7329,g7333,II14957,g7335,g7336,g7337,g7338,g7342,g7345,g7346,g7347,g7348,
    g7349,g7352,g7353,g7354,II14973,II14976,g7358,g7388,g7389,II14981,II14984,g7391,g7420,g7423,g7424,II14990,
    II14993,g7426,g7455,g7459,g7460,g7461,g7462,g7465,g7466,g7471,g7475,g7476,g7477,g7478,g7479,g7482,
    g7483,g7484,II15012,II15015,g7488,g7518,II15019,g7520,g7521,g7522,g7527,g7529,g7530,g7531,g7532,g7533,
    g7534,g7535,g7538,g7539,g7540,g7541,g7542,g7545,g7548,g7549,g7553,g7554,g7555,g7556,g7557,g7558,
    g7559,g7560,g7561,g7562,g7566,g7570,g7573,g7574,g7576,g7577,g7578,g7579,g7580,g7581,g7582,g7583,
    g7587,g7590,g7591,g7592,g7593,g7594,g7595,g7600,g7603,g7604,g7605,g7606,g7607,g7610,g7613,g7614,
    g7615,g7616,g7619,g7622,g7623,g7626,g7629,g7632,g7635,g7638,g7639,g7642,g7643,g7646,g7649,g7652,
    g7655,g7658,g7661,g7664,g7667,g7670,g7673,g7676,g7679,g7682,g7685,g7688,g7691,g7694,g7697,g7700,
    g7703,g7706,g7709,g7712,g7715,g7718,g7721,g7724,g7727,g7730,g7733,g7736,g7739,g7742,g7745,g7748,
    g7751,g7754,g7757,g7760,g7763,g7766,g7769,g7772,g7776,g7779,g7782,g7785,g7788,g7792,g7796,g7799,
    g7802,g7806,g7809,g7812,g7815,g7819,g7822,g7823,g7826,g7827,g7830,g7833,g7834,g7837,g7838,g7841,
    g7842,g7845,g7848,g7849,g7852,g7856,g7857,g7858,g7861,g7862,g7865,g7868,g7869,g7872,g7877,g7878,
    g7879,g7880,g7888,g7891,g7892,g7897,g7898,g7899,g7900,II15222,g7901,g7906,II15226,g7910,II15230,g7911,
    g7912,g7915,g7916,g7919,g7924,g7925,g7926,g7927,g7928,II15256,g7936,g7949,g7950,g7953,II15262,g7957,
    g7958,II15267,g7962,II15271,g7963,g7964,g7967,g7971,g7972,g7973,g7974,g7975,II15288,g7976,g7989,g7990,
    g7993,g7996,g7999,g8000,g8001,g8004,II15299,g8008,g8009,II15304,g8013,II15308,g8014,g8015,g8018,II15313,
    g8022,II15317,g8024,g8025,g8026,g8027,g8028,g8029,II15326,II15329,g8031,g8044,g8045,g8053,g8056,g8059,
    g8062,g8065,g8068,g8071,g8074,g8075,g8076,g8079,II15345,g8083,g8084,II15350,g8088,II15354,g8089,g8090,
    g8093,II15359,g8097,g8098,g8099,g8100,g8101,g8102,g8103,II15369,II15372,g8107,g8120,g8123,g8126,g8129,
    g8132,g8135,g8138,g8141,g8144,g8147,g8150,g8153,g8156,g8159,g8160,g8161,g8164,II15392,g8168,g8169,
    g8172,II15398,g8176,g8177,g8178,g8179,g8180,g8181,g8182,g8183,g8191,g8194,g8197,g8200,g8203,g8206,
    g8209,g8212,g8215,g8218,g8221,g8224,g8227,g8230,g8233,g8236,g8239,g8242,g8245,g8246,II15429,g8250,
    II15433,g8252,g8253,g8254,g8255,g8256,g8257,II15442,II15445,II15448,II15451,II15454,II15457,II15460,II15463,II15466,
    II15469,II15472,II15475,II15478,II15481,II15484,II15487,II15490,II15493,g8276,g8277,g8278,II15499,g8285,g8286,g8287,
    II15505,g8294,g8295,g8296,II15511,g8303,g8304,g8305,II15517,g8312,g8313,g8317,II15523,g8321,II15526,g8324,
    II15532,g8330,II15535,g8333,II15538,g8336,II15543,g8341,II15546,g8344,II15549,g8347,II15553,g8351,II15556,g8354,
    II15559,g8357,II15562,g8360,II15565,g8363,II15568,g8366,II15571,g8369,II15574,g8372,II15577,g8375,II15580,g8378,
    II15584,g8382,II15590,g8388,II15593,g8391,II15599,g8397,II15602,g8400,II15605,g8403,II15610,g8408,II15613,g8411,
    II15616,g8414,II15620,g8418,II15623,g8421,II15626,g8424,II15629,g8427,II15636,g8434,II15642,g8440,II15645,g8443,
    II15651,g8449,II15654,g8452,II15657,g8455,II15662,g8460,II15671,g8469,II15677,g8475,II15680,g8478,II15696,g8494,
    g8514,g8530,g8568,II15771,g8569,II15779,g8575,II15784,g8578,II15787,g8579,g8580,g8587,g8594,II15794,g8602,
    g8605,II15800,g8614,II15803,g8617,II15806,g8620,II15810,g8622,II15815,g8627,II15818,g8630,II15822,g8632,II15827,
    g8637,II15830,g8640,II15833,g8643,II15836,g8646,II15839,g8649,II15843,g8651,II15847,g8655,II15850,g8658,II15853,
    g8659,II15856,g8662,II15859,g8665,II15863,g8667,II15866,g8670,II15869,g8673,II15873,g8677,II15876,g8678,II15879,
    g8681,II15882,g8684,II15887,g8689,II15890,g8690,II15893,g8693,II15896,g8696,II15899,g8699,II15902,g8700,II15909,
    g8707,II15912,g8708,II15915,g8711,II15918,g8714,II15922,g8718,II15925,g8719,II15932,g8726,II15935,g8745,II15938,
    g8748,II15942,g8752,II15946,g8756,II15949,g8757,II15955,g8763,II15958,g8766,II15961,g8769,II15964,g8770,II15967,
    g8771,II15971,g8775,II15975,g8779,II15978,g8780,II15983,g8785,II15986,g8788,II15989,g8791,II15992,g8792,II15995,
    g8793,II15998,g8794,II16002,g8798,II16006,g8802,II16009,g8805,II16012,g8808,II16015,g8809,II16018,g8810,II16021,
    g8811,II16024,g8812,II16027,g8813,II16031,g8817,II16034,g8820,II16037,g8821,g8822,II16041,g8823,II16044,g8824,
    II16047,g8825,II16050,g8826,II16053,g8827,II16056,g8828,II16059,g8829,II16062,g8832,II16065,g8835,II16068,g8836,
    II16071,g8839,II16074,g8840,II16079,g8843,II16082,g8844,II16085,g8845,g8846,II16089,g8847,II16092,g8850,II16095,
    g8851,II16098,g8852,II16101,g8853,II16104,g8856,II16107,g8859,II16110,g8860,II16114,g8862,II16117,g8863,II16120,
    g8866,II16123,g8867,II16128,g8870,II16131,g8871,II16134,g8872,g8873,II16138,g8874,II16141,g8877,II16144,g8878,
    II16147,g8879,II16150,g8882,II16153,g8885,II16156,g8888,II16159,g8891,II16163,g8893,II16166,g8894,II16169,g8897,
    II16172,g8898,II16176,g8900,II16179,g8901,II16182,g8904,II16185,g8905,II16190,g8908,II16193,g8909,II16196,g8910,
    g8911,II16200,g8912,II16203,g8915,II16206,g8918,II16209,g8921,II16212,g8924,II16215,g8925,II16218,g8928,II16221,
    g8931,II16225,g8933,II16228,g8934,II16231,g8937,II16234,g8938,II16238,g8940,II16241,g8941,II16244,g8944,II16247,
    g8945,II16252,g8948,II16255,g8949,II16258,g8952,II16261,g8955,II16264,g8958,II16267,g8961,II16270,g8964,II16273,
    g8965,II16276,g8968,II16279,g8971,II16283,g8973,II16286,g8974,II16289,g8977,II16292,g8978,II16296,g8980,g8983,
    II16300,g8984,II16303,g8987,II16306,g8990,II16309,g8993,II16312,g8996,II16315,g8997,II16318,g9000,II16321,g9003,
    II16325,g9005,II16328,g9006,II16332,g9010,II16335,g9013,II16338,g9016,II16341,g9019,II16344,g9022,II16347,g9025,
    g9027,II16354,g9035,II16357,g9038,II16360,g9041,II16363,g9044,g9050,II16372,g9058,g9067,g9084,II16432,g9128,
    II16438,g9134,II16444,g9140,II16450,g9146,II16453,g9149,g9150,II16457,g9159,g9160,g9161,II16462,g9170,II16465,
    g9173,g9174,II16469,g9183,II16472,g9184,g9187,II16476,g9196,II16479,g9199,II16482,g9202,g9203,II16486,g9212,
    II16489,g9215,g9216,II16493,g9225,g9226,g9227,g9228,II16499,g9229,g9232,II16504,g9242,II16507,g9245,g9248,
    II16511,g9257,II16514,g9260,II16517,g9263,g9264,II16521,g9273,II16524,g9276,g9277,g9286,g9287,g9288,g9289,
    II16532,g9290,g9293,II16538,g9303,II16541,g9306,II16544,g9309,g9310,II16549,g9320,II16552,g9323,g9326,II16556,
    g9335,II16559,g9338,II16562,g9341,g9342,II16566,g9351,II16569,g9354,g9355,g9356,II16578,g9368,II16581,g9371,
    g9374,II16587,g9384,II16590,g9387,II16593,g9390,g9391,II16598,g9401,II16601,g9404,g9407,II16605,g9416,II16608,
    g9419,II16611,g9422,g9423,g9424,g9425,g9426,g9427,II16624,g9443,II16627,g9446,II16630,g9449,II16633,g9450,
    g9453,II16641,g9465,II16644,g9468,g9471,II16650,g9481,II16653,g9484,II16656,g9487,g9488,II16661,g9498,II16664,
    g9501,g9504,g9505,g9506,g9507,II16677,g9524,g9527,II16681,g9528,II16684,g9531,g9569,II16694,g9585,II16697,
    g9588,II16700,g9591,II16703,g9592,g9595,II16711,g9607,II16714,g9610,g9613,II16720,g9623,II16723,g9626,II16726,
    g9629,II16741,g9640,II16744,g9641,II16747,g9644,g9649,II16759,g9666,g9669,II16763,g9670,II16766,g9673,g9711,
    II16776,g9727,II16779,g9730,II16782,g9733,II16785,g9734,g9737,II16793,g9749,II16796,g9752,g9755,g9756,g9757,
    g9758,II16811,g9767,II16814,g9770,II16832,g9786,II16835,g9787,II16838,g9790,g9795,II16850,g9812,g9815,II16854,
    g9816,II16857,g9819,g9857,II16867,g9873,II16870,g9876,II16873,g9879,II16876,g9880,g9884,g9885,g9886,II16897,
    g9895,II16900,g9898,II16915,g9913,II16918,g9916,II16936,g9932,II16939,g9933,II16942,g9936,g9941,II16954,g9958,
    g9961,II16958,g9962,II16961,g9965,II16972,g10004,g10015,II16984,g10016,II16987,g10017,II16990,g10018,II16993,g10021,
    II17009,g10049,II17012,g10052,II17027,g10067,II17030,g10070,II17048,g10086,II17051,g10087,II17054,g10090,II17066,g10096,
    g10099,II17070,g7528,g10100,II17081,g10109,g10124,II17097,g10125,II17100,g10126,II17103,g10127,II17106,g10130,II17122,
    g10158,II17125,g10161,II17140,g10176,II17143,g10179,II17159,g10189,II17184,g10214,g10229,II17200,g10230,II17203,g10231,
    II17206,g10232,II17209,g10235,II17225,g10263,II17228,g10266,II17235,g10273,II17238,g10276,II17278,g10316,g10331,II17294,
    g10332,II17297,g10333,II17300,g10334,II17303,g10337,II17311,g10357,II17363,g10409,II17370,g10416,II17373,g10419,g10424,
    g10481,II17433,g10482,g10486,g10500,II17483,g10542,II17486,g10545,g10549,g10560,g10574,II17527,g10601,g10606,g10617,
    g10631,II17557,g10646,g10653,g10664,g10683,g10694,g10714,g10730,g10735,g10749,g10754,g10765,g10766,g10767,g10772,
    g10773,II17627,g7575,g10779,g10783,II17632,g10787,g10788,II17637,g10792,II17641,g10796,II17645,g10800,II17649,g10804,
    II17653,g10808,g10809,II17658,g10813,II17662,g10817,II17666,g10821,II17670,g10825,II17673,g10826,g10829,II17677,g10830,
    II17681,g10834,II17685,g10838,II17689,g10842,II17692,g10843,g10846,g10847,g10848,II17698,g10849,II17701,g10850,II17705,
    g10854,II17709,g10858,II17712,g10859,II17715,g10862,g10865,g10866,g10867,II17721,g10868,II17724,g10869,II17727,g10870,
    II17730,g10871,II17734,g10875,II17737,g10876,II17740,g10877,II17743,g10880,II17746,g10883,g10886,II17750,g10887,II17753,
    g10888,II17756,g10889,II17759,g10890,II17762,g10891,II17765,g10892,II17768,g10895,II17771,g10898,II17774,g10901,g10904,
    g10905,g10906,II17780,g10907,II17783,g10908,II17786,g10909,II17789,g10910,II17792,g10911,II17795,g10912,II17798,g10915,
    II17801,g10918,II17804,g10921,II17807,g10924,g10927,g10928,g10929,II17813,g10930,II17816,g10931,II17819,g10932,II17822,
    g10933,II17825,g10934,II17828,g10935,II17831,g10936,II17834,g10937,II17837,g10940,II17840,g10943,II17843,g10946,II17846,
    g10949,II17849,g10952,g10961,g10962,II17854,g10963,II17857,g10966,II17860,g10967,II17863,g10968,II17866,g10969,II17869,
    g10972,II17872,g10973,II17875,g10974,II17878,g10977,II17881,g10980,II17884,g10983,g10986,g10987,II17889,g10988,II17892,
    g10991,II17895,g10994,II17898,g10995,II17901,g10996,II17904,g10999,II17907,g11002,II17910,g11003,II17913,g11004,II17916,
    g11007,II17919,g11008,II17922,g11011,II17925,g11014,II17928,g11017,g11020,g11021,II17933,g11022,II17936,g11025,II17939,
    g11028,II17942,g11031,II17945,g11032,II17948,g11035,II17951,g11036,II17954,g11039,II17957,g11042,II17960,g11045,II17963,
    g11048,II17966,g11051,II17969,g11054,II17972,g11055,II17975,g11056,II17978,g7795,g11059,II17981,g11063,II17984,g11066,
    g11069,g11078,II17989,g11079,II17992,g11082,II17995,g11085,II17998,g11088,II18001,g11091,II18004,g11092,II18007,g11095,
    II18010,g11098,II18013,g11101,II18016,g11102,II18019,g11105,II18022,g11108,II18025,g11111,II18028,g11114,II18031,g11117,
    II18034,g11120,II18037,g11123,II18040,g11126,II18043,g11129,II18046,g11132,II18049,g11135,II18052,g11138,II18055,g11141,
    II18058,g11144,II18061,g11145,II18064,g11148,II18067,g11151,II18070,g11154,II18073,g11157,II18076,g11160,II18079,g11163,
    II18082,g11166,II18085,g11169,II18088,g11170,II18091,g11173,II18094,g11176,II18097,g11179,II18100,g11182,II18103,g11185,
    g11190,II18121,g11199,II18124,g11202,II18127,g11205,II18130,g11208,II18133,g11209,II18136,g11210,II18139,g11213,II18142,
    g11216,II18145,g11219,II18148,g11222,II18151,g11225,II18154,g11228,II18157,g11231,II18160,g11234,II18163,g11237,II18166,
    g11240,II18169,g11243,II18172,g11246,II18175,g11249,II18178,g11252,II18181,g11255,II18184,g11256,II18187,g11259,II18211,
    g11265,II18214,g11268,II18217,g11271,II18220,g11274,II18223,g11277,II18226,g11278,II18229,g11281,II18232,g11284,II18235,
    g11287,II18238,g11290,II18241,g11291,II18244,g11294,II18247,g11297,II18250,g11300,II18253,g11303,II18256,g11306,II18259,
    g11309,II18262,g11312,II18265,g11315,II18268,g11318,II18271,g11321,II18274,g11324,II18277,g11327,g11332,II18295,g11341,
    II18298,g11344,II18302,g11348,II18305,g11351,II18308,g11354,II18311,g11355,II18314,g11358,II18317,g11361,II18320,g11364,
    II18323,g11367,II18326,g11370,II18329,g11373,II18332,g11376,II18335,g11379,II18338,g11382,II18341,g11385,II18344,g11386,
    II18347,g11389,II18350,g11392,II18353,g11395,II18356,g11398,II18359,g11401,II18362,g11404,II18365,g11407,II18375,g11411,
    II18378,g11414,II18381,g11417,II18386,g11422,II18389,g11425,II18392,g11428,II18396,g11432,II18399,g11435,II18402,g11438,
    II18405,g11441,II18408,g11444,II18411,g11447,II18414,g11450,II18417,g11453,II18420,g11456,II18423,g11459,II18426,g11462,
    II18429,g11465,II18432,g11468,II18435,g11471,II18438,g11472,II18441,g11475,II18444,g11478,g11481,g11490,II18449,II18452,
    II18455,II18458,II18461,II18464,II18467,II18470,II18473,II18476,II18479,II18482,II18485,II18488,II18491,II18494,II18497,II18500,
    II18503,II18506,II18509,II18512,II18515,II18518,II18521,II18524,II18527,II18530,II18533,II18536,II18539,II18542,II18545,II18548,
    II18551,II18554,II18557,II18560,II18563,II18566,II18569,II18572,II18575,II18578,II18581,II18584,II18587,II18590,II18593,II18596,
    II18599,II18602,II18605,II18608,II18611,II18614,II18617,II18620,II18623,II18626,II18629,II18632,II18635,II18638,II18641,II18644,
    II18647,II18650,II18653,II18656,II18659,II18662,II18665,II18668,II18671,II18674,II18677,II18680,II18683,II18686,II18689,II18692,
    II18695,II18698,II18701,II18704,II18707,II18710,II18713,II18716,II18719,II18722,II18725,II18728,II18731,II18734,II18737,II18740,
    II18743,II18746,II18749,II18752,II18755,II18758,II18761,II18764,II18767,II18770,II18773,g11599,II18777,g11603,II18780,g11606,
    II18784,g11608,II18787,g11611,II18791,g11613,II18794,g11616,g11620,g11623,II18810,g11628,II18813,g11629,II18817,g11633,
    II18820,g11636,II18824,g11638,II18827,g11641,g11642,II18835,g11651,II18838,g11652,II18842,g11656,II18845,g11659,II18854,
    g11670,II18857,g11671,II18866,g11682,g11706,g11732,g11734,g11735,g11736,g11737,g11740,g11741,g11742,g11743,g11745,
    g11746,g11747,g11748,II18929,g10711,g11749,g11758,g11761,g11762,g11763,g11764,g11765,g11766,II18943,g11769,g11770,
    g11774,g11775,g11776,g11777,g11778,g11779,g11782,g11783,II18962,g11786,g11787,II18969,g11791,g11794,g11795,g11796,
    g11797,g11798,g11801,g11802,g11803,g11804,g11808,g11809,II18990,g11812,g11813,g11817,g11818,g11819,g11820,g11821,
    g11824,g11825,g11826,g11827,g11829,g11834,g11835,g11836,g11837,g11841,g11842,II19025,g11845,g11846,II19030,g11848,
    g11852,g11853,g11854,g11856,g11857,g11858,g11859,g11862,g11866,g11867,g11868,g11869,g11871,g11876,g11877,g11878,
    g11879,g11883,g11884,g11886,g11887,g11888,g11891,g11892,g11893,g11894,g11895,g11898,g11899,g11900,g11901,g11904,
    g11908,g11909,g11910,g11911,g11913,g11918,g11919,g11920,g11921,II19105,g11923,g11927,g11929,g11930,g11931,g11932,
    g11933,g11936,II19119,g11937,g11941,g11942,g11943,g11944,g11945,g11948,g11949,g11950,g11951,g11954,g11958,g11959,
    g11960,g11961,g11963,g11968,g11969,g11970,g11971,g11972,g11973,II19160,g11976,g11982,g11983,g11984,g11985,g11986,
    g11989,II19174,g11990,g11994,g11995,g11996,g11997,g11998,g12001,g12002,g12003,g12004,g12007,II19195,g12009,g12013,
    g12017,g12020,g12021,g12022,g12023,g12024,g12025,II19208,g12027,II19211,g12030,g12037,g12038,g12039,g12040,g12041,
    g12042,II19226,g12045,g12051,g12052,g12053,g12054,g12055,g12058,II19240,g12059,g12063,g12064,g12065,g12066,g12067,
    g12071,g12075,g12076,g12077,g12078,g12084,g12085,g12086,g12087,g12088,g12089,II19271,g12091,II19274,g12094,g12101,
    g12102,g12103,g12104,g12105,g12106,II19289,g12109,g12115,g12116,g12117,g12118,g12119,g12122,II19303,g12123,II19307,
    g12125,g12130,g12134,g12135,II19315,g12136,II19318,g12139,II19321,g12142,g12147,g12148,g12149,g12150,g12156,g12157,
    g12158,g12159,g12160,g12161,II19342,g12163,II19345,g12166,g12173,g12174,g12175,g12176,g12177,g12178,II19360,g12181,
    g12187,g12191,g12196,g12197,II19374,g12198,II19377,g12201,II19380,g12204,g12209,g12210,g12211,g12212,g12218,g12219,
    g12220,g12221,g12222,g12223,II19401,g12225,II19404,g12228,g12235,II19412,g12239,II19415,g12242,g12246,g12251,g12252,
    II19426,g12253,II19429,g12256,II19432,g12259,g12264,g12265,g12266,g12267,g12275,II19449,g12279,II19452,g12282,II19455,
    g12285,g12289,g12294,g12295,II19466,g12296,II19469,g12299,II19472,g12302,g12308,II19479,g12312,II19482,g12315,II19485,
    g12318,II19488,g12321,g12325,g12332,II19500,g12333,II19503,g12336,II19507,g12340,II19510,g12343,II19513,g12346,II19516,
    g12349,g12354,g8381,g12362,II19523,g12363,II19526,g12366,II19530,g12370,II19533,g12373,g12378,II19539,g12379,II19542,
    g12382,II19545,g12385,II19549,g12389,II19552,g8430,g12392,g12408,II19557,g12409,II19560,g12412,II19563,g12415,g12420,
    II19569,g12421,g12424,II19573,g12425,II19576,g12426,g12430,II19582,g12432,g12434,II19587,g12435,II19591,g12437,g12438,
    II19595,g10810,g12439,II19598,g12440,II19602,g12442,II19605,g10797,g12443,II19608,g10831,g12444,II19611,g12445,II19615,
    g10789,g12447,II19618,g10814,g12448,II19621,g10851,g12449,II19624,g12450,II19628,g10784,g12452,II19631,g10801,g12453,
    II19634,g10835,g12454,II19637,g10872,g12455,g12456,II19642,g10793,g12460,II19645,g10818,g12461,II19648,g10855,g12462,
    g12463,g12466,II19654,g10805,g12470,II19657,g10839,g12471,g12472,g12473,g12476,g12478,g12481,II19667,g10822,g12485,
    g12490,g12493,g12495,g12498,g12502,g12504,g12505,g12510,g12513,g12515,g12518,II19689,g12519,g12521,g12522,g12527,
    g12530,g12532,g12533,II19702,g12534,g12536,g12537,g12542,II19711,g12543,g12545,g12546,g12547,II19718,g12548,g12551,
    II19722,g12552,g12553,g12554,II19727,g12555,g12558,g12559,g12560,II19733,g12561,II19736,g12564,II19739,g12565,g12596,
    g12597,g12598,g12599,g12600,II19747,g12601,II19750,g12604,II19753,g12607,II19756,g12608,II19759,g12611,g12642,g12643,
    g12644,g12645,g12646,II19767,g12647,II19771,g10038,g12651,II19774,g12654,II19777,g12657,g12688,g12689,g12690,g12691,
    II19784,g12692,II19787,g12695,II19791,g12699,II19794,g10676,g12702,II19797,g10147,g12705,II19800,g12708,II19803,g12711,
    g12742,g12743,II19808,g12744,g12748,II19813,g10649,g12749,II19816,g10703,g12752,II19820,g12756,II19823,g10705,g12759,
    II19826,g10252,g12762,II19829,g12765,g12768,II19833,g12769,II19836,g12772,g12775,g12776,g12782,II19844,g8533,g12783,
    II19847,g10677,g12786,g12790,II19852,g10679,g12791,II19855,g10723,g12794,II19859,g12798,II19862,g10725,g12801,II19865,
    g10354,g12804,g12807,II19869,g12808,II19872,g12811,g12815,II19877,g8547,g12816,g12821,II19883,g8550,g12822,II19886,
    g10706,g12825,g12829,II19891,g10708,g12830,II19894,g10744,g12833,II19898,g12837,II19901,g10746,g12840,g12843,II19905,
    g12844,g12847,g12848,g12850,g12851,g12853,II19915,g8560,g12854,g12859,II19921,g8563,g12860,II19924,g10726,g12863,
    g12867,II19929,g10728,g12868,II19932,g10763,g12871,g12874,g12875,g12881,g12882,g12891,g12892,g12894,II19952,g8571,
    g12895,g12900,II19958,g8574,g12901,II19961,g10747,g12904,g12907,g12909,g12914,g12915,g12921,g12922,g12931,g12932,
    g12934,II19986,g8577,g12935,g12940,g12943,g12944,g12950,g12951,g12960,g12961,II20009,g12962,g12965,g12969,g12972,
    g12973,g12979,g12980,g12993,g12996,g12997,g12998,g13003,II20062,g10480,g13011,g13025,g13033,g13036,g13043,g13046,
    g13049,g13057,g13060,g13063,g13066,II20117,g13070,g13073,g13076,g13079,g13092,g13095,g13101,g13107,g13117,g13130,
    g13141,g13148,g13151,g13152,g13153,g13154,g13157,g13158,g13159,g13161,g13162,g13163,g13166,g13167,g13168,g13169,
    g13170,g13172,g13173,g13174,g13176,g13177,g13178,g13179,g13180,g13181,g13183,g13184,g13185,g13186,g13187,g13188,
    g13189,g13190,g13191,g13192,g13193,g13195,g13196,g13197,g13198,g13199,g13200,g13201,g13202,g13203,g13204,g13205,
    g13206,g13207,g13208,g13209,g13210,g13211,g13212,g13213,g13214,II20264,g13215,g13218,g13219,g13220,g13221,g13222,
    g13223,g13224,g13225,g13226,g13227,II20278,g13229,g13232,g13233,II20283,g13234,g13237,g13238,g13239,g13240,g13241,
    g13242,g13243,g13244,II20295,g13246,II20299,g13248,g13249,g13250,II20305,g13252,g13255,g13256,II20310,g13257,g13260,
    g13261,g13262,g13263,g13264,g13265,II20320,g13267,g13268,II20324,g13269,II20328,g13271,g13272,g13273,II20334,g13275,
    g13278,g13279,II20339,g13280,g13283,g13284,g13285,II20347,g13290,II20351,g13292,g13293,II20355,g13294,II20359,g13296,
    g13297,g13298,II20365,g13300,g13303,g13304,g13308,g13309,II20376,g13317,II20379,g13318,II20382,g13319,II20386,g13321,
    II20390,g13323,g13324,II20394,g13325,II20398,g13327,g13328,g13329,g13330,II20407,g13336,II20410,g13339,II20414,g13341,
    II20417,g13342,II20421,g13344,II20425,g13346,g13347,g13351,g13352,II20441,g13356,II20444,g13359,II20448,g13361,II20451,
    g13364,II20455,g13366,II20458,g13367,II20462,g13369,g13373,II20476,g13381,II20479,g13384,II20483,g13386,II20486,g13389,
    II20490,g13391,II20493,g13394,II20497,g13396,II20500,g13397,g13398,g13400,II20514,II20517,II20520,II20523,II20526,II20529,
    II20532,II20535,II20538,II20541,II20544,II20547,II20550,II20553,II20556,II20559,II20562,II20565,II20568,II20571,II20574,II20577,
    II20580,II20583,II20586,II20589,II20592,II20595,II20598,II20601,II20604,II20607,II20610,II20613,II20616,II20619,II20622,II20625,
    II20628,II20631,II20634,II20637,II20640,II20643,II20646,II20649,II20652,II20655,II20658,II20661,II20664,II20667,II20670,II20673,
    II20676,II20679,II20682,II20685,II20688,II20691,II20694,II20697,II20700,II20703,II20706,g13469,II20709,g13519,g13228,g13530,
    g13251,g13541,g13274,g13552,g13299,g13565,g12192,g13568,g11627,II20791,g13149,g13571,II20794,g13111,g13572,g13573,
    g12247,g13576,g11650,II20799,g13155,g13579,II20802,g13160,g13580,II20805,g13124,g13581,g13582,g12290,g13585,g11669,
    II20810,g13164,g13588,II20813,g13589,II20816,g12487,g13598,II20820,g13171,g13600,II20823,g13135,g13601,g13602,g12326,
    g13605,g11681,II20828,g13175,g13608,II20832,g12507,g13610,II20836,g13182,g13612,II20839,g13143,g13613,g13614,g11690,
    II20844,g12524,g13620,II20848,g13194,g13622,II20852,g12457,g13624,g13626,g11697,II20858,g12539,g13632,II20863,g12467,
    g13635,g13637,g11703,g13644,II20873,g12482,g13647,g13649,g11711,g13657,g13669,g13670,II20886,g12499,g13673,g13677,
    g13687,g13699,g13700,g13706,g13714,g13724,g13736,g13737,II20909,g13055,g13741,g13750,g13756,g13764,g13774,g13786,
    g13791,g13797,g13805,g13817,g13819,g13825,g13836,g13838,g13840,g13848,g11744,g13849,g13850,g13852,g13856,g11759,
    g13857,g11760,g13858,g13859,g13861,II20959,g11713,g13863,g13864,g11767,g13866,g11772,g13867,g11773,g13868,g13869,
    g13872,g11780,g13873,g12698,g13879,g11784,g13881,g11789,g13882,g11790,g13883,g13885,g11799,g13886,g12747,g13894,
    g11806,g13895,g12755,g13901,g11810,g13903,g11815,g13906,g11822,g13907,g12781,g13918,g11830,g13922,g11831,g13926,
    g11832,g13927,g12789,g13935,g11839,g13936,g12797,g13942,g11843,g13945,g11855,g13946,g12814,II21012,g12503,g13954,
    g13958,g11863,g13962,g11864,g13963,g12820,g13974,g11872,g13978,g11873,g13982,g11874,g13983,g12828,g13991,g11881,
    g13992,g12836,g13999,g11889,g14000,g11890,g14001,g12849,II21037,g12486,g14008,g14011,g11896,g14015,g11897,g14016,
    g12852,II21045,g12520,g14024,g14028,g11905,g14032,g11906,g14033,g12858,g14044,g11914,g14048,g11915,g14052,g11916,
    g14053,g12866,g14061,g11928,g14062,g12880,II21064,g13147,g14068,g14071,g11934,g14079,g11935,g14086,g11938,g14090,
    g11939,g14091,g11940,g14092,g12890,II21075,g12506,g14099,g14102,g11946,g14106,g11947,g14107,g12893,II21083,g12535,
    g14115,g14119,g11955,g14123,g11956,g14124,g12899,g14135,g11964,g14139,g11965,II21096,g14144,g14148,g12912,g14153,
    g12913,g14158,g11974,g14165,g11975,g14171,g11979,g14175,g11980,g14176,g11981,g14177,g12920,II21108,g13150,g14183,
    g14186,g11987,g14194,g11988,g14201,g11991,g14205,g11992,g14206,g11993,g14207,g12930,II21119,g12523,g14214,g14217,
    g11999,g14221,g12000,g14222,g12933,II21127,g12544,g14230,g14234,g12008,g14238,g12939,g14244,g12026,g14249,g12034,
    g14252,g12035,g14256,g12036,II21137,g14259,g14263,g12941,g14268,g12942,g14273,g12043,g14280,g12044,g14286,g12048,
    g14290,g12049,g14291,g12050,g14292,g12949,II21149,g13156,g14298,g14301,g12056,g14309,g12057,g14316,g12060,g14320,
    g12061,g14321,g12062,g14322,g12959,II21160,g12538,g14329,g14332,g12068,II21165,g13110,g14337,g14342,g12967,g14347,
    g12079,g14352,g12081,g14355,g12082,g14359,g12083,g14360,g12968,g14366,g12090,g14371,g12098,g14374,g12099,g14378,
    g12100,II21178,g14381,g14385,g12970,g14390,g12971,g14395,g12107,g14402,g12108,g14408,g12112,g14412,g12113,g14413,
    g12114,g14414,g12978,II21190,g13165,g14420,g14423,g12120,g14431,g12121,g14438,g12124,g14442,g11768,g14450,g12146,
    g14454,g12991,g14459,g12151,g14464,g12153,g14467,g12154,g14471,g12155,g14472,g12992,g14478,g12162,g14483,g12170,
    g14486,g12171,g14490,g12172,II21208,g14493,g14497,g12994,g14502,g12995,g14507,g12179,g14514,g12180,g14520,g12184,
    g14524,g12185,g14525,g12195,g14529,g11785,g14537,g12208,g14541,g13001,g14546,g12213,g14551,g12215,g14554,g12216,
    g14558,g12217,g14559,g13002,g14565,g12224,g14570,g12232,g14573,g12233,g14577,g12234,g14580,g12250,g14584,g11811,
    g14592,g12263,g14596,g13022,g14601,g12268,g14606,g12270,g14609,g12271,g14613,g12272,g14614,g12293,g14618,g11844,
    g14626,g12306,II21241,g13378,g14630,g14637,g12329,g14641,g11823,II21246,g11624,g14642,II21249,g11600,g14650,II21252,
    g11644,g14657,g14668,g11865,II21256,g11647,g14669,II21259,g11630,g14677,II21262,g14684,g14685,g12245,II21267,g11663,
    g14691,g14702,g11907,II21271,g11666,g14703,II21274,g11653,g14711,II21277,g14718,g14719,g12288,II21282,g11675,g14725,
    g14736,g11957,II21286,g11678,g14737,II21289,g14745,II21292,g14746,g14747,g12324,II21297,g11687,g14753,g14764,II21301,
    g14765,II21304,g14766,g14768,g12352,II21310,g14774,II21313,g14775,g14776,g12033,g14794,II21318,g14795,II21321,g14796,
    g14797,g12080,g14811,g12097,II21326,g14829,II21329,g14830,g14831,g11828,g14837,g12145,g14849,g12152,g14863,g12169,
    g14881,II21337,g14882,II21340,g14883,g14885,g11860,g14895,g12193,g14904,g11870,g14910,g12207,g14922,g12214,g14936,
    g12231,II21351,g14954,II21354,g14955,g14959,II21361,g13026,g14960,II21364,g13028,g14963,g14966,g11902,g14976,g12248,
    g14985,g11912,g14991,g12262,g15003,g12269,g15017,II21374,g15018,II21377,g15019,II21381,g15021,g15022,g11781,g15032,
    g15033,II21389,g12883,g15034,II21392,g13020,g15037,II21395,g13034,g15040,II21398,g13021,g15043,g15048,II21404,g13037,
    g15049,II21407,g13039,g15052,g15055,g11952,g15065,g12291,g15074,g11962,g15080,g12305,II21415,g15092,II21420,g15095,
    g15096,g11800,II21426,g11661,g15106,II21429,g13027,g15109,II21432,g13044,g15112,II21435,g11662,g15115,g15118,g11807,
    g15128,g15129,II21443,g12923,g15130,II21446,g13029,g15133,II21449,g13047,g15136,II21452,g13030,g15139,g15144,II21458,
    g13050,g15145,II21461,g13052,g15148,g15151,g12005,g15161,g12327,g15170,g15174,g15175,g15176,g15177,g12339,II21476,
    g11672,g15179,II21479,g13035,g15182,II21482,g13058,g15185,g15188,g11833,II21488,g11673,g15198,II21491,g13038,g15201,
    II21494,g13061,g15204,II21497,g11674,g15207,g15210,g11840,g15220,g15221,II21505,g12952,g15222,II21508,g13040,g15225,
    II21511,g13064,g15228,II21514,g13041,g15231,g15236,II21520,g13067,g15237,II21523,g13069,g15240,II21531,g11683,g15248,
    II21534,g13045,g15251,II21537,g13071,g15254,g15260,g15261,g15262,g15263,g12369,II21548,g11684,g15265,II21551,g13048,
    g15268,II21554,g13074,g15271,g15274,g11875,II21560,g11685,g15284,II21563,g13051,g15287,II21566,g13077,g15290,II21569,
    g11686,g15293,g15296,g11882,g15306,g15307,II21577,g12981,g15308,II21580,g13053,g15311,II21583,g13080,g15314,II21586,
    g13054,g15317,g15322,g15323,II21595,g11691,g15326,II21598,g13059,g15329,II21601,g13087,g15332,II21609,g11692,g15340,
    II21612,g13062,g15343,II21615,g13090,g15346,g15352,g15353,g15354,g15355,g12388,II21626,g11693,g15357,II21629,g13065,
    g15360,II21632,g13093,g15363,g15366,g11917,II21638,g11694,g15376,II21641,g13068,g15379,II21644,g13096,g15382,II21647,
    g11695,g15385,g15390,II21655,g11696,g15393,II21658,g13072,g15396,II21661,g13098,g15399,II21666,g13100,g15404,g15408,
    g15409,II21674,g11698,g15412,II21677,g13075,g15415,II21680,g13102,g15418,II21688,g11699,g15426,II21691,g13078,g15429,
    II21694,g13105,g15432,g15438,g15439,g15440,g15441,g12418,II21705,g11700,g15443,II21708,g13081,g15446,II21711,g13108,
    g15449,g15458,II21720,g11701,g15461,II21723,g13088,g15464,II21726,g13112,g15467,II21730,g13089,g15471,g15474,II21736,
    g11702,g15477,II21739,g13091,g15480,II21742,g13114,g15483,II21747,g13116,g15488,g15492,g15493,II21755,g11704,g15496,
    II21758,g13094,g15499,II21761,g13118,g15502,II21769,g11705,g15510,II21772,g13097,g15513,II21775,g13121,g15516,II21780,
    g13305,g15521,g15524,g15525,II21787,g11707,g15528,II21790,g13099,g15531,II21793,g13123,g15534,II21796,g11708,g15537,
    g15544,II21803,g11709,g15547,II21806,g13103,g15550,II21809,g13125,g15553,II21813,g13104,g15557,g15560,II21819,g11710,
    g15563,II21822,g13106,g15566,II21825,g13127,g15569,II21830,g13129,g15574,g15578,g15579,II21838,g11712,g15582,II21841,
    g13109,g15585,II21844,g13131,g15588,II21852,g11716,g15596,II21855,g13113,g15599,g15602,g15603,II21862,g11717,g15606,
    II21865,g13115,g15609,II21868,g13134,g15612,II21871,g11718,g15615,g15622,II21878,g11719,g15625,II21881,g13119,g15628,
    II21884,g13136,g15631,II21888,g13120,g15635,g15638,II21894,g11720,g15641,II21897,g13122,g15644,II21900,g13138,g15647,
    II21905,g13140,g15652,II21908,g13082,g15655,g15659,g15665,II21918,g11721,g15667,II21923,g11722,g15672,II21926,g13126,
    g15675,g15678,g15679,II21933,g11723,g15682,II21936,g13128,g15685,II21939,g13142,g15688,II21942,g11724,g15691,g15698,
    II21949,g11725,g15701,II21952,g13132,g15704,II21955,g13144,g15707,II21959,g13133,g15711,II21962,g13004,g15714,g15722,
    g15724,II21974,g11726,g15726,II21979,g11727,g15731,II21982,g13137,g15734,g15737,g15738,II21989,g11728,g15741,II21992,
    g13139,g15744,II21995,g13146,g15747,II21998,g11729,g15750,g15762,g15764,II22014,g11730,g15766,II22019,g11731,g15771,
    II22022,g13145,g15774,II22025,g11617,g15777,g15790,g15792,II22044,g11733,g15794,g15800,g15813,g15859,II22120,g15876,
    g15880,g15890,g15904,g15913,g15923,g15933,g15942,g15952,g15962,g15971,g15981,II22163,g12433,g15989,g15991,g15994,
    g15997,g16001,g16002,g16005,g16007,g16011,g16012,g16013,g16014,g16023,g16024,g16025,g16026,g16027,g16034,g16035,
    g16039,g16040,g16041,g16042,g16043,g16044,g16054,g16055,g16056,g16057,g16061,g16062,g16063,g16064,g16065,g16075,
    g11861,g16088,g16090,g16091,g16092,g16093,g16097,g16098,g16099,g16113,g11903,g16126,g16128,g16129,g16130,g16131,
    g16142,g16154,g12194,g16164,g11953,g16177,g16179,g16180,g16189,g16201,g16213,g12249,g16223,g12006,g16236,g16243,
    g16254,g16266,g16278,g12292,g16287,g16293,II22382,g16302,g16313,g16325,g16337,g12328,g16351,II22414,g16360,g16371,
    g16395,II22444,g16404,g16433,II22475,g16466,II22503,II22506,II22509,II22512,II22515,II22518,II22521,II22524,II22527,II22530,
    II22533,II22536,II22539,II22542,II22545,II22548,II22551,II22554,II22557,II22560,II22563,II22566,II22569,II22572,II22575,II22578,
    II22581,II22584,II22587,II22590,II22593,g16501,II22599,g16506,g16507,II22604,g16514,g16515,g16523,II22611,g16528,g16529,
    II22618,g16540,g16543,g16546,g16554,II22626,g16559,g16560,II22640,g16572,g16575,g16578,g16586,II22651,g16596,g16599,
    g16602,II22657,g16608,II22663,g16616,g16619,II22667,g16622,II22671,g16626,II22676,g16633,II22679,g16636,II22683,g16640,
    II22687,g16644,II22690,g16647,II22694,g16651,II22699,g16656,II22702,g16659,g16665,II22715,g16673,II22718,g16676,g16682,
    g16686,II22726,g16694,g16697,II22730,g16702,g16708,g16712,II22737,g16719,g16722,II22741,g16725,g16728,II22745,g16733,
    g16739,g16743,g16749,g15782,II22752,g16758,II22755,g16761,g16764,II22759,g16767,g16770,II22763,g16775,g16781,II22768,
    g16785,II22771,g16788,g16791,II22775,g16794,g16797,g16804,g15803,g16809,g15842,II22783,g16813,II22786,g16814,II22789,
    g16817,g16820,g16825,g15855,II22797,g16830,II22800,g16831,II22803,g16832,g16836,g15818,g16840,g15878,II22810,g16842,
    II22813,g16843,g16846,g15903,II22820,g16848,II22823,g16849,II22828,g16852,II22836,g16858,II22842,g16862,II22845,g16863,
    g16867,II22852,g16877,II22855,g16878,II22860,g16881,g16884,g16895,II22866,g16905,II22869,g16906,II22875,g16910,g16913,
    g16924,II22881,g16934,II22893,g16940,g16943,g16954,II22912,g16971,g16974,g17029,g17057,g17063,g17092,g17098,g17130,
    g17136,g17157,II23253,g17189,II23274,g17200,g17203,II23287,g17207,g17208,II23292,g17212,g17214,g17217,II23309,g16132,
    g17227,II23314,g15720,g17230,II23317,g16181,g17233,II23323,g15664,g17237,II23326,g15758,g17240,II23329,g15760,g17243,
    II23335,g16412,g17249,II23338,g15721,g17252,II23341,g15784,g17255,g17258,g16053,II23345,g15723,g17259,II23348,g15786,
    g17262,II23351,g15788,g17265,II23358,g16442,g17272,II23361,g15759,g17275,II23364,g15805,g17278,g17281,g16081,II23368,
    g16446,g17282,II23371,g15761,g17285,II23374,g15807,g17288,II23377,g15763,g17291,II23380,g15809,g17294,II23383,g15811,
    g17297,II23386,g17300,II23392,g13476,g17304,II23395,g15785,g17307,II23398,g15820,g17310,g17313,g16109,g17314,g16110,
    II23403,g13478,g17315,II23406,g15787,g17318,II23409,g15822,g17321,II23412,g13482,g17324,II23415,g15789,g17327,II23418,
    g15824,g17330,II23421,g15791,g17333,II23424,g15826,g17336,II23430,g13494,g17342,II23433,g15806,g17345,II23436,g15832,
    g17348,g17351,g16152,II23442,g13495,g17354,II23445,g15808,g17357,II23448,g15834,g17360,II23451,g13497,g17363,II23454,
    g15810,g17366,II23457,g15836,g17369,II23460,g13501,g17372,II23463,g15812,g17375,II23466,g15838,g17378,II23472,g13510,
    g17384,II23475,g15821,g17387,II23478,g15844,g17390,g17394,g16197,II23487,g13511,g17399,II23490,g15823,g17402,II23493,
    g15846,g17405,II23498,g13512,g17410,II23501,g15825,g17413,II23504,g15848,g17416,II23507,g13514,g17419,II23510,g15827,
    g17422,II23513,g15850,g17425,II23518,g15856,g17430,II23521,g13518,g17433,II23524,g15833,g17436,II23527,g15858,g17439,
    II23530,g17442,g17445,g16250,II23539,g13524,g17451,II23542,g15835,g17454,II23545,g15867,g17457,II23553,g13525,g17465,
    II23556,g15837,g17468,II23559,g15869,g17471,II23564,g13526,g17476,II23567,g15839,g17479,II23570,g15871,g17482,II23575,
    g15843,g17487,II23578,g15879,g17490,II23581,g13528,g17493,II23584,g15845,g17496,g17499,g16292,II23588,g17500,II23591,
    g17503,II23599,g15887,g17511,II23602,g13529,g17514,II23605,g15847,g17517,II23608,g15889,g17520,II23611,g17523,II23619,
    g13535,g17531,II23622,g15849,g17534,II23625,g15898,g17537,II23633,g13536,g17545,II23636,g15851,g17548,II23639,g15900,
    g17551,II23645,g13537,g17557,II23648,g15857,g17560,II23651,g13538,g17563,g17566,g16346,II23655,g17567,II23658,g17570,
    II23661,g16085,g17573,II23667,g15866,g17579,II23670,g15912,g17582,II23673,g13539,g17585,II23676,g15868,g17588,II23679,
    g17591,II23682,g17594,II23689,g15920,g17601,II23692,g13540,g17604,II23695,g15870,g17607,II23698,g15922,g17610,II23701,
    g17613,II23709,g13546,g17621,II23712,g15872,g17624,II23715,g15931,g17627,II23725,g13547,g17637,g17640,II23729,g17645,
    g17648,g16384,II23733,g17649,II23739,g13548,g17655,II23742,g15888,g17658,II23745,g13549,g17661,II23748,g17664,II23751,
    g17667,II23754,g16123,g17670,II23760,g15897,g17676,II23763,g15941,g17679,II23766,g13550,g17682,II23769,g15899,g17685,
    II23772,g17688,II23775,g17691,II23782,g15949,g17698,II23785,g13551,g17701,II23788,g15901,g17704,II23791,g15951,g17707,
    II23794,g17710,g17720,g15853,g17724,II23817,g13557,g17738,g17741,II23821,g17746,II23824,g17749,II23830,g13558,g17755,
    II23833,g15921,g17758,II23836,g13559,g17761,II23839,g17764,II23842,g17767,II23845,g16174,g17770,II23851,g15930,g17776,
    II23854,g15970,g17779,II23857,g13560,g17782,II23860,g15932,g17785,II23863,g17788,II23866,g17791,II23874,g15797,g17799,
    g17802,II23888,g17815,g17825,II23904,g13561,g17839,g17842,II23908,g17847,II23911,g17850,II23917,g13562,g17856,II23920,
    g15950,g17859,II23923,g13563,g17862,II23926,g17865,II23929,g17868,II23932,g16233,g17871,g17878,g15830,g17882,g17892,
    g17893,II23954,g17903,g17914,II23976,g17927,g17937,II23992,g13564,g17951,g17954,II23996,g17959,II23999,g17962,g17969,
    g15841,g17974,g17984,g17988,g17991,g17993,g18003,g18004,II24049,g18014,g18025,II24071,g18038,g18048,g18063,g15660,
    g18070,g15854,g18074,g18084,g18089,g18091,g18101,g18105,g18108,g18110,g18120,g18121,II24144,g18131,g18142,II24166,
    g18155,II24171,g16439,g18166,g18170,g15877,g18174,g18179,g18188,g18190,g18200,g18205,g18207,g18217,g18221,g18224,
    g18226,g18236,g18237,II24247,g18247,II24258,g16463,g18258,g18261,g15719,g18265,g18275,II24285,g15992,g18278,g18281,
    g18286,g18295,g18297,g18307,g18312,g18314,g18324,g18328,g18331,II24346,g15873,g18334,g18337,g15757,g18341,g18351,
    g18353,II24368,g15990,g18355,g18358,g18368,II24394,g15995,g18371,g18374,g18379,g18388,g18390,g18400,g18405,g18407,
    g15959,g18414,g15718,g18415,g15783,g18429,II24459,g13599,g18432,g18435,g18436,g18446,g18448,II24481,g15993,g18450,
    g18453,g18463,II24507,g15999,g18466,g18469,g18474,g18483,g18485,g15756,g18486,g15804,g18490,g18502,II24560,g13611,
    g18505,g18508,g18509,g18519,g18521,II24582,g15996,g18523,g18526,g18536,II24608,g16006,g18539,g18543,g15819,g18552,
    g18554,g18566,II24662,g13621,g18569,g18572,g18573,g18583,g18585,II24684,g16000,g18587,g18593,g15831,g18602,g18604,
    g18616,II24732,g13633,g18619,g18622,g18634,g18636,g18643,g18646,g16341,g18656,g18670,g18679,g18691,g18692,g18699,
    g18708,g18720,g18725,g13865,g18727,g18728,g18735,g18744,g18756,g18757,g18758,g18764,g18765,g18772,g18783,g18784,
    g18785,g18786,g18787,g18788,g18789,g18795,g18796,g18805,g18806,g18807,g18808,g18809,g18810,g18811,g18812,g18813,
    g18814,g18815,g18822,g18823,g18824,g18825,g18826,g18827,g18828,g18829,g18830,g18831,g18832,g18833,g18834,g18838,
    g18839,g18840,g18841,g18842,g18843,g18844,g18845,g18846,g18847,g18848,g18849,g18850,g18851,g18853,g18854,g18855,
    g18856,g18857,g18858,g18859,g18860,g18861,g18862,g18863,g18864,g18865,II24894,g18869,g18870,g18871,g18872,g18873,
    g18874,g18875,g18876,g18877,g18878,g18879,g18880,g18881,g18882,g18884,II24913,g18886,II24916,g18890,g18891,g18892,
    g18893,g18894,II24923,g18895,g18896,g18897,g18898,g18899,g18900,g18901,g18902,g18903,g18904,g18905,g18908,g18909,
    g18910,g18911,g18912,II24943,g18913,g18914,g18915,g18916,g18917,II24950,g18918,g18919,g18920,g18921,g18922,g18923,
    g18924,g18925,g18926,g18927,g18928,g18929,g18930,g18931,II24966,g18932,g18933,g18934,g18935,g18936,II24973,g18937,
    g18938,g18939,g18940,g18941,g18943,II24982,g18944,g18945,g18946,g18947,g18948,g18949,g18950,g18951,II24992,g18952,
    g18953,g18954,g18955,g18956,g18958,II25001,g18959,II25004,g18960,g18961,g18962,g18963,g18964,g18965,g18966,g18967,
    II25015,g18969,II25018,g18970,II25021,g18971,g18972,g18973,g18974,g18976,II25037,g18981,II25041,g18983,II25044,g18984,
    II25047,g18985,II25050,g18986,g18987,II25054,g18988,II25057,g18989,II25061,g18991,II25064,g18992,II25067,g18993,II25071,
    g18995,II25074,g18996,II25078,g18998,II25081,g18999,II25084,g19000,g19001,II25089,g19008,II25092,g19009,II25096,g19011,
    II25099,II25102,II25105,II25108,II25111,II25114,II25117,II25120,II25123,II25126,II25129,II25132,II25135,II25138,II25141,II25144,
    II25147,II25150,II25153,II25156,II25159,II25162,II25165,II25168,II25171,II25174,II25177,II25180,II25183,II25186,II25189,II25192,
    II25195,II25198,II25201,II25204,II25207,II25210,II25213,II25216,II25219,II25222,II25225,II25228,II25231,II25234,II25237,II25240,
    II25243,II25246,II25249,II25253,g17124,g19064,g19070,II25258,g19075,g19078,II25264,g17151,g19081,II25272,g17051,g19091,
    g19096,g18980,II25283,g17086,g19098,II25294,g19105,II25303,g19110,II25308,g19113,II25315,g19118,II25320,g19125,II25325,
    g19132,II25334,g19145,II25338,g19147,II25344,g19151,II25351,g19156,II25355,g18669,g19158,II25358,g18678,g19159,II25365,
    g18707,g19164,II25371,g18719,g19168,II25374,g18726,g19169,II25377,g18743,g19170,II25383,g18755,g19174,II25386,g18763,
    g19175,II25389,g18780,g19176,II25395,g18782,g19180,II25399,g18794,g19182,II25402,g18821,g19183,II25406,g18804,g19185,
    II25412,g18820,g19189,II25415,g18835,g19190,II25423,g18852,g19196,II25426,g18836,g19197,II25429,g18975,g19198,II25432,
    g18837,g19199,II25442,g18866,g19207,II25445,g18968,g19208,II25456,g18883,g19217,II25459,g18867,g19218,II25463,g18868,
    g19220,II25474,g18885,g19229,II25486,g18754,g19237,II25489,g18906,g19238,II25492,g18907,g19239,II25506,g18781,g19247,
    II25510,g18542,g19249,g19251,II25525,g18803,g19258,II25528,g18942,g19259,g19265,II25557,g18957,g19270,II25567,g17186,
    g19272,g19280,g19287,II25612,g17197,g19291,g19299,g19301,g19302,g17025,g19305,II25660,g17204,g19309,g19319,g19322,
    g19323,g17059,g19326,II25717,g17209,g19330,II25728,g17118,g19335,g19346,g19349,g19350,g17094,g19353,II25768,g17139,
    g19358,II25778,g17145,g19369,g19380,g19383,g19384,g17132,g19387,g16567,g19388,II25816,g17162,g19390,II25826,g17168,
    g19401,g19412,g19415,g19417,g16591,g19418,II25862,g17177,g19420,II25872,g17183,g19431,g19441,g17213,g19444,g17985,
    g19448,g19452,g19454,g16611,g19455,II25904,g17194,g19457,g19467,g19468,g17216,g19471,g18102,g19475,g19479,g19481,
    g16629,g19482,g19483,g19484,g19490,g19491,g17219,g19494,g18218,g19498,g19502,g19504,g19505,g19511,g19512,g17221,
    g19515,g18325,g19519,g19523,g19524,g19530,g19533,g19534,II25966,g16654,g19543,II25971,g16671,g19546,II25977,g16692,
    g19550,II25985,g16718,g19556,II25994,g16860,g19563,II26006,g16866,g19573,g19577,g19578,II26025,g16803,g19595,II26028,
    g16566,g19596,g19607,g19608,II26051,g16824,g19622,g19640,g19641,II26078,g16835,g19652,II26085,g18085,g19657,g19680,
    g19681,II26112,g16844,g19689,II26115,g16845,g19690,II26123,g19696,II26134,g18201,g19705,II26154,g16851,g19725,II26171,
    g19740,II26182,g18308,g19749,II26195,g16853,g19762,II26198,g16854,g19763,II26220,g19783,II26231,g18401,g19792,II26237,
    g16857,g19798,II26266,g19825,g19830,II26276,g16861,g19838,II26334,g18977,g19890,II26337,g16880,g19893,II26340,g19894,
    II26365,g18626,g19915,g19918,II26369,g19919,g19933,g18548,II26388,g19934,II26401,g17012,g19945,g19948,g17896,g19950,
    g18598,II26407,g19951,II26413,g16643,g19957,II26420,g17042,g19972,g19975,g18007,g19977,g18630,II26426,g16536,g19978,
    II26437,g16655,g19987,II26444,g17076,g20002,g20005,g18124,g20007,g18639,II26458,g20016,II26469,g16672,g20025,II26476,
    g17111,g20040,g20043,g18240,II26481,g18590,g20045,II26494,g20058,II26505,g16693,g20067,II26512,g16802,g20082,g20083,
    g17968,II26535,g20099,II26545,g16823,g20105,II26574,g20124,g20127,g18623,g20140,g20163,g17973,II26612,g20164,g20178,
    g20193,II26642,g20198,g20212,g20223,II26664,g20228,g20242,g20250,II26679,g20255,g20269,g20273,g20278,g20279,g20281,
    g20286,g20287,g20288,g20289,g20290,g20292,II26714,g20295,g20296,g20297,g20298,g20302,g20303,g20304,g20305,g20306,
    g20308,g20311,g20312,g20313,g20315,g20316,g20317,g20321,g20322,g20323,g20324,g20325,g20327,g20328,g20329,g20330,
    g20331,g20332,g20334,g20335,g20336,g20340,g20341,g20342,g20344,g20345,g20346,g20347,g20348,g20349,g20350,g20351,
    g20352,g20354,g20355,g20356,II26777,g17222,g20360,g20361,g20362,g20363,g20364,g20365,g20366,g20367,g20368,g20369,
    g20370,g20371,g20372,g20373,g20374,II26796,g17224,g20377,g20378,g20379,g20380,g20381,g20382,g20383,g20384,g20385,
    g20386,g20387,g20388,g20389,g20390,g20391,g20392,g20393,g20394,II26816,g17225,g20395,II26819,g17226,g20396,g20397,
    g20398,g20399,g20400,g20401,g20402,g20403,g20404,g20405,g20406,g20407,g20408,g20409,g20410,g20411,g20412,g20413,
    g20414,g20415,g20416,II26843,g17228,g20418,II26846,g17229,g20419,g20420,g20421,g20422,g20423,g20424,g20425,g20426,
    g20427,g20428,g20429,g20430,g20431,g20432,g20433,g20434,g20435,g20436,g20437,g20438,II26868,g17234,g20439,II26871,
    g17235,g20440,II26874,g17236,g20441,g20442,g20443,g20444,g20445,g20446,g20447,g20448,g20449,g20450,g20451,g20452,
    g20453,g20454,g20455,g20456,II26892,g17246,g20457,II26895,g17247,g20458,II26898,g17248,g20459,g20461,g20462,g20463,
    g20464,g20465,g20466,g20467,g20468,II26910,g17269,g20469,II26913,g17270,g20470,II26916,g17271,g20471,g20476,g20477,
    II26923,g17302,g20478,II26926,g17303,g20479,II26931,g17340,g20484,II26934,g17341,g20485,g20490,II26940,g17383,g20491,
    g20496,II26947,g17429,g20498,g20500,g20501,g20504,g20505,g20507,II26960,g20513,g20516,g20517,g20518,II26966,g20519,
    g20526,II26972,g20531,g20534,g20535,g20536,II26980,g20539,g20545,II26985,g20550,g20553,g20554,II26990,II26993,II26996,
    II26999,II27002,II27005,II27008,II27011,II27014,II27017,II27020,II27023,II27026,II27029,II27032,II27035,II27038,II27041,II27044,
    II27047,II27050,II27053,II27056,II27059,II27062,II27065,II27068,II27071,II27074,II27077,II27080,II27083,II27086,II27089,II27092,
    II27095,II27098,II27101,II27104,II27107,II27110,II27113,II27116,II27119,II27122,II27125,II27128,II27131,II27134,II27137,II27140,
    II27143,II27146,II27149,II27152,II27155,II27158,II27161,II27164,II27167,II27170,II27173,II27176,II27179,II27182,II27185,II27188,
    II27191,II27194,II27197,II27200,II27203,II27206,II27209,II27212,II27215,II27218,II27221,II27225,g20634,II27228,g20637,II27232,
    g20641,II27235,g20644,II27240,g20649,II27243,g20652,II27246,g20655,II27250,g20659,II27253,g20662,II27257,g20666,II27260,
    g20669,II27264,g20673,II27267,g20676,II27270,g20679,II27275,g20684,II27278,g20687,II27281,g20690,II27285,g20694,II27288,
    g20697,II27293,g20704,II27297,g20708,II27300,g20711,II27303,g20714,II27308,g20719,II27311,g20722,II27314,g20725,II27318,
    g20729,II27321,g20732,II27324,g20735,II27328,g20739,II27332,g20743,II27335,g20746,II27338,g20749,II27343,g20754,II27346,
    g20757,II27349,g20760,II27352,g20763,II27355,g20766,II27358,g20769,II27361,g20772,II27365,g20776,II27369,g20780,II27372,
    g20783,II27375,g20786,II27379,g20790,II27382,g20793,II27385,g20796,II27388,g20799,II27391,g20802,II27395,g20806,II27399,
    g20810,II27402,g20813,II27405,g20816,II27408,g20819,II27411,g20822,II27416,g20827,II27419,g20830,II27422,g20833,II27426,
    g20837,g20842,g20850,g20858,g20866,g20885,g19865,g20904,g19896,g20928,g19921,II27488,g20310,g20942,II27491,g20314,
    g20943,g20956,g19936,II27516,g20333,g20971,II27531,g20343,g20984,II27534,g20985,II27537,g20986,II27549,g20353,g20998,
    II27565,g21012,II27577,g20375,g21024,II27585,g20376,g21030,II27593,g21036,g21050,II27614,g21057,II27621,g20417,g21064,
    g21066,g21069,g21076,g21079,II27646,g21087,g21090,g21093,II27658,g21099,g21102,II27667,g21108,II27672,g21113,II27684,
    g21125,II27689,g21130,II27705,g21144,II27727,g21164,II27749,g19954,g21184,g21187,II27766,g19984,g21199,g21202,II27779,
    g20022,g21214,g21217,II27785,g20064,g21222,g21225,g21241,g21249,g21258,g21266,II27822,g21271,II27827,g21278,II27832,
    g21285,II27838,g21293,II27868,g19144,g21327,II27897,g19149,g21358,II27900,g21359,II27917,g19153,g21376,II27920,g19154,
    g21377,II27927,g21382,II27942,g19157,g21399,g21400,II27949,g21404,II27958,g21415,II27969,g19162,g21426,II27972,g19163,
    g21427,II27976,g21429,II27984,g21441,II27992,g21449,II28000,g19167,g21457,II28003,g21458,g21461,II28009,g20473,g21473,
    II28013,g21477,II28019,g21483,II28027,g21491,II28031,g19172,g21495,II28034,g19173,g21496,II28038,g21498,II28043,g21505,
    g21508,II28047,g20481,g21514,II28051,g21518,II28057,g21524,II28061,g19178,g21528,g21529,II28065,g21530,II28072,g21537,
    II28076,g21541,g21544,II28080,g20487,g21550,II28084,g21554,II28087,g19184,g21557,II28090,g20008,g21558,II28093,g21561,
    g21565,II28100,g21566,II28107,g21573,II28111,g21577,g21580,II28115,g20493,g21586,II28119,g21590,II28123,g21594,g21598,
    II28130,g21599,II28137,g21606,II28143,g21612,II28148,g21619,II28152,g21623,g21627,II28159,g21628,II28169,g21640,II28174,
    g21647,II28178,g21651,II28184,g19103,g21655,g21661,II28201,g21671,II28206,g21678,II28210,g20537,g21682,g21690,II28229,
    g21700,II28235,g20153,g21708,g21716,g21726,g21742,g21752,g21766,g21782,II28314,g19152,g21795,II28357,g20497,g21824,
    II28360,g21825,g21861,g21867,g21872,g21876,g21883,g21886,g21895,g21902,g21907,II28432,g21914,II28435,g21917,g21921,
    g21927,II28443,g21928,II28447,g21932,II28450,g21935,g21939,II28455,II28458,II28461,II28464,II28467,II28470,II28473,II28476,
    II28479,II28482,II28485,II28488,II28491,II28494,II28497,II28500,II28503,II28506,II28509,II28512,II28515,II28518,II28521,II28524,
    II28527,g21407,g21967,II28541,g21467,g21982,II28550,g21432,g21995,II28557,g22003,II28564,g21385,g22014,II28628,g21842,
    g22082,II28649,g21843,g22107,II28671,g21845,g22133,II28693,g21847,g22156,II28712,g21851,g22176,g22212,g22213,g22217,
    II28781,g21331,g22219,g22221,g22222,II28789,g21878,g22225,II28792,g21880,g22226,g22230,II28800,g21316,g22232,g22233,
    g22236,g22237,g22239,g22240,g22241,II28813,g21502,g22243,g22246,g22248,g22251,g22252,II28825,g21882,g22253,g22256,
    g22257,g22258,II28833,g21470,g22259,g22260,g22261,g22262,g22266,g22268,g22271,g22274,g22275,g22276,g22277,g22278,
    g22279,g22283,g22286,g22287,g22290,g22293,g22294,g22295,g22296,g22297,g22298,II28876,g21238,g22300,g22303,g22304,
    g22306,g22307,g22310,g22313,g22314,g22315,g22316,g21149,g22318,g22319,g21228,II28896,g21246,g22328,g22331,g22332,
    g22334,g22335,g22338,g22341,g21169,g22343,g22344,g21233,II28913,g21255,g22353,g22356,g22357,g22359,g22360,g22364,
    g21189,g22366,g22367,g21242,II28928,g21263,g22376,g22379,g22380,g22384,g21204,g22386,g22387,g21250,g22401,g21533,
    g22402,g21569,g22403,g21602,g22404,g21631,II28949,g21685,g22405,g22408,II28953,g21659,g22409,II28956,g21714,g22412,
    II28959,g21636,g22415,II28962,g21721,g22418,g22421,II28966,g20633,g22422,II28969,g21686,g22425,II28972,g21736,g22428,
    II28975,g21688,g22431,II28978,g21740,g22434,II28981,g21667,g22437,II28984,g21747,g22440,g22443,II28988,g20874,g22444,
    II28991,g20648,g22445,II28994,g21715,g22448,II28997,g21759,g22451,II29001,g20658,g22455,II29004,g21722,g22458,II29007,
    g21760,g22461,II29010,g21724,g22464,II29013,g21764,g22467,II29016,g21696,g22470,II29019,g21771,g22473,g22476,II29023,
    g20672,g22477,II29026,g21737,g22480,II29030,g20683,g22484,II29033,g21741,g22487,II29036,g21775,g22490,II29040,g20693,
    g22494,II29043,g21748,g22497,II29046,g21776,g22500,II29049,g21750,g22503,II29052,g21780,g22506,II29055,g21732,g22509,
    II29058,g20703,g22512,II29064,g20875,g22518,II29067,g20876,g22519,II29070,g20707,g22520,II29073,g21761,g22523,II29077,
    g20718,g22527,II29080,g21765,g22530,II29083,g21790,g22533,II29087,g20728,g22537,II29090,g21772,g22540,II29093,g21791,
    g22543,g22547,II29098,g20879,g22548,II29101,g20880,g22549,II29104,g20881,g22550,II29107,g21435,g22551,II29110,g20738,
    g22552,II29116,g20882,g22558,II29119,g20883,g22559,II29122,g20742,g22560,II29125,g21777,g22563,II29129,g20753,g22567,
    II29132,g21781,g22570,II29135,g21804,g22573,II29142,g20682,g22582,II29145,g20891,g22583,II29148,g20892,g22584,II29151,
    g20893,g22585,II29154,g20894,g22586,g22588,II29159,g20896,g22589,II29162,g20897,g22590,II29165,g20898,g22591,II29168,
    g20775,g22592,II29174,g20899,g22598,II29177,g20900,g22599,II29180,g20779,g22600,II29183,g21792,g22603,g22609,II29191,
    g20901,g22611,II29194,g20902,g22612,II29197,g20903,g22613,II29203,g20717,g22619,II29206,g20910,g22620,II29209,g20911,
    g22621,II29212,g20912,g22622,II29215,g20913,g22623,g22625,II29220,g20915,g22626,II29223,g20916,g22627,II29226,g20917,
    g22628,II29229,g20805,g22629,II29235,g20918,g22635,II29238,g20919,g22636,II29243,g20921,g22639,II29246,g20922,g22640,
    II29249,g20923,g22641,II29252,g20924,g22642,g22645,II29259,g20925,g22647,II29262,g20926,g22648,II29265,g20927,g22649,
    II29271,g20752,g22655,II29274,g20934,g22656,II29277,g20935,g22657,II29280,g20936,g22658,II29283,g20937,g22659,g22661,
    II29288,g20939,g22662,II29291,g20940,g22663,II29294,g20941,g22664,II29301,g20944,g22669,II29304,g20945,g22670,II29307,
    g20946,g22671,II29310,g20947,g22672,II29313,g20948,g22673,II29317,g20949,g22675,II29320,g20950,g22676,II29323,g20951,
    g22677,II29326,g20952,g22678,g22681,II29333,g20953,g22683,II29336,g20954,g22684,II29339,g20955,g22685,II29345,g20789,
    g22691,II29348,g20962,g22692,II29351,g20963,g22693,II29354,g20964,g22694,II29357,g20965,g22695,II29360,g21796,g22696,
    II29366,g20966,g22702,II29369,g20967,g22703,II29372,g20968,g22704,II29375,g20969,g22705,II29378,g20970,g22706,II29383,
    g20972,g22709,II29386,g20973,g22710,II29389,g20974,g22711,II29392,g20975,g22712,II29395,g20976,g22713,II29399,g20977,
    g22715,II29402,g20978,g22716,II29405,g20979,g22717,II29408,g20980,g22718,g22721,II29415,g20981,g22723,II29418,g20982,
    g22724,II29421,g20983,g22725,II29426,g20989,g22728,II29429,g20990,g22729,II29432,g20991,g22730,II29435,g20992,g22731,
    II29439,g20993,g22733,II29442,g20994,g22734,II29445,g20995,g22735,II29448,g20996,g22736,II29451,g20997,g22737,II29456,
    g20999,g22740,II29459,g21000,g22741,II29462,g21001,g22742,II29465,g21002,g22743,II29468,g21003,g22744,II29472,g21004,
    g22746,II29475,g21005,g22747,II29478,g21006,g22748,II29481,g21007,g22749,II29484,g21903,g22750,g22753,II29490,g21009,
    g22756,II29493,g21010,g22757,II29496,g21011,g22758,II29500,g21015,g22760,II29503,g21016,g22761,II29506,g21017,g22762,
    II29509,g21018,g22763,II29513,g21019,g22765,II29516,g21020,g22766,II29519,g21021,g22767,II29522,g21022,g22768,II29525,
    g21023,g22769,II29530,g21025,g22772,II29533,g21026,g22773,II29536,g21027,g22774,II29539,g21028,g22775,II29542,g21029,
    g22776,g22777,II29547,g21031,g22785,II29550,g21032,g22786,g22787,II29556,g21033,g22790,II29559,g21034,g22791,II29562,
    g21035,g22792,II29566,g21039,g22794,II29569,g21040,g22795,II29572,g21041,g22796,II29575,g21042,g22797,II29579,g21043,
    g22799,II29582,g21044,g22800,II29585,g21045,g22801,II29588,g21046,g22802,II29591,g21047,g22803,g22805,g21894,g22806,
    g21615,II29600,g21720,g22812,II29603,g21051,g22824,II29606,g21364,g22825,II29610,g21052,g22827,II29613,g21053,g22828,
    g22829,II29619,g21054,g22832,II29622,g21055,g22833,II29625,g21056,g22834,II29629,g21060,g22836,II29632,g21061,g22837,
    II29635,g21062,g22838,II29638,g21063,g22839,II29641,g20825,g22840,g22843,g21889,g22847,g21643,II29653,g21746,g22852,
    II29656,g21070,g22864,II29660,g21071,g22866,II29663,g21072,g22867,g22868,II29669,g21073,g22871,II29672,g21074,g22872,
    II29675,g21075,g22873,g22875,g21884,g22882,g21674,II29687,g21770,g22887,II29690,g21080,g22899,II29694,g21081,g22901,
    II29697,g21082,g22902,II29700,g20700,g22903,g22907,g21711,g22917,g21703,II29712,g21786,g22922,II29715,g21094,g22934,
    II29724,g22945,II29727,g20877,g22948,g22949,g21665,g22954,g21739,g22958,g21694,g22962,g21763,g22966,g21730,II29736,
    g20884,g22970,g22971,g21779,g22975,g21756,II29741,g21346,g22979,g22980,g21794,g22986,g22988,g22989,g22991,g22995,
    g22996,g22998,g23001,g23002,g23006,g23007,g23008,g23012,g23015,g23016,g23020,g23021,g23024,g23028,g23031,g23032,
    g23036,g23037,g23038,g23041,g23045,g23048,g23049,II29797,g23050,II29802,g23055,g23056,g23057,g23060,g23064,II29812,
    g23065,II29817,g23068,g23069,g23074,g23075,II29827,g23078,g23079,g23082,g23087,g23088,II29841,g23094,g23095,g23098,
    g23103,II29852,g23105,g23112,g23115,II29863,g23116,II29872,g23125,II29881,g23134,g23140,g23141,g23142,g23143,g23144,
    g23145,g23146,g23147,II29897,II29900,II29903,II29906,II29909,II29912,II29915,II29918,II29921,II29924,II29927,II29930,II29933,
    II29936,II29939,II29942,II29945,II29948,II29951,II29954,II29957,II29960,II29963,II29966,II29969,II29972,II29975,II29978,II29981,
    II29984,II29987,II29990,II29993,II29996,II29999,II30002,II30005,II30008,II30011,II30014,II30017,II30020,II30023,II30026,II30029,
    II30032,II30035,II30038,II30041,II30044,II30047,II30050,II30053,II30056,II30059,II30062,II30065,II30068,II30071,II30074,II30077,
    II30080,II30083,II30086,II30089,II30092,II30095,II30098,II30101,II30104,II30107,II30110,II30113,II30116,II30119,II30122,II30125,
    II30128,II30131,II30134,II30137,II30140,II30143,II30146,II30149,II30152,II30155,II30158,II30161,II30164,II30167,II30170,II30173,
    II30176,II30179,II30182,II30185,II30188,II30191,II30194,II30197,II30200,II30203,II30206,II30209,II30212,II30215,II30218,II30221,
    II30224,II30227,II30230,II30233,II30236,II30239,II30242,II30245,II30248,II30251,II30254,II30257,II30260,II30263,II30266,II30269,
    II30272,II30275,II30278,II30281,II30284,II30287,II30290,II30293,II30296,II30299,II30302,II30305,II30308,II30311,II30314,II30317,
    II30320,II30323,II30326,II30329,II30332,II30335,II30338,II30341,II30344,II30347,II30350,II30353,II30356,II30359,II30362,II30365,
    II30368,II30371,II30374,II30377,II30380,II30383,II30386,II30389,II30392,II30395,II30398,II30401,II30404,II30407,g23403,g23052,
    g23410,g23071,g23415,g23084,g23420,g23089,g23424,g23100,g23429,g23107,g23435,g23120,II30467,g23000,g23438,II30470,
    g23117,g23439,g23441,g23129,g23444,II30476,g22876,g23448,II30480,g23014,g23452,II30483,g23126,g23453,II30486,g23022,
    g23454,II30489,g22911,g23455,II30493,g23030,g23459,II30496,g23137,g23460,II30501,g23039,g23463,II30504,g22936,g23464,
    II30508,g23047,g23468,II30511,g21970,g23469,g23470,g22188,II30516,g23058,g23472,II30519,g22942,g23473,II30525,g23067,
    g23481,g23482,g22197,II30531,g23076,g23485,II30536,g23081,g23492,g23493,g22203,II30544,g23092,g23500,II30547,g23093,
    g23501,II30552,g23097,g23508,g23509,g22209,II30560,g23110,g23516,II30563,g23111,g23517,II30568,g23114,g23524,II30575,
    g23123,g23531,II30578,g23124,g23532,II30586,g23132,g23542,II30589,g23133,g23543,II30594,g22025,g23546,II30598,g22027,
    g23548,II30601,g22028,g23549,II30607,g22029,g23553,II30611,g22030,g23555,II30614,g22031,g23556,II30617,g22032,g23557,
    II30623,g22033,g23561,II30626,g22034,g23562,II30632,g22035,g23566,II30636,g22037,g23568,II30639,g22038,g23569,II30642,
    g22039,g23570,II30648,g22040,g23574,II30651,g22041,g23575,II30654,g22042,g23576,II30660,g22043,g23580,II30663,g22044,
    g23581,II30669,g22045,g23585,II30673,g22047,g23587,II30676,g22048,g23588,II30679,g22049,g23589,II30686,g23136,g23594,
    II30689,g22054,g23595,II30692,g22055,g23596,II30695,g22056,g23597,II30701,g22057,g23601,II30704,g22058,g23602,II30707,
    g22059,g23603,II30713,g22060,g23607,II30716,g22061,g23608,II30722,g22063,g23612,II30725,g22064,g23613,II30728,g22065,
    g23614,II30735,g22066,g23619,II30738,g22067,g23620,II30741,g22068,g23621,II30748,g21969,g23626,II30751,g22073,g23627,
    II30754,g22074,g23628,II30757,g22075,g23629,II30763,g22076,g23633,II30766,g22077,g23634,II30769,g22078,g23635,II30776,
    g22079,g23640,II30779,g22080,g23641,II30782,g22081,g23642,II30786,g22454,g23644,II30797,g22087,g23661,II30800,g22088,
    g23662,II30803,g22089,g23663,II30810,g22090,g23668,II30813,g22091,g23669,II30816,g22092,g23670,II30823,g21972,g23675,
    II30826,g22097,g23676,II30829,g22098,g23677,II30832,g22099,g23678,II30838,g22100,g23682,II30841,g22101,g23683,II30844,
    g22102,g23684,II30847,g22103,g23685,II30854,g22104,g23690,II30857,g22105,g23691,II30860,g22106,g23692,II30864,g22493,
    g23694,II30875,g22112,g23711,II30878,g22113,g23712,II30881,g22114,g23713,II30888,g22115,g23718,II30891,g22116,g23719,
    II30894,g22117,g23720,II30901,g21974,g23725,II30905,g22122,g23727,II30908,g22123,g23728,II30911,g22124,g23729,II30914,
    g22125,g23730,II30917,g23731,II30922,g22126,g23736,II30925,g22127,g23737,II30928,g22128,g23738,II30931,g22129,g23739,
    II30938,g22130,g23744,II30941,g22131,g23745,II30944,g22132,g23746,II30948,g22536,g23748,II30959,g22138,g23765,II30962,
    g22139,g23766,II30965,g22140,g23767,II30973,g22141,g23773,II30976,g22142,g23774,II30979,g22143,g23775,II30985,g22992,
    g23779,II30988,g22145,g23782,II30991,g22146,g23783,II30994,g22147,g23784,II30997,g22148,g23785,II31000,g23786,II31005,
    g22149,g23791,II31008,g22150,g23792,II31011,g22151,g23793,II31014,g22152,g23794,II31021,g22153,g23799,II31024,g22154,
    g23800,II31027,g22155,g23801,II31031,g22576,g23803,II31043,g22161,g23821,II31050,g22162,g23826,II31053,g22163,g23827,
    II31056,g22164,g23828,II31062,g23003,g23832,II31065,g22166,g23835,II31068,g22167,g23836,II31071,g22168,g23837,II31074,
    g22169,g23838,II31077,g23839,II31082,g22170,g23844,II31085,g22171,g23845,II31088,g22172,g23846,II31091,g22173,g23847,
    g23853,II31102,g22177,g23856,II31109,g22178,g23861,II31112,g22179,g23862,II31115,g22180,g23863,II31121,g23017,g23867,
    II31124,g22182,g23870,II31127,g22183,g23871,II31130,g22184,g23872,II31133,g22185,g23873,II31136,g23874,II31141,g23879,
    II31144,g22935,g23882,g23885,g22062,g23887,II31152,g22191,g23890,II31159,g22192,g23895,II31162,g22193,g23896,II31165,
    g22194,g23897,II31171,g23033,g23901,g23905,g22046,g23908,II31181,g22200,g23911,II31188,g21989,g23916,g23918,g22036,
    II31195,g22578,g23923,g23940,II31205,g22002,g23943,II31213,g22615,g23955,II31226,g22651,g23984,II31232,g22026,g24000,
    II31235,g22218,g24001,II31244,g22687,g24014,II31250,g22953,g24030,II31253,g22231,g24033,II31257,g22234,g24035,g24047,
    g23023,II31266,g22242,g24051,II31270,g22247,g24053,II31274,g22249,g24055,g24060,g23040,II31282,g22263,g24064,II31286,
    g22267,g24066,II31290,g22269,g24068,g24073,g23059,II31298,g22280,g24077,II31302,g22284,g24079,g24084,g23077,II31310,
    g22299,g24088,g24094,g22339,g24095,g22362,g24096,g24097,g22382,g24098,g24099,g24101,g24102,g24103,g22397,g24104,
    g24105,g24106,g24107,g24108,g24110,g24111,g24112,g24113,g24114,g24115,g22381,g24121,g24122,g24123,g24124,g24125,
    g24127,g24128,g24129,g24130,g24131,g24132,g24133,g24134,g22396,g24140,g24141,g24142,g24143,g24144,g24146,g24147,
    g24148,g24149,g24150,g24151,g24152,g24153,g22399,g24159,g24160,g24161,g24162,g24163,g24164,g24165,g24166,g24167,
    g24168,g22400,g24175,g24176,g24177,g24180,II31387,g22811,g24183,g24210,g24220,II31417,g24233,II31426,g24240,II31436,
    g24248,g24251,II31445,g24255,II31451,II31454,II31457,II31460,II31463,II31466,II31469,II31472,II31475,II31478,II31481,II31484,
    II31487,II31490,II31493,II31496,II31499,II31502,II31505,II31508,II31511,II31514,II31517,II31520,II31523,II31526,II31529,II31532,
    II31535,II31538,II31541,II31544,II31547,II31550,II31553,II31556,II31559,II31562,II31565,II31568,II31571,II31574,II31577,II31580,
    II31583,II31586,II31589,II31592,II31595,II31598,II31601,II31604,II31607,II31610,II31613,II31616,II31619,II31622,II31625,II31628,
    II31631,II31634,II31637,II31640,II31643,II31646,II31649,II31652,II31655,II31658,II31661,II31664,II31667,II31670,II31673,II31676,
    II31679,II31682,II31685,II31688,II31691,II31694,II31697,II31700,II31703,II31706,II31709,II31712,II31715,II31718,II31721,II31724,
    II31727,II31730,II31733,II31736,II31739,II31742,II31745,II31748,II31751,II31754,II31757,II31760,II31763,II31766,II31769,II31772,
    II31775,II31778,II31781,II31784,II31787,II31790,II31793,II31796,II31799,II31802,II31805,II31808,II31811,II31814,II31817,II31820,
    II31823,II31826,II31829,II31832,II31835,II31838,II31841,II31844,II31847,II31850,II31853,II31856,II31859,II31862,II31865,II31868,
    II31871,II31874,II31877,II31880,II31883,II31886,II31889,II31892,II31895,II31898,II31901,II31904,II31907,II31910,II31913,II31916,
    II31919,II31922,II31925,II31928,II31931,II31934,II31937,II31940,II31943,II31946,II31949,g24482,II32042,g23399,g24518,II32057,
    g23406,g24531,II32067,g24174,g24539,II32074,g23413,g24544,II32081,g24178,g24549,II32085,g24179,g24551,II32092,g23418,
    g24556,II32098,g24181,g24560,II32102,g24182,g24562,II32109,g24206,g24567,II32112,g24207,g24568,II32116,g24208,g24570,
    II32120,g24209,g24572,II32126,g24212,g24576,II32129,g24213,g24577,II32133,g24214,g24579,II32137,g24215,g24581,II32140,
    g24216,g24582,II32143,g24218,g24583,II32146,g24219,g24584,II32150,g24222,g24586,II32153,g24223,g24587,II32156,g24225,
    g24588,II32159,g24226,g24589,II32164,g24228,g24592,II32167,g24230,g24593,II32170,g24231,g24594,II32175,g24235,g24597,
    II32178,g24237,g24598,II32181,g24238,g24599,II32184,g23497,g24600,II32189,g24243,g24605,II32193,g23513,g24607,II32198,
    g24250,g24612,II32203,g23528,g24619,II32210,g23539,g24630,g24648,g24668,g24687,g24704,II32248,g23919,II32251,g24735,
    II32281,g23950,g24763,II32320,g23979,g24784,II32365,g24009,g24805,g24815,II32388,g23385,g24816,II32419,g24043,g24827,
    g24834,II32439,g23392,g24835,g24850,II32487,g23400,g24851,II32506,g23324,g24856,g24864,II32535,g23407,g24865,II32556,
    g23329,g24872,II32583,g23330,g24879,II32604,g23339,g24886,g24893,g23486,II32642,g23348,g24903,g24912,g23495,g24916,
    g23502,g24929,g23511,g24933,g23518,g24939,g23660,g24941,g23526,g24945,g23533,II32704,g23357,g24949,g24950,g23710,
    g24952,g23537,II32716,g23358,g24956,II32719,g23359,g24957,g24958,g23478,g24962,g23764,g24969,g23489,g24973,g23819,
    g24982,g23505,g24993,g23521,g25087,g25094,g25095,II32829,g24059,g25103,g25104,g25105,II32835,g24072,g25109,g25110,
    g25111,g25115,g25116,II32844,g25118,II32847,g24083,g25119,g25120,II32851,g25121,II32854,g24092,g25122,II32857,g25123,
    II32860,g25124,g25126,II32868,II32871,II32874,II32877,II32880,II32883,II32886,II32889,II32892,II32895,II32898,II32901,II32904,
    II32907,II32910,II32913,II32916,II32919,II32922,II32925,II32928,II32931,II32934,II32937,II32940,II32943,II32946,II32949,II32952,
    II32955,II32958,II32961,II32964,II32967,II32970,II32973,II32976,II32979,II32982,II32985,II32988,II32991,II32994,II32997,II33000,
    II33003,II33006,II33009,II33013,g25179,II33016,g25180,g25274,g25283,g25291,II33128,g24975,g25296,g25301,g25305,g24880,
    II33136,g24986,g25306,g25313,g24868,g25314,g24897,II33145,g24997,g25315,g25319,g24857,g25322,g24883,g25323,g24920,
    II33154,g25005,g25324,II33157,g25027,g25327,g25329,g24844,g25330,g24873,g25332,g24900,g25333,g24937,g25335,g24832,
    II33168,g25042,g25336,g25338,g24860,g25339,g24887,g25341,g24923,g25347,g24817,g25349,g24848,II33182,g25056,g25350,
    g25352,g24875,g25353,g24904,II33188,g24814,g25354,g25355,g24797,g25361,g24837,g25363,g24862,II33198,g25067,g25364,
    g25366,g24889,g25367,g24676,g25368,g24778,II33205,g24833,g25369,g25370,g24820,g25376,g24852,g25378,g24877,g25379,
    g25383,g24766,g25384,g24695,g25385,g24801,II33219,g24849,g25386,g25387,g24839,g25393,g24866,g25394,g24753,g25395,
    g25399,g24787,g25400,g24712,g25401,g24823,II33232,g24863,g25402,g25403,g24854,g25404,g24771,g25405,g25409,g24808,
    g25410,g24723,g25411,g24842,g25412,g24791,g25413,g25417,g24830,g25419,g24812,II33246,g24890,II33249,g25421,g25422,
    g25430,g24616,g25431,II33257,g24909,II33260,g25436,g25437,g24627,g25438,II33265,g24925,II33268,g25443,g25444,g24641,
    g25445,g25449,g24660,II33278,g25088,g25454,II33282,g25096,g25458,II33286,g24426,g25462,II33289,g25106,g25463,II33293,
    g25008,g25467,II33297,g24430,g25471,II33300,g25112,g25472,II33304,g25004,g25476,II33307,g25011,g25479,II33312,g25014,
    g25484,II33316,g24434,g25488,II33321,g24442,g25493,II33324,g25009,g25496,II33327,g25017,g25499,II33330,g25019,g25502,
    II33335,g25010,g25507,II33338,g25021,g25510,II33343,g25024,g25515,II33347,g24438,g25519,II33352,g24443,g25524,II33355,
    g25012,g25527,II33358,g25028,g25530,II33361,g25013,g25533,II33364,g25029,g25536,II33368,g24444,g25540,II33371,g25015,
    g25543,II33374,g25031,g25546,II33377,g25033,g25549,II33382,g25016,g25554,II33385,g25035,g25557,II33390,g25038,g25562,
    II33396,g24447,g25573,II33399,g25018,g25576,II33402,g24448,g25579,II33405,g25020,g25582,II33408,g25040,g25585,II33411,
    g24491,g25588,II33415,g24449,g25590,II33418,g25022,g25593,II33421,g25043,g25596,II33424,g25023,g25599,II33427,g25044,
    g25602,II33431,g24450,g25606,II33434,g25025,g25609,II33437,g25046,g25612,II33440,g25048,g25615,II33445,g25026,g25620,
    II33448,g25050,g25623,g25630,g24478,II33457,g24451,g25634,II33460,g24452,g25637,II33463,g25030,g25640,II33466,g25053,
    g25643,II33469,g24498,g25646,II33472,g24499,g25647,II33476,g24453,g25652,II33479,g25032,g25655,II33482,g24454,g25658,
    II33485,g25034,g25661,II33488,g25054,g25664,II33491,g24501,g25667,II33495,g24455,g25669,II33498,g25036,g25672,II33501,
    g25057,g25675,II33504,g25037,g25678,II33507,g25058,g25681,II33511,g24456,g25685,II33514,g25039,g25688,II33517,g25060,
    g25691,II33520,g25062,g25694,g25698,II33526,g24457,g25700,II33529,g25041,g25703,II33532,g24507,g25706,II33535,g24508,
    g25707,II33539,g24458,g25711,II33542,g24459,g25714,II33545,g25045,g25717,II33548,g25064,g25720,II33551,g24510,g25723,
    II33554,g24511,g25724,II33558,g24460,g25729,II33561,g25047,g25732,II33564,g24461,g25735,II33567,g25049,g25738,II33570,
    g25065,g25741,II33573,g24513,g25744,II33577,g24462,g25746,II33580,g25051,g25749,II33583,g25068,g25752,II33586,g25052,
    g25755,II33589,g25069,g25758,II33593,g24445,g25762,II33596,g24446,g25763,II33600,g24463,g25767,II33603,g24519,g25770,
    g25771,II33608,g24464,g25773,II33611,g25055,g25776,II33614,g24521,g25779,II33617,g24522,g25780,II33621,g24465,g25784,
    II33624,g24466,g25787,II33627,g25059,g25790,II33630,g25071,g25793,II33633,g24524,g25796,II33636,g24525,g25797,II33640,
    g24467,g25802,II33643,g25061,g25805,II33646,g24468,g25808,II33649,g25063,g25811,II33652,g25072,g25814,II33655,g24527,
    g25817,II33659,g24469,g25821,II33662,g24532,g25824,g25825,II33667,g24470,g25827,II33670,g25066,g25830,II33673,g24534,
    g25833,II33676,g24535,g25834,II33680,g24471,g25838,II33683,g24472,g25841,II33686,g25070,g25844,II33689,g25074,g25847,
    II33692,g24537,g25850,II33695,g24538,g25851,II33700,g24474,g25856,II33703,g24545,g25859,g25860,II33708,g24475,g25862,
    II33711,g25073,g25865,II33714,g24547,g25868,II33717,g24548,g25869,II33723,g24477,g25877,II33726,g24557,g25880,II33732,
    g24473,g25886,II33737,g24476,g25891,g25895,g25899,g24928,g25903,g25907,g24940,g25911,g25915,g24951,g25919,g25923,
    g24963,g25937,g25939,g25942,g25945,g25952,II33790,g25976,II33798,g25982,II33801,II33804,II33807,II33810,II33813,II33816,
    II33819,II33822,II33825,II33828,II33831,II33834,II33837,II33840,II33843,II33846,II33849,II33852,II33855,II33858,II33861,II33864,
    II33867,II33870,II33873,II33876,II33879,II33882,II33885,II33888,II33891,II33894,II33897,II33900,II33903,II33906,II33909,II33912,
    II33915,II33918,II33954,g25343,g26056,II33961,g25357,g26063,II33968,g25372,g26070,II33974,g25389,g26076,II33984,g25932,
    g26086,II33990,g25870,g26092,II33995,g25935,g26102,II33999,g25490,II34002,g26105,II34009,g25882,g26114,II34012,g25938,
    g26118,II34017,g25887,g26121,II34020,g25940,g26125,II34026,g25892,g26131,II34029,g25520,II34032,g26136,II34041,g25566,
    II34044,g26150,II34051,g25204,g26159,II34056,g25206,g26164,II34059,g25207,g26165,II34063,g25209,g26167,II34068,g25211,
    g26172,II34071,g25212,g26173,II34074,g25213,g26174,II34077,g25954,g26175,II34080,g25539,g26178,II34083,g25214,g26181,
    II34086,g25215,g26182,II34091,g25217,g26187,g26189,II34096,g25218,g26190,II34099,g25219,g26191,II34102,g25220,g26192,
    II34105,g25221,g26193,II34108,g25222,g26194,II34111,g25223,g26195,II34114,g25958,g26196,II34118,g25605,g26202,II34121,
    g25224,g26205,II34124,g25225,g26206,II34128,g25227,g26208,g26209,II34132,g25228,g26210,II34135,g25229,g26211,II34140,
    g25230,g26214,II34143,g25231,g26215,II34146,g25232,g26216,II34150,g25233,g26220,II34153,g25234,g26221,II34156,g25235,
    g26222,II34159,g25964,g26223,II34162,g25684,g26226,II34165,g25236,g26229,II34168,g25237,g26230,II34172,g25239,g26232,
    g26237,II34180,g25240,g26238,II34183,g25241,g26239,II34189,g25242,g26245,II34192,g25243,g26246,II34195,g25244,g26247,
    II34198,g25245,g26248,II34201,g25246,g26249,II34204,g25247,g26250,II34207,g25969,g26251,II34210,g25761,g26254,II34220,
    g25248,g26264,g26275,II34230,g25249,g26276,II34233,g25250,g26277,II34238,g25251,g26280,II34241,g25252,g26281,II34244,
    g25253,g26282,II34254,g25185,g26294,II34266,g25255,g26308,g26313,II34274,g25256,g26314,II34277,g25257,g26315,II34296,
    g25189,g26341,II34306,g25259,g26349,II34313,g25265,g26354,II34316,g25191,g26355,II34321,g25928,g26358,II34327,g25260,
    g26364,II34343,g25194,g26385,II34353,g25927,g26393,II34358,g25262,g26398,II34363,g25930,g26401,II34369,g25263,g26407,
    II34385,g25197,g26428,II34388,g25200,g26429,II34392,g25266,g26433,II34395,g25929,g26434,II34400,g25267,g26439,II34405,
    g25933,g26442,II34411,g25268,g26448,II34421,g25203,g26461,II34425,g25270,g26465,II34428,g25931,g26466,II34433,g25271,
    g26471,II34438,g25936,g26474,II34444,g25272,g26480,g26481,g25764,II34449,g25205,g26485,II34453,g25279,g26489,II34456,
    g25934,g26490,II34461,g25280,g26495,II34464,g25199,g26496,g26497,g25818,II34469,g25210,g26501,II34473,g25288,g26505,
    II34476,g25201,g26506,II34479,g25202,g26507,g26508,g25312,g26512,g25853,g26516,g25320,g26520,g25874,g26521,g25331,
    g26525,g25340,g26533,g26538,g26539,g26540,g26542,g26543,g26544,g26546,II34505,g25450,g26548,g26549,g26550,g26551,
    g26552,g26554,g26555,g26556,g26558,g26561,g26562,g26563,g26564,g26565,g26566,g26567,g26568,g26570,g26571,g26572,
    g26574,II34535,g25451,g26576,g26577,g26578,g26579,g26580,g26581,g26582,g26584,g26585,g26586,g26587,g26588,g26589,
    g26590,g26591,g26593,g26594,g26595,g26597,g26598,g26599,g26600,g26601,g26602,g26603,g26604,g26605,g26606,g26608,
    g26609,g26610,g26611,g26612,g26613,g26614,g26615,g26617,II34579,g25452,g26618,g26619,g26620,g26621,g26622,g26623,
    g26624,g26625,g26626,g26627,g26628,g26629,g26631,g26632,g26633,g26634,g26635,g26636,g26637,g26638,g26639,g26640,
    g26641,g26642,g26643,g26644,g26645,g26646,g26647,g26648,g26649,g26650,g26651,g26652,g26653,g26654,g26656,g26657,
    g26658,g26662,II34641,II34644,II34647,II34650,II34653,II34656,II34659,II34662,II34665,II34668,II34671,II34674,II34677,II34680,
    II34683,II34686,II34689,II34692,II34695,II34698,II34701,II34704,II34707,II34710,II34713,II34716,II34719,II34722,II34725,II34728,
    II34731,II34734,II34737,II34740,II34743,II34746,II34749,II34752,II34755,II34758,II34761,II34764,II34767,II34770,II34773,II34776,
    II34779,II34782,II34785,II34788,II34791,II34794,II34797,II34800,II34803,II34806,II34809,II34812,II34815,II34818,II34821,II34824,
    II34827,II34830,II34833,II34836,II34839,II34842,II34845,II34848,II34851,II34854,II34857,II34860,II34863,II34866,II34872,g26217,
    g26757,II34879,g26240,g26762,II34901,g26295,g26782,II34909,g26265,g26788,II34916,g26793,II34921,g26796,II34946,g26534,
    g26819,II34957,g26541,g26828,II34961,g26545,g26830,II34964,g26547,g26831,II34967,g26553,g26832,II34971,g26557,g26834,
    II34974,g26168,g26835,II34977,g26559,g26836,II34980,g26458,g26837,II34983,g26569,g26840,II34986,g26160,g26841,II34990,
    g26573,g26843,II34993,g26575,g26844,II34997,g26482,g26846,II35000,g26336,g26849,II35003,g26592,g26850,II35007,g26596,
    g26852,II35011,g26304,g26854,II35014,g26498,g26855,II35017,g26616,g26858,II35028,g26513,g26861,II35031,g26529,g26864,
    II35049,g26530,g26868,II35053,g26655,g26872,II35064,g26531,g26875,II35067,g26659,g26876,II35072,g26661,g26881,II35076,
    g26532,g26883,II35079,g26664,g26884,II35083,g26665,g26886,II35087,g26667,g26890,II35092,g26669,g26895,II35095,g26670,
    g26896,II35099,g26672,g26900,II35106,g26675,g26909,II35109,g26676,g26910,II35116,g26025,g26921,g26922,g26283,g26935,
    g26327,g26944,g26374,g26950,g26417,II35136,g26660,g26953,g26954,II35141,g26666,g26956,g26957,II35146,g26671,g26959,
    g26960,II35153,g26677,g26964,II35172,g26272,g26983,g26987,g27010,g27036,g27064,II35254,g26048,g27075,II35283,g26031,
    g27102,II35297,g26199,g27114,II35301,g26037,g27116,II35313,g27126,II35319,g26183,g27132,g27133,g27134,g27135,g27136,
    g27137,g27138,g27139,g27140,g27141,g27142,g27143,II35334,g26106,g27145,g27146,g27148,II35341,g26120,g27150,g27151,
    g27153,II35347,g27154,g27155,II35351,g27156,II35355,g26130,g27158,g27159,II35360,g27161,g27162,II35364,g27163,g27164,
    II35369,g26144,g27166,g27167,II35373,g27168,II35376,g27171,g27172,g27173,II35383,g27176,g27177,II35389,g27180,II35394,
    g27183,II35399,g27186,II35404,II35407,II35410,II35413,II35416,II35419,II35422,II35425,II35428,II35431,II35434,II35437,II35440,
    II35443,II35446,II35449,II35452,II35455,II35458,II35461,II35464,II35467,II35470,II35473,II35476,II35479,II35482,II35485,II35488,
    II35491,II35494,II35497,II35500,II35503,II35506,II35509,II35512,II35515,II35518,II35521,II35524,II35527,II35530,II35533,II35536,
    II35539,II35542,II35545,II35548,II35551,II35554,g27349,II35667,g27120,g27353,II35673,g27123,g27357,II35678,g27129,g27360,
    II35681,g26869,g27361,II35686,g27131,g27366,II35689,g26878,g27367,II35695,g26887,g27373,II35698,g26897,g27376,II35708,
    g26974,II35711,g27381,g27383,g27384,II35723,g27385,g27386,II35727,g26902,g27387,II35731,g26892,g27391,II35737,g26915,
    g27397,II35741,g27118,g27401,II35744,g26906,g27404,II35750,g26928,g27410,II35756,g27117,g27416,II35759,g27121,g27419,
    II35762,g26918,g27422,II35768,g26941,g27428,II35772,g26772,g27432,II35777,g27119,g27437,II35780,g27124,g27440,II35783,
    g26931,g27443,g27449,II35791,g26779,g27451,II35796,g27122,g27456,II35799,g27130,g27459,II35803,g26803,g27463,g27465,
    II35809,g26785,g27467,II35814,g27125,g27472,II35817,g27475,II35821,g26804,g27479,II35824,g26805,g27480,II35829,g26806,
    g27483,g27484,II35834,g26792,g27486,II35837,g26911,g27489,II35841,g26807,g27493,II35844,g26808,g27494,II35849,g26776,
    g27497,II35852,g27498,II35856,g26809,g27502,II35859,g26810,g27503,II35863,g26811,g27505,g27506,II35868,g26812,g27508,
    II35872,g26925,g27510,II35876,g26813,g27514,II35879,g26814,g27515,II35883,g26781,g27517,II35886,g27518,II35890,g26815,
    g27522,II35893,g26816,g27523,II35897,g26817,g27525,II35900,g26786,g27526,II35915,g26818,g27533,II35919,g26938,g27535,
    II35923,g26820,g27539,II35926,g26821,g27540,II35930,g26789,g27542,II35933,g27543,II35937,g26822,g27547,II35940,g26823,
    g27548,II35953,g26824,g27553,II35957,g26947,g27555,II35961,g26825,g27559,II35964,g26826,g27560,II35968,g26795,g27562,
    II35983,g26827,g27569,II36008,g26798,g27586,g27589,g27590,g27144,g27595,g27149,g27599,g27147,g27604,g27157,g27608,
    g27152,g27613,g27165,g27617,g27160,g27622,g27174,II36032,g27113,g27632,II36042,g27662,II36046,g27667,II36052,g27674,
    II36060,II36063,II36066,II36069,II36072,II36075,II36078,II36081,II36084,II36087,II36090,II36093,II36096,II36099,II36102,II36105,
    II36108,II36111,II36114,II36117,II36120,II36123,II36126,II36129,II36132,II36135,II36138,II36141,II36144,II36147,II36150,II36153,
    II36156,II36159,II36162,g27748,II36213,g27571,g27776,II36217,g27580,g27780,II36221,g27784,II36224,g27785,II36227,g27594,
    g27786,II36230,g27583,g27787,II36234,g27791,II36237,g27792,II36240,g27603,g27793,II36243,g27587,g27794,II36246,g27797,
    II36250,g27612,g27799,II36253,g27800,II36264,g27621,g27805,II36267,g27395,g27806,II36280,g27390,g27817,II36283,g27408,
    g27820,II36296,g27626,g27831,II36307,g27400,g27839,II36311,g27426,g27843,II36321,g27627,g27847,II36327,g27413,g27858,
    II36330,g27447,g27861,II36337,g27628,g27872,II36341,g27431,g27879,II36347,g27630,g27889,II36354,g27903,II36358,g27672,
    g27905,II36362,g27907,II36367,g27678,g27910,II36371,g27912,II36379,g27682,g27918,II36382,g27563,g27919,II36390,g27243,
    g27927,II36393,g27572,g27928,II36397,g27574,g27932,II36404,g27450,g27939,II36407,g27581,g27942,II36411,g27582,g27946,
    II36417,g27462,g27952,II36420,g27253,g27955,II36423,g27466,g27956,II36426,g27584,g27959,II36432,g27585,g27965,g27969,
    II36438,g27255,g27971,II36441,g27256,g27972,II36444,g27482,g27973,II36447,g27257,g27976,II36450,g27485,g27977,II36454,
    g27588,g27981,II36459,g27258,g27986,II36462,g27259,g27987,II36465,g27260,g27988,II36468,g27261,g27989,g27990,II36473,
    g27262,g27992,II36476,g27263,g27993,II36479,g27504,g27994,II36483,g27264,g27998,II36486,g27507,g27999,II36490,g27265,
    g28003,II36493,g27266,g28004,II36496,g27267,g28005,II36499,g27268,g28006,II36502,g27269,g28007,II36507,g27270,g28010,
    II36510,g27271,g28011,II36513,g27272,g28012,II36516,g27273,g28013,g28014,II36521,g27274,g28016,II36524,g27275,g28017,
    II36527,g27524,g28018,II36530,g27276,g28021,II36533,g27277,g28022,II36536,g27278,g28023,II36539,g27279,g28024,II36542,
    g27280,g28025,II36545,g27281,g28026,II36551,g27282,g28030,II36554,g27283,g28031,II36557,g27284,g28032,II36560,g27285,
    g28033,II36563,g27286,g28034,II36568,g27287,g28037,II36571,g27288,g28038,II36574,g27289,g28039,II36577,g27290,g28040,
    g28041,II36582,g27291,g28043,II36585,g27292,g28044,II36588,g27293,g28045,II36598,g27294,g28047,II36601,g27295,g28048,
    II36604,g27296,g28049,II36609,g27297,g28052,II36612,g27298,g28053,II36615,g27299,g28054,II36618,g27300,g28055,II36621,
    g27301,g28056,II36627,g27302,g28060,II36630,g27303,g28061,II36633,g27304,g28062,II36636,g27305,g28063,II36639,g27306,
    g28064,II36644,g27307,g28067,II36647,g27308,g28068,II36650,g27309,g28069,II36653,g27310,g28070,II36656,g27311,g28071,
    II36659,g27312,g28072,II36663,g27313,g28074,II36673,g27314,g28076,II36676,g27315,g28077,II36679,g27316,g28078,II36684,
    g27317,g28081,II36687,g27318,g28082,II36690,g27319,g28083,II36693,g27320,g28084,II36696,g27321,g28085,II36702,g27322,
    g28089,II36705,g27323,g28090,II36708,g27324,g28091,II36711,g27325,g28092,II36714,g27326,g28093,II36718,g27327,g28095,
    II36721,g27328,g28096,II36724,g27329,g28097,II36728,g27330,g28099,II36738,g27331,g28101,II36741,g27332,g28102,II36744,
    g27333,g28103,II36749,g27334,g28106,II36752,g27335,g28107,II36755,g27336,g28108,II36758,g27337,g28109,II36761,g27338,
    g28110,II36766,g27339,g28113,II36769,g27340,g28114,II36772,g27341,g28115,II36776,g27342,g28117,II36786,g27343,g28119,
    II36789,g27344,g28120,II36792,g27345,g28121,II36797,g27346,g28124,II36800,g27347,g28125,II36803,g27348,g28126,g28128,
    g27528,II36808,g27354,g28132,g28133,g27550,g28137,g27566,g28141,g27576,g28149,g28150,g28151,g28152,g28153,g28154,
    g28155,g28156,g28158,g28159,g28160,g28161,g28162,g28163,g28164,g28165,g28166,g28167,g28168,g28169,g28170,g28172,
    g28173,g28174,g28175,g28177,g28178,II36848,g28179,g28186,g28187,g28190,II36860,g28194,II36864,g28200,II36867,II36870,
    II36873,II36876,II36879,II36882,II36885,II36888,II36891,II36894,II36897,II36900,II36903,II36906,II36909,II36912,II36915,II36918,
    II36921,II36924,II36927,II36930,II36933,II36936,II36939,II36942,II36945,II36948,II36951,II36954,II36957,II36960,II36963,II36966,
    II36969,II36972,II36975,II36978,II36981,II36984,II36987,II36990,II36993,II36996,II36999,II37002,II37005,II37008,II37011,II37014,
    II37017,II37020,II37023,II37026,II37029,II37032,II37035,II37038,II37041,II37044,II37047,II37050,II37053,II37056,II37059,II37062,
    II37065,II37068,II37071,II37074,II37077,II37080,II37083,II37086,II37089,II37092,II37095,II37098,II37101,II37104,II37107,II37110,
    II37113,II37116,II37119,II37122,II37125,II37128,II37131,II37134,II37137,II37140,II37143,II37146,II37149,II37152,II37155,II37158,
    II37161,II37164,II37167,II37170,II37173,II37176,II37179,II37182,II37185,II37188,II37191,II37194,II37197,II37200,II37203,II37228,
    g28341,II37232,g28343,II37238,g28347,II37252,g28359,II37260,g28365,II37266,g28369,II37269,g28145,g28370,II37273,g28372,
    II37277,g28146,g28374,II37280,g28375,II37284,g28147,g28377,II37291,g28148,g28382,II37319,g28390,II37330,g28393,II37334,
    g28395,g28419,II37379,g28199,g28432,II37386,g28437,II37394,g27718,g28443,II37400,g28447,II37410,g27722,g28455,II37415,
    g28458,II37426,g27724,g28467,g28483,g28491,g28496,II37459,g27759,g28498,g28500,II37467,g27760,g28524,II37471,g27761,
    g28526,II37474,g27762,g28527,II37481,g27763,g28552,II37484,g27764,g28553,g28554,II37488,g27765,g28555,II37494,g27766,
    g28579,II37497,g27767,g28580,g28581,g28582,II37502,g27768,g28583,II37508,g27769,g28607,g28608,g28609,g28610,II37514,
    g27771,g28611,g28612,g28046,g28616,g28617,g28618,g28619,g28075,g28623,g28624,g28625,g28100,g28629,g28630,g28118,
    g28638,g28639,g28640,g28641,g28642,g28643,g28644,g28645,g28646,g28647,g28648,g28649,g28650,g28651,g28652,g28653,
    g28655,II37566,II37569,II37572,II37575,II37578,II37581,II37584,II37587,II37590,II37593,II37596,II37599,II37602,II37605,II37608,
    II37611,II37614,II37617,II37620,II37623,II37626,II37629,II37632,II37635,II37638,II37641,II37644,II37647,II37650,II37653,II37656,
    II37659,II37662,II37665,g28720,g28495,g28721,g28490,g28723,g28528,g28725,g28499,g28727,g28489,g28730,g28470,g28734,
    g28525,g28740,g28488,II37702,g28512,g28741,II37712,g28751,II37716,g28540,g28755,II37725,g28764,II37729,g28567,g28768,
    II37736,g28775,II37740,g28595,g28779,II37746,g28785,II37752,g28791,II37757,g28796,II37760,g28799,II37765,g28804,II37768,
    g28807,II37771,g28810,II37775,g28814,II37778,g28817,II37781,g28820,II37784,g28823,II37787,g28826,II37790,g28829,II37793,
    g28832,II37796,g28634,g28833,II37800,g28635,g28835,II37804,g28636,g28837,II37808,g28637,g28839,g28855,g28409,g28859,
    g28413,g28863,g28417,g28867,g28418,II37842,g28501,g28871,II37846,g28877,II37851,g28668,g28882,II37854,g28529,g28883,
    II37858,g28889,II37863,g28894,II37868,g28321,g28899,II37871,g28556,g28900,II37875,g28906,II37880,g28911,II37885,g28916,
    II37891,g28325,g28924,II37894,g28584,g28925,II37897,g28928,II37901,g28932,II37906,g28937,II37912,g28945,II37917,g28328,
    g28950,II37920,g28951,II37924,g28955,II37928,g28959,II37934,g28967,II37939,g28972,II37942,g28975,II37946,g28979,II37950,
    g28983,II37956,g28993,II37961,g28998,II37965,g29002,II37968,g29005,II37973,g29010,II37978,g29019,II37982,g29023,II37986,
    g29027,II37991,g29032,II37994,g29035,II37999,g29042,II38003,g29046,II38007,g29050,II38011,g29054,II38014,g29057,II38018,
    g28342,g29061,II38024,g29065,II38028,g29069,II38032,g28344,g29073,II38035,g28345,g29074,II38038,g28346,g29075,II38042,
    g29077,II38046,g28348,g29081,II38049,g28349,g29082,II38053,g28350,g29084,II38056,g28351,g29085,II38059,g28352,g29086,
    II38064,g28353,g29089,II38068,g28354,g29091,II38071,g28355,g29092,II38074,g28356,g29093,II38077,g28357,g29094,II38080,
    g28358,g29095,II38085,g28360,g29098,II38088,g28361,g29099,II38091,g28362,g29100,II38094,g28363,g29101,II38097,g28364,
    g29102,II38101,g28366,g29104,II38104,g28367,g29105,II38107,g28368,g29106,II38111,g28371,g29108,II38119,g28420,g29117,
    II38122,g28421,g29118,II38125,g28425,g29119,II38128,g29120,II38136,II38139,II38142,II38145,II38148,II38151,II38154,II38157,
    II38160,II38163,II38166,II38169,II38172,II38175,II38178,II38181,II38184,II38187,II38190,II38193,II38196,II38199,II38202,II38205,
    II38208,II38211,II38214,II38217,II38220,II38223,II38226,II38229,II38232,II38235,II38238,II38241,II38245,g28920,g29168,II38250,
    g28941,g29171,II38258,g28963,g29177,II38272,g29013,g29189,II38275,g28987,g29190,II38278,g29191,g29192,g28954,II38282,
    g29193,II38321,g29113,g29230,II38330,g29237,II38339,g29244,II38342,g28886,g29245,II38345,g29109,g29246,II38348,g28874,
    g29247,II38352,g29110,g29249,II38355,g29039,g29250,II38360,g29111,g29253,II38363,g29016,g29254,II38369,g29112,g29258,
    g29266,II38386,g29267,g29268,g29269,II38391,g29270,g29271,g29272,II38396,g29273,g29274,g29275,II38401,g29276,g29277,
    II38405,g29278,II38408,g29279,g29280,II38412,g29281,g29282,g29283,g29285,g29286,g29287,II38421,g29288,g29290,g29291,
    g29292,II38428,g28732,g29293,g29295,g29296,II38434,g28735,g29297,II38437,g28736,g29298,II38440,g28738,g29299,g29301,
    II38447,g28744,g29304,II38450,g28745,g29305,II38453,g28746,g29306,II38456,g28747,g29307,II38459,g28749,g29308,II38462,
    g29309,II38466,g28754,g29311,II38471,g28758,g29314,II38474,g28759,g29315,II38477,g28760,g29316,II38480,g28761,g29317,
    II38483,g28990,g29318,II38486,g28763,g29319,II38491,g28767,g29322,II38496,g28771,g29325,II38499,g28772,g29326,II38502,
    g28773,g29327,II38505,g28774,g29328,II38510,g28778,g29331,II38515,g28782,g29334,II38518,g28783,g29335,II38524,g28788,
    g29339,II38536,g29349,II38539,g29350,g29356,g29358,II38548,g28903,g29359,g29360,g29361,g29362,g29363,g29364,g29365,
    g29366,g29367,g29368,g29369,g29370,g29371,g29372,g29373,g29374,g29375,g29376,g29377,g29378,g29379,g29380,g29381,
    g29382,g29383,g29384,g29385,g29386,g29387,g29388,g29389,g29390,g29391,g29392,g29393,g29394,g29395,g29396,g29397,
    g29398,II38591,g29400,II38594,g29401,g29402,II38599,g29404,II38602,g29405,II38606,g29407,II38609,g29408,II38613,g29410,
    II38617,g29412,II38620,II38623,II38626,II38629,II38632,II38635,II38638,II38641,II38644,II38647,II38650,II38653,II38656,II38659,
    II38662,II38665,II38668,II38671,II38674,II38677,II38680,II38683,II38686,II38689,II38692,II38695,II38698,II38701,II38704,II38707,
    II38710,II38713,II38716,II38719,II38722,II38725,II38728,II38731,II38734,II38737,II38740,II38743,II38746,II38749,II38752,II38755,
    II38758,II38761,II38764,II38767,II38770,g29491,II38801,g29495,II38804,g29353,g29496,II38807,g29497,II38817,g29354,g29499,
    II38827,g29355,g29501,II38838,g29357,g29504,II38848,g29167,g29506,II38851,g29169,g29507,II38854,g29170,g29508,II38857,
    g29172,g29509,II38860,g29173,g29510,II38863,g29178,g29511,II38866,g29179,g29512,II38869,g29181,g29513,II38872,g29182,
    g29514,II38875,g29184,g29515,II38878,g29185,g29516,II38881,g29187,g29517,II38885,g29519,II38898,g29194,g29530,II38905,
    g29197,g29535,II38909,g29198,g29537,II38916,g29201,g29542,II38920,g29204,g29544,II38924,g29205,g29546,II38931,g29209,
    g29551,II38936,g29212,g29554,II38940,g29213,g29556,II38947,g29218,g29561,II38951,g29221,g29563,II38958,g29226,g29568,
    II38975,g29348,g29583,II38999,II39002,II39005,II39008,II39011,II39014,II39017,II39020,II39023,II39026,II39029,II39032,II39035,
    II39038,II39041,II39044,II39047,II39050,II39053,II39056,II39059,II39062,II39065,II39068,II39071,II39074,II39077,II39080,II39083,
    II39086,II39089,g29658,g29574,g29659,g29571,g29660,g29578,g29661,g29576,g29662,g29570,g29664,g29552,g29666,g29577,
    g29668,g29569,g29673,II39121,g29579,g29689,II39124,g29606,g29690,II39127,g29608,g29691,II39130,g29580,g29692,II39133,
    g29609,g29693,II39136,g29611,g29694,II39139,g29612,g29695,II39142,g29581,g29696,II39145,g29613,g29697,II39148,g29616,
    g29698,II39151,g29617,g29699,II39154,g29582,g29700,II39157,g29618,g29701,II39160,g29620,g29702,II39164,g29621,g29704,
    II39168,g29623,g29708,g29716,g29498,g29724,g29500,g29726,g29503,g29739,g29505,II39234,II39237,II39240,II39243,II39246,
    II39249,II39252,II39255,II39258,II39261,II39264,II39267,II39270,II39273,II39276,II39279,g29823,g29663,g29829,g29665,g29835,
    g29667,g29840,g29669,g29844,g29670,g29848,g29761,g29849,g29671,g29853,g29672,g29857,g29676,g29861,g29677,g29865,
    g29678,g29869,g29679,g29873,g29680,g29877,g29681,g29881,g29682,g29885,g29683,g29889,g29684,g29893,g29685,g29897,
    g29686,g29901,g29687,g29905,g29688,II39398,g29932,II39401,g29933,II39404,g29934,II39407,g29935,II39411,g29937,II39414,
    g29938,II39418,g29940,II39423,g29943,II39454,II39457,II39460,II39463,II39466,II39469,II39472,II39475,g30036,g29912,g30040,
    g29914,g30044,g29916,g30048,g29920,II39550,g30052,II39573,g29936,g30076,II39577,g29939,g30078,II39585,g29941,g30084,
    II39622,II39625,II39628,II39631,II39635,g30055,g30124,II39638,g30056,g30125,II39641,g30057,g30126,II39647,g30058,g30130,
    g30134,g30010,g30139,g30011,g30143,g30012,g30147,g30013,g30151,g30014,g30155,g30015,g30159,g30016,g30163,g30017,
    g30167,g30018,g30171,g30019,g30175,g30020,g30179,g30021,g30183,g30022,g30187,g30023,g30191,g30024,g30195,g30025,
    g30199,g30026,g30203,g30027,g30207,g30028,g30211,g30029,II39674,g30072,g30215,g30229,g30030,g30233,g30031,g30237,
    g30032,g30241,g30033,II39761,g30306,II39764,g30060,g30307,II39767,g30061,g30308,II39770,g30063,g30309,II39773,g30064,
    g30310,II39776,g30066,g30311,II39779,g30053,g30312,II39782,g30054,g30313,II39785,II39788,II39791,II39794,II39797,II39800,
    II39803,II39806,II39809,II39812,II39815,II39818,II39821,g30267,g30326,II39825,g30268,g30328,II39828,g30269,g30329,II39832,
    g30270,g30331,II39835,g30271,g30332,II39840,g30272,g30335,II39843,g30273,g30336,II39848,g30274,g30339,II39853,g30275,
    g30342,II39856,g30276,g30343,II39859,g30277,g30344,II39863,g30278,g30346,II39866,g30279,g30347,II39870,g30280,g30349,
    II39873,g30281,g30350,II39878,g30282,g30353,II39881,g30283,g30354,II39886,g30284,g30357,II39889,g30285,g30358,II39892,
    g30286,g30359,II39895,g30287,g30360,II39899,g30288,g30362,II39902,g30289,g30363,II39906,g30290,g30365,II39909,g30291,
    g30366,II39913,g30292,g30368,II39916,g30293,g30369,II39919,g30294,g30370,II39922,g30295,g30371,II39926,g30296,g30373,
    II39930,g30297,g30375,II39933,g30298,g30376,II39936,g30299,g30377,II39939,g30300,g30378,II39942,g30301,g30379,II39945,
    g30302,g30380,II39948,g30303,g30381,II39951,g30304,g30382,g30383,II39976,g30245,g30408,II39982,g30305,g30412,II39985,
    g30246,g30435,II39991,g30247,g30439,II39997,g30248,g30443,II40002,g30249,g30446,II40008,g30250,g30450,II40016,g30251,
    g30456,II40021,g30252,g30459,II40027,g30253,g30463,II40032,g30254,g30466,II40039,g30255,g30471,II40044,g30256,g30474,
    II40051,g30257,g30479,II40054,g30258,g30480,II40059,g30259,g30483,II40066,g30260,g30488,II40071,g30261,g30491,II40075,
    g30262,g30493,II40078,g30263,g30494,II40083,g30264,g30497,II40086,g30265,g30498,II40091,g30266,g30501,II40098,II40101,
    II40104,II40107,II40110,II40113,II40116,II40119,II40122,II40125,II40128,II40131,II40134,II40137,II40140,II40143,II40146,II40149,
    II40152,II40155,II40158,II40161,II40164,II40167,II40170,II40173,II40176,II40179,II40182,II40185,II40188,II40191,II40194,II40197,
    II40200,II40203,II40206,II40209,II40212,II40215,II40218,II40221,II40224,II40227,II40230,II40233,II40236,II40239,II40242,II40245,
    II40248,II40251,II40254,II40257,II40260,II40263,II40266,II40269,II40272,II40275,g30567,g30403,g30568,g30402,g30569,g30406,
    g30570,g30404,g30571,g30401,g30572,g30399,g30573,g30405,g30574,g30400,g30575,II40288,g30455,g30578,II40291,g30468,
    g30579,II40294,g30470,g30580,II40297,g30482,g30581,II40300,g30485,g30582,II40303,g30487,g30583,II40307,g30500,g30585,
    II40310,g30503,g30586,II40313,g30505,g30587,II40317,g30338,g30591,II40320,g30341,g30592,II40326,g30356,g30600,II40420,
    II40423,II40426,II40429,II40432,II40435,II40438,II40441,II40444,II40447,II40450,II40453,II40456,g30668,g30722,II40459,g30669,
    g30723,II40462,g30670,g30724,II40465,g30671,g30725,II40468,g30672,g30726,II40471,g30673,g30727,II40475,g30674,g30729,
    II40478,g30675,g30730,II40481,g30676,g30731,II40484,g30677,g30732,II40487,g30678,g30733,II40490,g30679,g30734,II40495,
    g30680,g30737,II40498,g30681,g30738,II40501,g30682,g30739,II40504,g30683,g30740,II40507,g30684,g30741,II40510,g30686,
    g30742,II40515,g30687,g30745,II40518,g30688,g30746,II40521,g30689,g30747,II40524,g30690,g30748,II40527,g30691,g30749,
    II40531,g30692,g30751,II40534,g30693,g30752,II40537,g30694,g30753,II40542,g30695,g30756,g30765,g30685,II40555,g30699,
    g30767,II40565,g30700,g30769,II40568,g30701,g30770,II40578,g30702,g30772,II40581,g30703,g30773,II40584,g30704,g30774,
    II40594,g30705,g30776,II40597,g30706,g30777,II40600,g30707,g30778,II40611,g30708,g30781,II40614,g30709,g30782,II40618,
    g30566,g30784,II40634,g30792,II40637,g30793,II40640,g30794,II40643,g30795,II40647,g30797,II40651,g30799,II40654,g30800,
    II40658,g30802,II40661,g30635,g30803,II40664,g30636,g30804,II40667,g30637,g30805,II40670,g30638,g30806,II40673,g30639,
    g30807,II40676,g30640,g30808,II40679,g30641,g30809,II40682,g30642,g30810,II40685,g30643,g30811,II40688,g30644,g30812,
    II40691,g30645,g30813,II40694,g30646,g30814,II40697,g30647,g30815,II40700,g30648,g30816,II40703,g30649,g30817,II40706,
    g30650,g30818,II40709,g30651,g30819,II40712,g30652,g30820,II40715,g30653,g30821,II40718,g30654,g30822,II40721,g30655,
    g30823,II40724,g30656,g30824,II40727,g30657,g30825,II40730,g30658,g30826,II40733,g30659,g30827,II40736,g30660,g30828,
    II40739,g30661,g30829,II40742,g30662,g30830,II40745,g30663,g30831,II40748,g30664,g30832,II40751,g30665,g30833,II40754,
    g30666,g30834,II40757,g30667,g30835,II40760,II40763,II40766,II40769,II40772,II40775,II40778,II40781,II40784,II40787,II40790,
    II40793,II40796,II40799,II40802,II40805,II40808,II40811,II40814,II40817,II40820,II40823,II40826,II40829,II40832,II40835,II40838,
    II40841,II40844,II40847,II40850,II40853,II40856,II40859,II40862,II40865,II40868,II40871,II40874,II40877,II40880,II40883,II40886,
    II40889,II40892,II40895,II40898,II40901,II40904,II40907,II40910,II40913,II40916,II40919,II40922,II40925,II40928,II40931,II40934,
    II40937,II40940,II40943,II40946,II40949,II40952,II40955,II40958,II40961,II40964,II40967,II40970,II40973,II40976,II40979,II40982,
    II40985,II40988,II40991,II40994,II40997,II41024,g30928,II41035,g30796,g30937,II41038,g30798,g30938,II41041,g30801,g30939,
    II41044,II41047,II41050,II41053,g30962,g30958,g30963,g30957,g30964,g30961,g30965,g30959,g30966,g30956,g30967,g30954,
    g30968,g30960,g30969,g30955,g30971,g30970,II41090,g30972,II41093,g30973,II41096,g30974,II41099,g30975,II41102,g30976,
    II41105,g30977,II41108,g30978,II41111,g30979,II41114,II41117,II41120,II41123,II41126,II41129,II41132,II41135,II41138,g30988,
    II41141,g5630,g5649,g5650,g5658,g5676,g5677,g5678,g5687,g5688,g5696,g5709,g5710,g5711,g5728,g5729,
    g5730,g5739,g5740,g5748,g5757,g5758,g5767,g5768,g5769,g5786,g5787,g5788,g5797,g5798,g5807,g5816,
    g5817,g5826,g5827,g5828,g5845,g5846,g5847,g5863,g5872,g5873,g5882,g5883,g5884,g5910,g5919,g5920,
    g5949,g8327,g8328,g8329,g8339,g8340,g8350,g8385,g8386,g8387,g8394,g8395,g8396,g8406,g8407,g8417,
    g8431,g8432,g8433,g8437,g8438,g8439,g8446,g8447,g8448,g8458,g8459,g8463,g8464,g8465,g8466,g8467,
    g8468,g8472,g8473,g8474,g8481,g8482,g8483,g8484,g8485,g8486,g8487,g8488,g8489,g8490,g8491,g8492,
    g8493,g8497,g8498,g8499,g8500,g8501,g8502,g8503,g8504,g8505,g8506,g8507,g8508,g8509,g8510,g8511,
    g8512,g8513,g8515,g8516,g8517,g8518,g8519,g8520,g8521,g8522,g8523,g8524,g8525,g8526,g8527,g8528,
    g8529,g8531,g8532,g8534,g8535,g8536,g8537,g8538,g8539,g8540,g8541,g8542,g8543,g8544,g8545,g8546,
    g8548,g8549,g8551,g8552,g8553,g8554,g8555,g8556,g8557,g8558,g8559,g8561,g8562,g8564,g8565,g8566,
    g8567,g8570,g8572,g8573,g8576,g8601,g8612,g8613,g8621,g8625,g8626,g8631,g8635,g8636,g8650,g8654,
    g8666,g8676,g8687,g8688,g8703,g8704,g8705,g8706,g8717,g8722,g8723,g8724,g8725,g8751,g8755,g8760,
    g8761,g8762,g8774,g8778,g8783,g8784,g8797,g8801,g8816,g8841,g8842,g8861,g8868,g8869,g8892,g8899,
    g8906,g8907,g8932,g8939,g8946,g8947,g8972,g8979,g9004,g9009,g9026,g9033,g9034,g9047,g9048,g9049,
    g9056,g9057,g9061,g9062,g9063,g9064,g9065,g9066,g9073,g9074,g9075,g9076,g9077,g9078,g9079,g9080,
    g9081,g9082,g9083,g9090,g9091,g9092,g9093,g9094,g9095,g9096,g9097,g9098,g9099,g9100,g9101,g9102,
    g9103,g9104,g9105,g9106,g9107,g9108,g9109,g9110,g9111,g9112,g9113,g9114,g9115,g9116,g9117,g9118,
    g9119,g9120,g9121,g9122,g9123,g9124,g9125,g9126,g9127,g9131,g9132,g9133,g9137,g9138,g9139,g9143,
    g9145,g9241,g9301,g9302,g9319,g9364,g9365,g9366,g9367,g9382,g9383,g9400,g9438,g9439,g9440,g9441,
    g9442,g9461,g9462,g9463,g9464,g9479,g9480,g9497,g9518,g9519,g9520,g9521,g9522,g9523,g9534,g9580,
    g9581,g9582,g9583,g9584,g9603,g9604,g9605,g9606,g9621,g9622,g9630,g9631,g9632,g9633,g9634,g9635,
    II16735,II16736,g9636,g9639,g9647,g9648,g9660,g9661,g9662,g9663,g9664,g9665,g9676,g9722,g9723,g9724,
    g9725,g9726,g9745,g9746,g9747,g9748,g9759,g9760,g9761,g9762,g9763,g9764,g9765,g9766,g9773,g9774,
    g9775,g9776,g9777,g9778,g9779,g9780,g9781,II16826,II16827,g9782,g9785,g9793,g9794,g9806,g9807,g9808,
    g9809,g9810,g9811,g9822,g9868,g9869,g9870,g9871,g9872,g9887,g9888,g9889,g9890,g9891,g9892,g9893,
    g9894,g9901,g9902,g9903,g9904,g9905,g9906,g9907,g9908,g9909,g9910,g9911,g9912,g9919,g9920,g9921,
    g9922,g9923,g9924,g9925,g9926,g9927,II16930,II16931,g9928,g9931,g9939,g9940,g9952,g9953,g9954,g9955,
    g9956,g9957,g9968,g10007,g10008,g10009,g10010,g10011,g10012,g10013,g10014,g10024,g10035,g10036,g10037,g10041,
    g10042,g10043,g10044,g10045,g10046,g10047,g10048,g10055,g10056,g10057,g10058,g10059,g10060,g10061,g10062,g10063,
    g10064,g10065,g10066,g10073,g10074,g10075,g10076,g10077,g10078,g10079,g10080,g10081,II17042,II17043,g10082,g10085,
    g10093,g10094,g10101,g10102,g10103,g10104,g10105,g10106,g10107,g10108,g10112,g10113,g10114,g10115,g10116,g10117,
    g10118,g10119,g10120,g10121,g10122,g10123,g10133,g10144,g10145,g10146,g10150,g10151,g10152,g10153,g10154,g10155,
    g10156,g10157,g10164,g10165,g10166,g10167,g10168,g10169,g10170,g10171,g10172,g10173,g10174,g10175,g10182,g10183,
    g10184,II17156,g10186,g10192,g10193,g10194,g10195,g10196,g10197,g10198,g10199,g10200,g10201,g10202,g10203,g10204,
    g10205,g10206,g10207,g10208,g10209,g10210,g10211,g10212,g10213,g10217,g10218,g10219,g10220,g10221,g10222,g10223,
    g10224,g10225,g10226,g10227,g10228,g10238,g10249,g10250,g10251,g10255,g10256,g10257,g10258,g10259,g10260,g10261,
    g10262,g10269,g10270,g10271,g10272,g10279,g10280,g10281,g10282,g10283,g10284,g10285,g10286,g10287,g10288,g10289,
    g10290,g10291,g10292,g10293,g10294,g10295,g10296,g10297,g10298,g10299,g10300,g10301,g10302,g10303,g10304,g10305,
    g10306,g10307,g10308,g10309,g10310,g10311,g10312,g10313,g10314,g10315,g10319,g10320,g10321,g10322,g10323,g10324,
    g10325,g10326,g10327,g10328,g10329,g10330,g10340,g10351,g10352,g10353,g10360,g10361,g10362,g10363,g10364,g10365,
    g10366,g10367,g10368,g10369,g10370,g10371,g10372,g10373,g10374,g10375,g10376,g10377,g10378,g10379,g10380,g10381,
    g10382,g10383,g10384,g10385,g10386,g10387,g10388,g10389,g10390,g10391,g10392,g10393,g10394,g10395,g10396,g10397,
    g10398,g10399,g10400,g10401,g10402,g10403,g10404,g10405,g10406,g10407,g10408,g10412,g10413,g10414,g10415,g10422,
    g10423,g10430,g10431,g10432,g10433,g10434,g10435,g10436,g10437,g10438,g10439,g10440,g10441,g10442,g10443,g10444,
    g10445,g10446,g10447,g10448,g10449,g10450,g10451,g10452,g10453,g10454,g10455,g10456,g10457,g10458,g10459,g10460,
    g10461,g10462,g10463,g10464,g10465,g10466,g10467,g10468,g10469,g10470,g10471,g10472,g10473,g10474,g10475,g10476,
    g10477,g10478,g10479,II17429,g10485,g10492,g10493,g10494,g10495,g10496,g10497,g10498,g10499,g10506,g10507,g10508,
    g10509,g10510,g10511,g10512,g10513,g10514,g10515,g10516,g10517,g10518,g10519,g10520,g10521,g10522,g10523,g10524,
    g10525,g10526,g10527,g10528,g10529,g10530,g10531,g10532,g10533,g10534,g10535,g10536,g10537,g10538,g10539,g10540,
    g10541,g10548,g10555,g10556,g10557,g10558,g10559,g10566,g10567,g10568,g10569,g10570,g10571,g10572,g10573,g10580,
    g10581,g10582,g10583,g10584,g10585,g10586,g10587,g10588,g10589,g10590,g10591,g10592,g10593,g10594,g10595,g10596,
    g10597,g10598,g10599,g10600,g10604,g10605,g10612,g10613,g10614,g10615,g10616,g10623,g10624,g10625,g10626,g10627,
    g10628,g10629,g10630,g10637,g10638,g10639,g10640,g10641,g10642,g10643,g10644,g10645,g10650,g10651,g10652,g10659,
    g10660,g10661,g10662,g10663,g10670,g10671,g10672,g10673,g10674,g10675,g10678,g10680,g10681,g10682,g10689,g10690,
    g10691,g10692,g10693,g10704,g10707,g10709,g10710,II17599,g10724,g10727,g10729,g10745,g10748,g10764,g11347,g11420,
    g11421,g11431,g11607,g11612,g11637,g11771,g11788,g11805,g11814,g11816,g11838,g11847,g11851,g11880,g11885,g11922,
    g11926,g11966,g11967,g12012,g12069,g12070,g12128,g12129,g12186,g12273,g12274,g12307,g12330,g12331,g12353,g12376,
    g12419,g12429,g12477,g12494,g12514,g12531,g12650,II19937,II19938,g12876,g12908,II19971,II19972,g12916,g12938,II19996,
    II19997,g12945,g12966,II20021,II20022,g12974,g12989,g12990,g13000,g13009,g13010,g13023,g13031,g13032,g13042,II20100,
    g13056,II20131,II20132,g13247,g13266,g13270,g13289,g13291,g13295,g13316,g13320,g13322,g13326,g13335,g13340,g13343,
    g13345,g13355,g13360,g13365,g13368,g13385,g13390,g13395,g13477,g13479,g13480,g13481,g13483,g13484,g13485,g13486,
    g13487,g13488,g13489,g13490,g13491,g13492,g13493,g13496,g13498,g13499,g13500,g13502,g13503,g13504,g13505,g13506,
    g13513,g13515,g13516,g13517,g13527,g13609,g13619,g13623,g13625,g13631,g13634,g13636,g13642,g13643,g13645,g13646,
    g13648,g13654,g13655,g13656,g13671,g13672,g13674,g13675,g13676,g13701,g13702,g13703,g13704,g13705,g13738,g13739,
    g13740,g13755,g13787,g13788,g13789,g13790,g13796,g13815,g13816,g13818,g13824,g13833,g13834,g13835,g13837,g13839,
    g13845,g13846,g13847,g13851,g13853,g13854,g13855,g13860,g13862,g13870,g13871,g13878,g13880,g13884,g13892,g13900,
    g13902,g13904,g13905,g13913,g13914,g13933,g13941,g13943,g13944,g13952,g13953,g13969,g13970,g13989,g13997,g13998,
    g14006,g14007,g14022,g14023,g14039,g14040,g14059,g14067,g14097,g14098,g14113,g14114,g14130,g14131,g14143,g14182,
    g14212,g14213,g14228,g14229,g14297,g14327,g14328,g14336,g14419,g14690,g14724,g14752,g14767,g13245,g14773,g14884,
    g14894,g14956,g14957,g14958,g14975,g15020,g15030,g15031,g15046,g15047,g15064,g15093,g15094,g15104,g15105,g15126,
    g15127,g15142,g15143,g15160,g15171,g15172,g15173,g15178,g15196,g15197,g15218,g15219,g15234,g15235,g15243,g15244,
    g15245,g15246,g15247,g15257,g15258,g15259,g15264,g15282,g15283,g15304,g15305,g15320,g15321,g15324,g15325,g15335,
    g15336,g15337,g15338,g15339,g15349,g15350,g15351,g15356,g15374,g15375,g15388,g15389,g15391,g15392,g15402,g15403,
    g15407,g15410,g15411,g15421,g15422,g15423,g15424,g15425,g15435,g15436,g15437,g15442,g15452,g15453,g15459,g15460,
    g15470,g15475,g15476,g15486,g15487,g15491,g15494,g15495,g15505,g15506,g15507,g15508,g15509,g15519,g15520,g15526,
    g15527,g15545,g15546,g15556,g15561,g15562,g15572,g15573,g15577,g15580,g15581,g15591,g15592,g15593,g15594,g15595,
    g15604,g15605,g15623,g15624,g15634,g15639,g15640,g15650,g15651,g15658,g15666,g15670,g15671,g15680,g15681,g15699,
    g15700,g15710,g15717,g15725,g15729,g15730,g15739,g15740,g15753,g15754,g15755,g15765,g15769,g15770,II22028,g15780,
    g15781,g15793,g15801,g15802,g15817,g15828,g15829,g15840,g15852,II22136,g15902,g15998,g16003,g16004,g16008,g16009,
    g16010,g16015,g16016,g16017,g16018,g16019,g16028,g16029,g16030,g16031,g16032,g16033,g16045,g16046,g16047,g16048,
    g16049,g16050,g16051,g16052,g16066,g16067,g16068,g16069,g16070,g16071,g16072,g16073,g16074,g16089,g16100,g16101,
    g16102,g16103,g16104,g16105,g16106,g16107,g16108,g16111,g16112,g16119,g16127,g16133,g16134,g16135,g16136,g16137,
    g16138,g16139,g16140,g16141,g16153,g16158,g16159,g16160,g16161,g16162,g16163,g16170,g16178,g16182,g16183,g16184,
    g16185,g16186,g16187,g16188,g16198,g16199,g16200,g16211,g16212,g16217,g16218,g16219,g16220,g16221,g16222,g16229,
    g16237,g16238,g16239,g16240,g16241,g16242,g16251,g16252,g16253,g16262,g16263,g16264,g16265,g16276,g16277,g16282,
    g16283,g16284,g16285,g16286,g16288,g16289,g16290,g16291,g16298,g16299,g16300,g16301,g16309,g16310,g16311,g16312,
    g16321,g16322,g16323,g16324,g16335,g16336,g16342,g16343,g16344,g16345,g16347,g16348,g16349,g16350,g16356,g16357,
    g16358,g16359,g16367,g16368,g16369,g16370,g16379,g16380,g16381,g16382,g16383,g16385,g16386,g16387,g16388,g16389,
    g16390,g16391,g16392,g16393,g16394,g16400,g16401,g16402,g16403,g16411,g16413,g16414,g16415,g16416,g16417,g16418,
    g16419,g16420,g16421,g16422,g16423,g16424,g16425,g16426,g16427,g16428,g16429,g16430,g16431,g16432,g16438,g16443,
    g16444,g16445,g16447,g16448,g16449,g16450,g16451,g16452,g16453,g16454,g16455,g16456,g16457,g16458,g16459,g16460,
    g16461,g16462,g16505,g16513,g16527,g16535,g16558,g16590,g16607,g16625,g16639,g16650,g16850,g16855,g16856,g16859,
    g16864,g16865,g16879,g16894,g16907,g16908,g16909,g16923,g16938,g16939,g16953,g16964,g16966,g16967,g16968,g16969,
    g16970,g16984,g16987,g16988,g16989,g16990,g16991,g16993,g16994,g16997,g16998,g16999,g17001,g17015,g17017,g17018,
    g17021,g17022,g17023,g17028,g17031,g17045,g17047,g17048,g17055,g17056,g17062,g17065,g17079,g17081,g17082,g17084,
    g17090,g17091,g17097,g17100,g17114,g17116,g17117,g17122,g17128,g17129,g17135,g17138,g17143,g17144,g17149,g17155,
    g17156,g17161,g17166,g17167,g17172,g17176,g17181,g17182,g17193,g17268,g17301,g17339,g17352,g17353,g17381,g17382,
    g17393,g17395,g17396,g17397,g17398,g17408,g17409,g17428,g17446,g17447,g17448,g17449,g17450,g17460,g17461,g17462,
    g17463,g17464,g17474,g17475,g17485,g17486,g17506,g17508,g17509,g17510,g17526,g17527,g17528,g17529,g17530,g17540,
    g17541,g17542,g17543,g17544,g17554,g17555,g17556,g17576,g17577,g17578,g17597,g17598,g17599,g17600,g17616,g17617,
    g17618,g17619,g17620,g17630,g17631,g17632,g17633,g17634,g17635,g17636,g17652,g17653,g17654,g17673,g17674,g17675,
    g17694,g17695,g17696,g17697,g17713,g17714,g17715,g17716,g17717,g17718,g17719,g17734,g17735,g17736,g17737,g17752,
    g17753,g17754,g17773,g17774,g17775,g17794,g17795,g17796,g17797,g17798,g17812,g17813,g17814,g17824,g17835,g17836,
    g17837,g17838,g17853,g17854,g17855,g17874,g17875,g17876,g17877,g17900,g17901,g17902,g17912,g17924,g17925,g17926,
    g17936,g17947,g17948,g17949,g17950,g17965,g17966,g17967,g17989,g17990,g18011,g18012,g18013,g18023,g18035,g18036,
    g18037,g18047,g18058,g18059,g18060,g18061,g18062,g18088,g18106,g18107,g18128,g18129,g18130,g18140,g18152,g18153,
    g18154,g18164,g18165,g18169,g18204,g18222,g18223,g18244,g18245,g18246,g18256,g18311,g18329,g18330,g18333,g18404,
    II24619,g18547,II24689,g18597,II24738,g18629,II24758,g18638,g18645,g18647,g18648,g18649,g18650,g18651,g18652,g18653,
    g18654,g18655,g18665,g18666,g18667,g18668,g18688,g18689,g18690,g18717,g18718,g18753,g18982,g18990,g18994,g18997,
    g19007,g19010,g19063,g19079,g19080,g19087,g17215,g19088,g19089,g19090,g19092,g19093,g17218,g19094,g19095,II25280,
    g19097,g19099,g19100,g17220,g19101,g19102,II25291,g19104,g19106,g19107,g17223,g19108,II25300,g19109,g19111,g19112,
    II25311,g19116,g19117,g19124,g19131,g19142,g17159,g19143,g17174,g19146,g17191,g19148,g17202,g19150,g19155,g19161,
    g19166,g19228,g16662,g19236,g16935,g19241,g19248,g19252,g19254,g19260,g19267,g19282,g19284,g19285,g19289,g19303,
    g19307,g19316,g19317,g19320,g19324,g19328,g19347,g19351,g19355,g19356,g19381,g19385,g19413,g19449,g19476,g19499,
    g19520,g19531,g19540,g19541,g19544,g19545,g19547,g19548,g19549,g19551,g19552,g16829,g19553,g19554,g19555,g19557,
    g19558,g19559,g19560,g19561,g19562,g19564,g19565,g19566,g19567,g19568,g19569,g19570,g19571,g19572,g19574,g19575,
    g19576,g19584,g19585,g19586,g19587,g19588,g19589,g19590,g19591,g19592,g19593,g19594,g19597,g19598,g19599,g19600,
    g19601,g19602,g19603,g19604,g19605,g19606,g19614,g19615,g19616,g19617,g19618,g19619,g19620,g19621,g19623,g19624,
    g19625,g19626,g19627,g19628,g19629,g19630,g19631,g19632,g19633,g19634,g19635,g19636,g19637,g19638,g19639,g19647,
    g19648,g19649,g19650,g19651,g19653,g19654,g19655,g19656,g19660,g19661,g19662,g19663,g19664,g19665,g19666,g19667,
    g19668,g19669,g19670,g19671,g19672,g19673,g19674,g19675,g19676,g19677,g19678,g19679,g19687,g19688,g19691,g16841,
    g19692,g19693,g19694,g19695,g19697,g19698,g19699,g19700,g19701,g19702,g19703,g19704,g19708,g19709,g19710,g19711,
    g19712,g19713,g19714,g19715,g19716,g19717,g19718,g19719,g19720,g19721,g19722,g19723,g19724,g19726,g16847,g19727,
    g19728,g19729,g19730,g19731,g19732,g19733,g19734,g19735,g19736,g19737,g19738,g19739,g19741,g19742,g19743,g19744,
    g19745,g19746,g19747,g19748,g19752,g19753,g19754,g19755,g19756,g19757,g19758,g19759,g19760,g19761,g19764,g19765,
    g19766,g19767,g19768,g19769,g19770,g19771,g19772,g19773,g19774,g19775,g19776,g19777,g19778,g19779,g19780,g19781,
    g19782,g19784,g19785,g19786,g19787,g19788,g19789,g19790,g19791,g19795,g19796,g19797,II26240,g19799,g19802,g19803,
    g19804,g19805,g19806,g19807,g19808,g19809,g19810,g19811,g19812,g19813,g19814,g19815,g19816,g19817,g19818,g19819,
    g19820,g19821,g19822,g19823,g19824,g19826,g19827,g19828,g19829,g19836,g19837,g19839,g19840,g19841,II26282,g19842,
    II26285,g19843,g19846,g19847,g19848,g19849,g19850,g19851,g19852,g19853,g19854,g19855,g19856,g19857,g19858,g19859,
    g19860,g19861,g19862,g19863,g19864,g19868,g16498,g19869,g19870,II26311,g19871,g19872,g19873,g19874,II26317,g19875,
    II26320,g19876,g19879,g19880,g19881,g19882,g19883,g19884,g19885,g19886,g19887,g19888,g19889,g19895,g19899,g16520,
    g19900,g19901,II26348,g19902,g19903,g19904,g19905,II26354,g19906,II26357,g19907,g19910,g19911,g19912,g19913,g19914,
    g19920,g19924,g16551,g19925,g19926,II26377,g19927,g19928,g19929,g19930,II26383,g19931,g19932,g19935,g19939,g16583,
    g19940,g19941,II26396,g19942,g19943,g19944,g19949,g19952,g19953,II26416,g18553,g18491,g18431,g19970,g18354,g18276,
    g19971,g19976,II26432,g18277,g18189,g18090,g19982,g17992,g17913,g19983,II26440,g18603,g18555,g18504,g20000,g18449,
    g18369,g20001,g20006,g20011,g20012,g20013,g20014,II26464,g18370,g18296,g18206,g20020,g18109,g18024,g20021,II26472,
    g18635,g18605,g18568,g20038,g18522,g18464,g20039,g20044,g20048,g20049,g20050,g20051,g20052,g20053,II26500,g18465,
    g18389,g18313,g20062,g18225,g18141,g20063,II26508,g18644,g18637,g18618,g20080,g18586,g18537,g20081,g20084,g20085,
    g20086,g20087,g20088,g20089,g20090,g20091,g20092,II26525,g20093,II26528,g20094,II26541,g18538,g18484,g18406,g20103,
    g18332,g18257,g20104,g20106,g20107,g20108,g20109,g20110,g20111,g20112,g20113,g20114,g20115,II26558,g20116,II26561,
    g20117,II26564,g20118,II26567,g20119,g20131,g20132,g20133,g20134,g20135,g20136,g20137,g20138,g20139,g20144,g16679,
    g20145,II26590,g20146,II26593,g20147,II26596,g20148,II26599,g20149,g20156,g20157,g20158,g20159,g20160,g20161,g20162,
    II26615,g20177,g20182,g16705,g20183,II26621,g20184,II26624,g20185,II26627,g20186,II26630,g20187,g20188,g20189,g20190,
    g20191,g20192,II26639,g20197,II26645,g20211,g20216,g16736,g20217,II26651,g20218,II26654,g20219,g20220,g20221,g20222,
    II26661,g20227,II26667,g20241,g20246,g16778,g20247,g20248,g20249,II26676,g20254,II26682,g20268,g20270,g20271,g20272,
    II26690,g20277,II26695,g20280,g20282,g20283,g20284,g20285,II26708,g20291,g20293,g20294,II26726,g20307,g20309,II26745,
    g20326,g20460,g20472,g20480,g20486,g20492,g20499,g20502,g20503,g17507,g20506,g20512,g20525,g20538,g20640,g20647,
    g20665,g20809,g20826,g20836,g20840,g21049,g21067,g21068,g21077,g21078,g21085,g21086,g21091,g21092,g21097,g21098,
    g21103,g21107,g21111,g21112,g21121,g20054,g21122,g21123,g21124,g21128,g21129,II27695,g19318,g19300,g19286,g21136,
    g19271,g19261,g21137,g21138,g21140,g20095,g21141,g21142,g21143,II27711,g19262,g19414,g19386,g21152,g19357,g19334,
    g21153,g21154,g21155,II27717,g19345,g19321,g19304,g21156,g19290,g19276,g21157,g21158,g21160,g20120,g21161,g21162,
    g21163,II27733,g19277,g19451,g19416,g21172,g19389,g19368,g21173,g21174,g21175,II27739,g19379,g19348,g19325,g21176,
    g19308,g19295,g21177,g21178,g21180,g20150,g21181,g21182,g21188,II27755,g19296,g19478,g19453,g21192,g19419,g19400,
    g21193,g21194,g21195,II27761,g19411,g19382,g19352,g21196,g19329,g19313,g21197,g21198,g21203,II27772,g19314,g19501,
    g19480,g21207,g19456,g19430,g21208,g21209,g21210,g21218,g21226,g21229,g21234,g21243,g21245,g20299,g21251,g21252,
    g21254,g20318,g21259,g21260,g21262,g20337,g21267,g21268,g21270,g20357,g21276,g21277,g21283,g21284,g21290,g21291,
    g21292,g21298,g21299,g21300,g21301,g21302,g21303,g21304,g21305,g21306,g21307,g21308,g21309,g21310,g21311,g21312,
    g21313,g21314,g21315,g21319,g21320,g21321,g21322,g21323,g21324,g21325,g21326,g21328,g21329,g21330,g21334,g21335,
    g21336,g21337,g21338,g21339,g21340,g21341,g21342,g21343,g21344,g21345,g21349,g21350,g21351,g21352,g21353,g21354,
    g21355,g21356,g21357,g21360,g21361,g21362,g21363,g21367,g21368,g21369,g21370,g21371,g21372,g21373,g21374,g21375,
    g21378,g21379,g21380,g21381,g21388,g21389,g21390,g21391,g21392,g21393,g21394,g21395,g21396,g21397,g21398,g21401,
    g21402,g21403,g21410,g21411,g21412,g21413,g21414,g21418,g21419,g21420,g21421,g21422,g21423,g21424,g21425,g21428,
    g21438,g21439,g21440,g21444,g21445,g21446,g21447,g21448,g21452,g21453,g21454,g21455,g21456,g21476,g21480,g21481,
    g21482,g21486,g21487,g21488,g21489,g21490,g21494,g21497,g21517,g21521,g21522,g21523,g21527,II28068,g21553,II28096,
    g21564,II28103,g21589,g21593,II28126,g21597,II28133,g21610,g21611,g21622,II28155,g21626,II28162,g21635,g21639,g21650,
    II28181,g21654,g21658,g21666,g21670,g21681,g21687,g21695,g21699,g21707,g21723,g21731,g21735,g21749,g21757,g21758,
    g21773,g21805,g21812,g21818,g21822,g21891,g21892,g19288,g21899,g21900,g19306,g21906,g21911,g21912,g19327,g21913,
    g21920,g21925,g21926,g19354,g21931,g21938,g21990,g22004,g22015,g22020,II28582,g19141,g21133,g21116,g21104,g21095,
    g21084,II28594,g21167,g21147,g21134,g21117,g21105,g21096,II28609,g21183,g21168,g21148,g21135,g21118,g21106,g22187,
    g22196,g22201,g22202,g22206,g22207,g22208,g22211,g22214,g22215,g22220,g22223,g22224,g22228,g22229,g22235,g22238,
    g22244,g22245,g22250,g22254,g22255,g22264,g22265,g22270,g22272,g22273,g22281,g22282,g22285,g22289,g22291,g22292,
    g22305,g22309,g22311,g22312,g22333,g22337,g22340,g22358,g22363,g22383,g22398,g22483,g22515,g22516,g22517,g22526,
    g22546,g22555,g22556,g22557,g22566,g22577,g22581,g22587,g22595,g22596,g22597,g22606,g22607,g22610,g22614,g22618,
    g22624,g22632,g22633,g22634,g22637,g20841,g22638,g22643,g22646,g22650,g22654,g22660,g22665,g20920,g22666,g22667,
    g22674,g22679,g22682,g22686,g22690,g22699,g22700,g22701,g22707,g22714,g22719,g22722,g22726,g22727,g22732,g22738,
    g22745,g22754,g22759,g22764,g22770,g22788,g22793,g22798,g22804,g22830,g22835,g22841,g22842,g22869,g22874,g22906,
    g22984,g23104,g23106,g23118,g23119,g23127,g23128,g23138,g23139,g23409,g23414,g23419,g22755,g23423,g23428,g22789,
    g23432,g23434,g22831,g23440,g22870,g23451,g23458,g23462,g23467,g23471,g23476,g23483,g23484,g23494,g23496,g23510,
    g23512,g23525,g23527,g23536,g23538,g23544,g23547,g23550,g23551,g23552,g23554,g23558,g23559,g23560,g23563,g23564,
    g23565,g23567,g23571,g23572,g23573,g23577,g23578,g23579,g23582,g23583,g23584,g23586,g23590,g23591,g23592,g23593,
    g22845,g23598,g23599,g23600,g23604,g23605,g23606,g23609,g23610,g23611,g23615,g23616,g23617,g22810,g23618,g22608,
    g23622,g23623,g23624,g23625,g22880,g23630,g23631,g23632,g23636,g23637,g23638,g23639,g23643,g23659,g22784,g23664,
    g23665,g23666,g22851,g23667,g22644,g23671,g23672,g23673,g23674,g22915,g23679,g23680,g23681,g23686,g23687,g22668,
    g23689,g23693,g23709,g22826,g23714,g23715,g23716,g22886,g23717,g22680,g23721,g23722,g23723,g23724,g22940,g23726,
    g23734,g23735,g23740,g23741,g22708,g23743,g23747,g23763,g22865,g23768,g23769,g23770,g22921,g23771,g22720,g23772,
    g23776,g23777,g23778,g23789,g23790,g23795,g23796,g22739,g23798,g23802,g23818,g22900,g23820,g23822,g23824,g23825,
    g23829,g23830,g23831,g23842,g23843,g23848,g23849,g22771,g23851,g23852,g19179,g23854,g23855,g23857,g23859,g23860,
    g23864,g23865,g23866,g23877,g23878,g23886,g23888,g23889,g23891,g23893,g23894,g23898,g23899,g23900,g23904,g23907,
    g23909,g23910,g23912,g23914,g23915,g23917,g23939,g23941,g23942,g23944,g23971,g23972,g24029,g24211,g24217,g24221,
    g24224,g24229,g24236,g24241,g24246,g24247,g24253,g24256,g24427,g24429,g24431,g24432,g24433,g24435,g24436,g24437,
    g24439,g24440,g24441,g23545,g21119,g21227,g24529,g24540,g24541,g24542,g24550,g24552,g24553,g24554,g24559,g24561,
    g24563,g24564,g24565,g24569,g24571,g24573,g24574,g24578,g24580,g24585,g24590,g24591,g24595,g24596,g24603,g24604,
    g24610,g24611,g24644,g24664,g24683,g24700,g24745,g15454,g24746,g24747,g24748,g24749,g15540,g24750,g24751,g24752,
    g24754,g24755,g24757,g24758,g15618,g24759,g24760,g24761,g24762,g24767,g24768,g24769,g24772,g24773,g24774,g24775,
    g15694,g24776,g24777,g24779,g24780,g24781,g24788,g24789,g24790,g24792,g24793,g24794,g24795,g24232,g24796,g24798,
    g24799,g24802,g24803,g24804,g24809,g24810,g24811,g24813,g24818,g24821,g24822,g24824,g24825,g24826,g24831,g24100,
    g24838,g24840,g24841,g24843,g24846,g24109,g24853,g24855,g24858,g24861,g24126,g24867,g24869,g24870,g24874,g24876,
    g24145,g24878,g24881,g24882,g24884,g24885,g24888,g24898,g24899,g24901,g24902,g24905,g24906,g24907,g24908,g24921,
    g24922,g24924,g24938,g24964,g24974,g25086,g25102,g25117,g25128,g25178,g24623,g25181,g24636,g25182,g24681,g25184,
    g24694,g25187,g24633,g25188,g24652,g25192,g24711,g25193,g24653,g25196,g24672,g25198,g24691,g25269,g25277,g25278,
    g25281,g25282,g25286,g25287,g25289,g25290,g25294,g25295,g25299,g25300,g25304,g25309,g25310,g25318,g24682,g25321,
    g25075,g25328,g25334,g25337,g25342,g25346,g25348,g25351,g25356,g25360,g25362,g25365,g25371,g25375,g25377,g25388,
    g25392,g25453,g25457,g25461,g25466,g25470,g24479,g25475,g25482,g24480,g25483,g24481,g25487,g24485,g25505,g25506,
    g25513,g24487,g25514,g24488,g25518,g24489,g25552,g25553,g25560,g24494,g25561,g24495,g25565,g24496,g25618,g25619,
    g25626,g24504,g25627,g24505,g25628,g21008,g25629,g25697,g25881,g25951,g24800,g25953,g24783,g25957,g24782,g25961,
    g24770,g25963,g24756,g25968,g24871,g25972,g24859,g25973,g24847,g25975,g24606,g25977,g24845,g25978,g24836,g25980,
    g24663,g25981,g24819,g26023,g26024,g26026,g26027,g25418,g26028,g26029,g26030,g25429,g26032,g26033,g26034,g26035,
    g25523,g26036,g26038,g25589,g26039,g25668,g26040,g25745,g26051,g26052,g25941,g26053,g26054,g25944,g26060,g25943,
    g26061,g26062,g25947,g26067,g25946,g26068,g26069,g25949,g26074,g25948,g26075,g26080,g25950,g26082,g26085,g26091,
    g26157,g26158,g26163,g26166,g26171,g26186,g26188,g26207,g26212,g26213,g26231,g26233,g26234,g26235,g26236,g26243,
    g26244,g26257,g26258,g26259,g26260,g25254,g26261,g26262,g26263,g26268,g26269,g26270,g26271,g26278,g26279,g26288,
    g26289,g26290,g26291,g26292,g26293,g26298,g26299,g26300,g26301,g25258,g26302,g26303,g26307,g26309,g26310,g26311,
    g26312,g26316,g26317,g26318,g26319,g26324,g26325,g26326,g26332,g26333,g26334,g26335,g26339,g26340,g26342,g26343,
    g26344,g26345,g25261,g26346,g26347,g26348,g26350,g26351,g26352,g26353,g26357,g26361,g26362,g26363,g26365,g26366,
    g26371,g26372,g26373,g26379,g26380,g26381,g26382,g26383,g26384,g26386,g26387,g26388,g26389,g25264,g26390,g26391,
    g26392,g26396,g26397,g26400,g26404,g26405,g26406,g26408,g26409,g26414,g26415,g26416,g26422,g26423,g26424,g26425,
    g26426,g26427,g26432,g26437,g26438,g26441,g26445,g26446,g26447,g26449,g26450,g26455,g26456,g26457,g26464,g26469,
    g26470,g26473,g26477,g26478,g26479,g26488,g26493,g26494,g26504,g26663,g26668,g26673,g12431,g26674,g26754,g26755,
    g26083,g26756,g26113,g26758,g16614,g26759,g26356,g26760,g26137,g26761,g26154,g26763,g26764,g16632,g26765,g26399,
    g26766,g26767,g26087,g26768,g26440,g26769,g26770,g26059,g26771,g26773,g26145,g26774,g26472,g26775,g26099,g26777,
    g26066,g26778,g26780,g26119,g26783,g26073,g26784,g26787,g26129,g26790,g26079,g26791,g26794,g26143,g26797,g26148,
    g26829,g26833,g26842,g26845,g26851,g26853,g26860,g26866,g26955,g26958,g26961,g26962,g26963,g26965,g23320,g26966,
    g26967,g26968,g26969,g26970,g21976,g26971,g23325,g26972,g26973,g26977,g26978,g26979,g23331,g26980,g23360,g26981,
    g26982,g21983,g26984,g23335,g26985,g26986,g26993,g26994,g26995,g21991,g26996,g26997,g22050,g26998,g26999,g27000,
    g23340,g27001,g23364,g27002,g27003,g21996,g27004,g23344,g27005,g27006,g27007,g27008,g27009,g23368,g27016,g27017,
    g27018,g22005,g27019,g27020,g22069,g27021,g27022,g27023,g23349,g27024,g23372,g27025,g27026,g22009,g27027,g27028,
    g27029,g27030,g22083,g27031,g27032,g27033,g27034,g27035,g23377,g27042,g27043,g27044,g22016,g27045,g27046,g22093,
    g27047,g27048,g27049,g23353,g27050,g23381,g27052,g27053,g27054,g27055,g27056,g27057,g27058,g22108,g27059,g27060,
    g27061,g27062,g27063,g23388,g27070,g27071,g27072,g22021,g27073,g27074,g22118,g27076,g27077,g27079,g27080,g27081,
    g27082,g27083,g27084,g27085,g22134,g27086,g27087,g27088,g27089,g27090,g23395,g27091,g27092,g27093,g27095,g27096,
    g27097,g27098,g27099,g27100,g27101,g22157,g27103,g27104,g27105,g27107,g27108,g27109,g27110,g27111,g27112,g27115,
    g27178,g26110,g27181,g16570,g27182,g26151,g27185,g26126,g27187,g16594,g27240,g26905,g27241,g26934,g27242,g27244,
    g26914,g27245,g26877,g27246,g26988,g27247,g27011,g27248,g27037,g27249,g27065,g27355,g27356,g27358,g27359,g27364,
    g27365,g27370,g27371,g27372,g27394,g27396,g27407,g27409,g27425,g27427,g27446,g27448,g27495,g23945,g27509,g27516,
    g23974,g27530,g27534,g27541,g24004,g27552,g27554,g27561,g24038,g27568,g27570,g27578,g27656,g27657,g27659,g27660,
    g27661,g27666,g27671,g26885,g27673,g27679,g27680,g27681,g27719,g27496,g27720,g27481,g27721,g27579,g27723,g27464,
    g27725,g27532,g27726,g27531,g27727,g27414,g27728,g27564,g27729,g27435,g27730,g27454,g27731,g27470,g27732,g27492,
    g27733,g27513,g27734,g27538,g27737,g27558,g27770,g27772,g27773,g27774,g27775,g27779,g27783,g27790,g27904,g27908,
    g27909,g27913,g27914,g27915,g27922,g27923,g27924,g27926,g27931,g27935,g27936,g27938,g27945,g27949,g27951,g27963,
    g27968,g27970,g27984,g27985,g27991,g28008,g28009,g28015,g28027,g28028,g28035,g28036,g28042,g28050,g28051,g28057,
    g28058,g28065,g28066,g28073,g28079,g28080,g28086,g28087,g28094,g28098,g28104,g28105,g28111,g28112,g28116,g28122,
    g28123,g28127,g28171,g28176,g28188,g28193,g27573,g28319,g27855,g28320,g27854,g28322,g27937,g28323,g27838,g28324,
    g27810,g28326,g27865,g28327,g27900,g28329,g27823,g28330,g27864,g28331,g27802,g28332,g27883,g28333,g27882,g28334,
    g27842,g28335,g27814,g28336,g27896,g28337,g28002,g28338,g28029,g28339,g28059,g28340,g28088,g28373,g28376,g28378,
    g28379,g27868,g28380,g28381,g28157,g28383,g28385,g28387,g28389,g28396,g28398,g28399,g28401,g28402,g28404,g28405,
    g28407,g28408,g28411,g28412,g28416,g28422,g28423,g28424,g28426,g28427,g28428,g28429,g28430,g28431,g28433,g28434,
    g28435,g28436,g28438,g28439,g28440,g28441,g28442,g28444,g28445,g28446,g28448,g28450,g28451,g28452,g28453,g28454,
    g28456,g28457,g28459,g28460,g28462,g28463,g28464,g28465,g28466,g28468,g28469,g28471,g28472,g28474,g28475,g28476,
    g28477,g28478,g28479,g28480,g28481,g28484,g28485,g28486,g28487,g28492,g28493,g28494,g28497,g28657,g27925,g28659,
    g27917,g28660,g27916,g28662,g27911,g28663,g27906,g28664,g27997,g28665,g27827,g28666,g27980,g28667,g27964,g28669,
    g27897,g28670,g27798,g28671,g27962,g28672,g27950,g28707,g12436,g28708,g28392,g28709,g28400,g28710,g28403,g28711,
    g28415,g28712,g28406,g28713,g28410,g28714,g28394,g28715,g28414,g28716,g28449,g28717,g28461,g28718,g28473,g28719,
    g28482,g28722,g28523,g28724,g28551,g28726,g28578,g28729,g28606,g28834,g28836,g28838,g28840,g28841,g27834,g28843,
    g28844,g27850,g28846,g28847,g28848,g27875,g28849,g28850,g28851,g27892,g28852,g28853,g28854,g28880,g28881,g28892,
    g28893,g28897,g28898,g28909,g28910,g28914,g28915,g28919,g28923,g28931,g28935,g28936,g28940,g28944,g28948,g28949,
    g28958,g28962,g28966,g28970,g28971,g28986,g28996,g28997,g29022,g29130,g28397,g29174,g29031,g29175,g29009,g29176,
    g29097,g29180,g28982,g29183,g29064,g29186,g29063,g29188,g29083,g29196,g29200,g29203,g29208,g29211,g29217,g29220,
    g29225,g29229,g29232,g29233,g29234,g29235,g29236,g29238,g29239,g29240,g29241,g29242,g29243,g29248,g29251,g29252,
    g29255,g29256,g29257,g29259,g29260,g29261,g29262,g29263,g29264,g29284,g29001,g29289,g29030,g29294,g29053,g29300,
    g29072,g29302,g29026,g29310,g28978,g29312,g29049,g29320,g29088,g29321,g29008,g29323,g29068,g29329,g29096,g29330,
    g29038,g29332,g29080,g29336,g29045,g29337,g29103,g29338,g29060,g29341,g29062,g29342,g29107,g29344,g29076,g29346,
    g29087,g29411,g29090,g29464,g29465,g29466,g29265,g29467,g29340,g29468,g29343,g29469,g29345,g29470,g29347,g29471,
    g29472,g29473,g29474,g29475,g29476,g29477,g29478,g29479,g29480,g29481,g29482,g29483,g29484,g29485,g29486,g29487,
    g29488,g29489,g29490,g29502,g29518,g28728,g29520,g28731,g29521,g28733,g29522,g27735,g29523,g28737,g29524,g28739,
    g29525,g29195,g29526,g27741,g29527,g28748,g29528,g28750,g29529,g29199,g29531,g29202,g29532,g27746,g29533,g28762,
    g29534,g29206,g29536,g29207,g29538,g29210,g29539,g27754,g29540,g26041,g29541,g29214,g29543,g29215,g29545,g29216,
    g29547,g29219,g29548,g28784,g29549,g26043,g29550,g29222,g29553,g29223,g29555,g29224,g29557,g28789,g29558,g28790,
    g29559,g26045,g29560,g29227,g29562,g29228,g29564,g28794,g29565,g28795,g29566,g26047,g29567,g29231,g29572,g28802,
    g29573,g28803,g29575,g28813,g29607,g29610,g29614,g29615,g29619,g29622,g29624,g29625,g29626,g29790,g29792,g29793,
    g29810,g29748,g29811,g29703,g29812,g29762,g29813,g29760,g29814,g29728,g29815,g29727,g29816,g29759,g29817,g29709,
    g29818,g29732,g29819,g29751,g29820,g29717,g29821,g29731,g29822,g29705,g29827,g29741,g29828,g29740,g29833,g29725,
    g29834,g29713,g29839,g29747,g29909,g29735,g29910,g29779,g29942,g29771,g29944,g29782,g29945,g29773,g29946,g29778,
    g29947,g29785,g29948,g29775,g29949,g29781,g29950,g29788,g29951,g29777,g29952,g29784,g29953,g29791,g29954,g29770,
    g29955,g29787,g29956,g29780,g29957,g29772,g29958,g29783,g29959,g29774,g29960,g29786,g29961,g29776,g29962,g29789,
    g29963,g29758,g29964,g29757,g29965,g29756,g29966,g29755,g29967,g29754,g29968,g29765,g29969,g29721,g29970,g29764,
    g29971,g29763,g29980,g29981,g29982,g29983,g29984,g29985,g29986,g29987,g29988,g29989,g29990,g29991,g29992,g12441,
    g29993,g29994,g29995,g29996,g29997,g29918,g29998,g29922,g29999,g29924,g30000,g29930,g30001,g30002,g30003,g30004,
    g29926,g30005,g30006,g29928,g30007,g30008,g29919,g30009,g29929,g30077,g30079,g30080,g30081,g30082,g30083,g30085,
    g30086,g30087,g30088,g30089,g30090,g30091,g30092,g30093,g30094,g30095,g30096,g30097,g30098,g30099,g30100,g30101,
    g30102,g30103,g30104,g30105,g30106,g30107,g30108,g30109,g30110,g30111,g30112,g30113,g30114,g30115,g30116,g29921,
    g30117,g30118,g30123,g30070,g30127,g30065,g30128,g30062,g30129,g30071,g30131,g30059,g30132,g30068,g30133,g30067,
    g30138,g30069,g30216,g30217,g30218,g30219,g30220,g30221,g30222,g30223,g30224,g30225,g30226,g30227,g30327,g30330,
    g30333,g30334,g30337,g30340,g30345,g30348,g30351,g30352,g30355,g30361,g30364,g30367,g30372,g30228,g30374,g30387,
    g30388,g30389,g30390,g30391,g30392,g30393,g30394,g30395,g30396,g30397,g30398,g30407,g30409,g30410,g30411,g30436,
    g30437,g30438,g30440,g30441,g30442,g30444,g30445,g30447,g30448,g30449,g30451,g30452,g30453,g30454,g30457,g30458,
    g30460,g30461,g30462,g30464,g30465,g30467,g30469,g30472,g30473,g30475,g30476,g30477,g30478,g30481,g30484,g30486,
    g30489,g30490,g30492,g30495,g30496,g30499,g30502,g30504,g30696,g30697,g30698,g30728,g30605,g30735,g30629,g30736,
    g30584,g30743,g30610,g30744,g30609,g30750,g30593,g30754,g30614,g30755,g30632,g30757,g30601,g30758,g30613,g30759,
    g30588,g30760,g30622,g30761,g30621,g30762,g30608,g30763,g30597,g30764,g30628,g30766,g30617,g30916,g30785,g30917,
    g12446,g30918,g30780,g30919,g30786,g30920,g30787,g30921,g30791,g30922,g30788,g30923,g30789,g30924,g30783,g30925,
    g30790,g30944,g30935,g30945,g30931,g30946,g30930,g30947,g30936,g30948,g30929,g30949,g30933,g30950,g30932,g30951,
    g30934,g30953,g30952,g9144,g10778,g12377,g12407,g12886,g12926,g12955,g12984,g16539,g16571,g16595,g16615,g19181,
    g17729,g17979,g19186,g18419,g17887,g19187,g19188,g17830,g18096,g19191,g17807,g19192,g18183,g18270,g19193,g18492,
    g17998,g19194,g19195,g17942,g18212,g19200,g18346,g18424,g19201,g19202,g17919,g19203,g18290,g18363,g19204,g18556,
    g18115,g19205,g19206,g18053,g18319,g19209,g18079,g19210,g19211,g18441,g18497,g19212,g19213,g18030,g19214,g18383,
    g18458,g19215,g18606,g18231,g19216,g19221,g19222,g18195,g19223,g19224,g18514,g18561,g19225,g19226,g18147,g19227,
    g18478,g18531,II25477,g17024,g17000,g16992,g19230,g16985,g16965,g19231,g19232,g18302,g19233,g19234,g18578,g18611,
    g19235,II25495,g17158,g17137,g17115,g19240,g17083,g17050,g19242,II25500,g17058,g17030,g17016,g19243,g16995,g16986,
    g19244,g19245,g18395,g19246,g19250,II25516,g17173,g17160,g17142,g19253,g17121,g17085,g19255,II25521,g17093,g17064,
    g17046,g19256,g17019,g16996,g19257,g19263,g19264,II25549,g17190,g17175,g17165,g19266,g17148,g17123,g19268,II25554,
    g17131,g17099,g17080,g19269,g17049,g17020,g19275,g19278,g19279,II25588,g17201,g17192,g17180,g19281,g17171,g17150,
    g19283,g19294,g19297,g19298,g19312,g19315,g19333,g19450,g19477,g19500,g19503,g19521,g19522,g19532,g19542,II26429,
    g19981,II26455,g20015,II26461,g20019,II26491,g20057,II26497,g20061,II26532,g20098,II26538,g20102,II26571,g20123,g21120,
    g21139,g21159,g21179,g21244,g21253,g21261,g21269,g21501,g20522,g21536,g21540,g20542,g21572,g21576,g19067,g21605,
    g21609,g19084,g21634,g21774,g19121,g21787,II28305,g21788,g21789,g19128,II28318,g21799,g21800,g21801,II28323,g21802,
    g21803,g19135,g21806,II28330,g21807,g21808,g21809,II28335,g21810,g21811,g19138,g21813,II28341,g21814,g21815,g21816,
    II28346,g21817,g21819,II28351,g21820,g21821,g21823,II28365,g21844,II28369,g21846,II28374,g21849,II28380,g21856,g22175,
    g22190,g22199,g22205,g12451,g23319,g22385,g23688,g23742,g23797,g23850,g24239,g24244,g22317,g24245,g24252,g22342,
    g24254,g24257,g22365,g24258,g24965,g23922,g24978,g23954,g24989,g23983,g25000,g24013,g25183,g25186,g25190,g25195,
    g26320,g25852,g26367,g25873,g26410,g25885,g26451,g25890,g27738,g27743,g27751,g27756,II15167,II15168,II15169,g7855,
    II15183,II15184,II15185,g7875,II15190,II15191,II15192,g7876,II15204,II15205,II15206,g7895,II15211,II15212,II15213,g7896,
    II15237,II15238,II15239,g7922,II15244,II15245,II15246,g7923,II15276,II15277,II15278,g7970,II16879,II16880,II16881,g9883,
    II16965,II16966,II16967,g10003,II17059,II17060,II17061,g10095,II17149,II17150,II17151,g10185,II18106,II18107,II18108,g11188,
    II18113,II18114,II18115,g11189,II18190,II18191,II18192,g11262,II18197,II18198,II18199,g11263,II18204,II18205,II18206,g11264,
    II18280,II18281,II18282,g11330,II18287,II18288,II18289,g11331,II18368,II18369,II18370,g11410,II18799,II18800,II18801,g11621,
    II20031,II20032,II20033,g12988,II20048,II20049,II20050,g12999,II20429,II20430,II20431,g13348,II20465,II20466,II20467,g13370,
    II20504,II20505,II20506,g13399,II20743,II20744,II20745,g13507,g13893,g13915,g13934,g13957,g13971,g13990,g14027,g14041,
    g14060,g14118,g14132,g14233,g12780,g12819,g12857,g13401,g12898,g13286,g13313,g11622,g13332,g11643,g13375,g11660,
    II22062,II22063,II22064,g15814,g13024,g13310,g13331,g13353,g13354,g13374,g13404,II22282,II22283,II22284,II22316,II22317,
    II22318,II22630,g15978,II22631,II22632,II22705,g15661,II22706,II22707,II22884,II22885,II22886,II22900,II22901,II22902,II22917,
    II22918,II22919,II22924,II22925,II22926,II22936,II22937,II22938,II22945,II22946,II22947,II22952,II22953,II22954,II22962,II22963,
    II22964,II22972,II22973,II22974,II22981,II22982,II22983,II22988,II22989,II22990,II22998,II22999,II23000,II23008,II23009,II23010,
    II23018,II23019,II23020,II23027,II23028,II23029,II23034,II23035,II23036,II23045,II23046,II23047,II23055,II23056,II23057,II23065,
    II23066,II23067,II23074,II23075,II23076,II23082,II23083,II23084,II23093,II23094,II23095,II23103,II23104,II23105,II23113,II23114,
    II23115,II23123,II23124,II23125,II23131,II23132,II23133,II23142,II23143,II23144,II23152,II23153,II23154,II23161,II23162,II23163,
    II23171,II23172,II23173,II23179,II23180,II23181,II23190,II23191,II23192,II23198,II23199,II23200,II23207,II23208,II23209,II23217,
    II23218,II23219,II23225,II23226,II23227,II23233,II23234,II23235,II23242,II23243,II23244,II23256,II23257,II23258,II23264,II23265,
    II23266,II23277,II23278,II23279,II23806,II23807,II23808,II23878,II23879,II23880,II23893,II23894,II23895,II23941,II23942,II23943,
    II23958,II23959,II23960,II23966,II23967,II23968,II23981,II23982,II23983,II24005,II24006,II24007,II24015,II24016,II24017,II24028,
    II24029,II24030,II24036,II24037,II24038,II24053,II24054,II24055,II24061,II24062,II24063,II24076,II24077,II24078,II24091,II24092,
    II24093,II24102,II24103,II24104,II24110,II24111,II24112,II24123,II24124,II24125,II24131,II24132,II24133,II24148,II24149,II24150,
    II24156,II24157,II24158,II24178,II24179,II24180,II24186,II24187,II24188,II24194,II24195,II24196,II24205,II24206,II24207,II24213,
    II24214,II24215,II24226,II24227,II24228,II24234,II24235,II24236,II24251,II24252,II24253,II24263,II24264,II24265,II24271,II24272,
    II24273,II24278,II24279,II24280,II24290,II24291,II24292,II24298,II24299,II24300,II24306,II24307,II24308,II24317,II24318,II24319,
    II24325,II24326,II24327,II24338,II24339,II24340,II24351,II24352,II24353,II24361,II24362,II24363,II24372,II24373,II24374,II24380,
    II24381,II24382,II24387,II24388,II24389,II24399,II24400,II24401,II24407,II24408,II24409,II24415,II24416,II24417,II24426,II24427,
    II24428,II24436,II24437,II24438,II24443,II24444,II24445,II24452,II24453,II24454,II24464,II24465,II24466,II24474,II24475,II24476,
    II24485,II24486,II24487,II24493,II24494,II24495,II24500,II24501,II24502,II24512,II24513,II24514,II24520,II24521,II24522,II24530,
    II24531,II24532,II24537,II24538,II24539,II24544,II24545,II24546,II24553,II24554,II24555,II24565,II24566,II24567,II24575,II24576,
    II24577,II24586,II24587,II24588,II24594,II24595,II24596,II24601,II24602,II24603,II24611,II24612,II24613,II24624,II24625,II24626,
    II24632,II24633,II24634,II24639,II24640,II24641,II24646,II24647,II24648,II24655,II24656,II24657,II24667,II24668,II24669,II24677,
    II24678,II24679,II24694,II24695,II24696,II24702,II24703,II24704,II24709,II24710,II24711,II24716,II24717,II24718,II24725,II24726,
    II24727,II24743,II24744,II24745,II24751,II24752,II24753,II24763,II24764,II24765,II25030,II25031,II25032,II25532,II25533,II25534,
    II25539,II25540,II25541,II25560,II25561,II25562,II25571,II25572,II25573,II25578,II25579,II25580,II25595,II25596,II25597,II25605,
    II25606,II25607,II25616,II25617,II25618,II25623,II25624,II25625,II25633,II25634,II25635,II25643,II25644,II25645,II25653,II25654,
    II25655,II25664,II25665,II25666,II25671,II25672,II25673,II25681,II25682,II25683,II25690,II25691,II25692,II25700,II25701,II25702,
    II25710,II25711,II25712,II25721,II25722,II25723,II25731,II25732,II25733,II25740,II25741,II25742,II25750,II25751,II25752,II25761,
    II25762,II25763,II25771,II25772,II25773,II25781,II25782,II25783,II25790,II25791,II25792,II25800,II25801,II25802,II25809,II25810,
    II25811,II25819,II25820,II25821,II25829,II25830,II25831,II25838,II25839,II25840,II25846,II25847,II25848,II25855,II25856,II25857,
    II25865,II25866,II25867,II25880,II25881,II25882,II25888,II25889,II25890,II25897,II25898,II25899,II25913,II25914,II25915,II25921,
    II25922,II25923,II25938,II25939,II25940,g19219,II28189,II28190,II28191,g21660,II28217,II28218,II28219,g21689,II28247,II28248,
    II28249,g21725,II28271,II28272,II28273,g21751,g21848,g21850,g21855,g21857,g21858,g21859,g21860,g21862,g21863,g21864,
    g21865,g21866,g21868,g21869,g21870,g21871,g21873,g21874,g21875,g21877,g21879,g21881,g21885,g21888,g21048,g21065,
    II28726,g21887,II28727,II28728,II28741,g21890,II28742,II28743,II28753,g21893,II28754,II28755,II28765,g21901,II28766,II28767,
    g21211,g21219,g21230,g21235,g22809,g22844,g22846,g22850,g22879,g22881,g22885,g22914,g22916,g22920,g22939,g22941,
    g23066,g23051,g23080,g23070,g22999,g22174,g23096,g23083,g23013,g22189,g23113,g23099,g23029,g22198,g23046,g22204,
    g21980,g21975,g21987,g21981,g23135,g22288,g22000,g21988,g23376,g21968,g22308,g22013,g22001,g23387,g21971,g22336,
    g23394,g21973,g22361,g23402,II30790,II30791,II30792,II30868,II30869,II30870,II30952,II30953,II30954,II31035,II31036,II31037,
    g23906,g23936,g23937,g23938,g23953,g23968,g23969,g23970,g23973,g23982,g23997,g23998,g23999,g24002,g24003,g24012,
    g24027,g24028,g24034,g24036,g24037,g24046,g24052,g24054,g24056,g24057,g24058,g24065,g24067,g24069,g24070,g24071,
    g24078,g24080,g24081,g24082,g24089,g24090,g24091,g24093,II32265,II32266,II32267,II32284,II32285,II32286,II32295,II32296,
    II32297,II32308,II32309,II32310,II32323,II32324,II32325,II32333,II32334,II32335,II32345,II32346,II32347,II32355,II32356,II32357,
    II32368,II32369,II32370,II32378,II32379,II32380,II32391,II32392,II32393,II32400,II32401,II32402,II32409,II32410,II32411,II32422,
    II32423,II32424,II32430,II32431,II32432,II32443,II32444,II32445,II32451,II32452,II32453,II32460,II32461,II32462,II32468,II32469,
    II32470,II32478,II32479,II32480,II32490,II32491,II32492,II32498,II32499,II32500,II32509,II32510,II32511,II32518,II32519,II32520,
    II32526,II32527,II32528,II32538,II32539,II32540,II32546,II32547,II32548,II32559,II32560,II32561,II32567,II32568,II32569,II32575,
    II32576,II32577,II32586,II32587,II32588,II32595,II32596,II32597,II32607,II32608,II32609,II32615,II32616,II32617,II32624,II32625,
    II32626,II32633,II32634,II32635,II32645,II32646,II32647,II32659,II32660,II32661,II32668,II32669,II32670,II32677,g23823,II32678,
    II32679,II32686,II32687,II32688,II32695,g23858,II32696,II32697,II32708,g23892,II32709,II32710,II32724,g23913,II32725,II32726,
    g24517,g24530,g24543,g24555,II35020,II35021,II35022,g26859,II35034,II35035,II35036,g26865,II35042,II35043,II35044,g26867,
    II35057,II35058,II35059,g26874,g25699,g25569,g25631,g25772,g25648,g25708,g25826,g25725,g25781,g25861,g25798,g25835,
    II35123,g26107,g26096,II35124,II35125,II35701,II35702,II35703,g27379,II35714,II35715,II35716,g27382,g26989,g27012,g27038,
    g27066,II35904,g27051,II35905,II35906,II35944,g27078,II35945,II35946,II35974,g27094,II35975,II35976,II35992,g27106,II35993,
    II35994,g27415,g27436,g27455,g27471,II36256,g27527,II36257,II36258,g27801,II36270,g27549,II36271,II36272,g27809,II36289,
    g27565,II36290,II36291,g27830,II36300,II36301,II36302,II36314,g27575,II36315,II36316,g27846,II36591,g27529,II36592,II36593,
    II36666,g27551,II36667,II36668,II36731,g27567,II36732,II36733,II36779,g27577,II36780,II36781,II37295,II37296,II37297,g28384,
    II37303,II37304,II37305,g28386,II37311,II37312,II37313,g28388,II37322,II37323,II37324,g28391,II37356,g27824,g27811,II37357,
    II37358,II37813,II37814,II37815,g28842,II37822,II37823,II37824,g28845,II38378,II38379,II38380,II38810,g29303,II38811,II38812,
    II38820,g29313,II38821,II38822,II38831,g29324,II38832,II38833,II38841,g29333,II38842,II38843,II39323,II39324,II39325,g29911,
    II39331,II39332,II39333,g29913,II39339,II39340,II39341,g29915,II39347,II39348,II39349,g29917,II39359,g29766,II39360,II39361,
    g29923,II39367,g29767,II39368,II39369,g29925,II39375,g29768,II39376,II39377,g29927,II39384,g29718,g29710,II39385,II39386,
    II39391,g29769,II39392,II39393,g29931,II39532,II39533,II39534,g30034,II39539,II39540,II39541,g30035,II39689,II39690,II39691,
    II40558,II40559,II40560,g30768,II40571,II40572,II40573,g30771,II40587,II40588,II40589,g30775,II40603,II40604,II40605,g30779,
    II40627,g30602,g30594,II40628,II40629,II41010,II41011,II41012,g30926,II41017,II41018,II41019,g30927,II41064,II41065,II41066,
    g16020,g16036,g16058,g16082,g16094,g16120,g16171,g16230,g18352,g18430,g18447,g18503,g18520,g18567,g18584,g18617,
    g19160,g19165,g19171,g19177,g20878,g20895,g20914,g20938,g21083,g21618,g21646,g21677,g21706,g21738,g21762,g21778,
    g21793,g22144,g22165,g22181,g22186,g22195,g22210,g22216,g22227,g22985,g22987,g22990,g22997,g23009,g23025,g23042,
    g23061,g23386,g23393,g23401,g23408,g23427,g23433,g23461,g23477,g24227,g24234,g24242,g24249,g24428,g24486,g24490,
    g24492,g24493,g24497,g24500,g24502,g24503,g24506,g24509,g24512,g24514,g24515,g24516,g24520,g24523,g24526,g24528,
    g24533,g24536,g24546,g24558,g24566,g24575,g24613,g24622,g24624,g24637,g24638,g24656,g24657,g24675,g24708,g24717,
    g24720,g24728,g24731,g24736,g24739,g24742,g25076,g25077,g25078,g25081,g25082,g25085,g25091,g25099,g25125,g25127,
    g25129,g25208,g25216,g25226,g25238,g25273,g25311,g25426,g25962,g25967,g25974,g25979,g26042,g26044,g26046,g26049,
    g26050,g26055,g26081,g26084,g26090,g26103,g26140,g26560,g26583,g26607,g26630,g26799,g26800,g26801,g26802,g26873,
    g26882,g26891,g26901,g27175,g27179,g27184,g27188,g27250,g27251,g27252,g27254,g27478,g27501,g27521,g27546,g27629,
    g27631,g27655,g27658,g27736,g27742,g27747,g27755,g27869,g27886,g28185,g28189,g28191,g28192,g28654,g28656,g28658,
    g28661,g29126,g29127,g29128,g29129,g29399,g29403,g29406,g29409,g29736,g29744,g30618,g30625,extra0,extra1,extra2,
    extra3,extra4,extra5,extra6,extra7,extra8,extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,extra17,extra18,
    extra19;

  DFF_X1 DFF_0( .CK(CK), .Q(g2814), .D(g16475) );
  DFF_X1 DFF_1( .CK(CK), .Q(g2817), .D(g20571) );
  DFF_X1 DFF_2( .CK(CK), .Q(g2933), .D(g20588) );
  DFF_X1 DFF_3( .CK(CK), .Q(g2950), .D(g21951) );
  DFF_X2 DFF_4( .CK(CK), .Q(g2883), .D(g23315) );
  DFF_X2 DFF_5( .CK(CK), .Q(g2888), .D(g24423) );
  DFF_X2 DFF_6( .CK(CK), .Q(g2896), .D(g25175) );
  DFF_X1 DFF_7( .CK(CK), .Q(g2892), .D(g26019) );
  DFF_X1 DFF_8( .CK(CK), .Q(g2903), .D(g26747) );
  DFF_X1 DFF_9( .CK(CK), .Q(g2900), .D(g27237) );
  DFF_X1 DFF_10( .CK(CK), .Q(g2908), .D(g27715) );
  DFF_X1 DFF_11( .CK(CK), .Q(g2912), .D(g24424) );
  DFF_X1 DFF_12( .CK(CK), .Q(g2917), .D(g25174) );
  DFF_X1 DFF_13( .CK(CK), .Q(g2924), .D(g26020) );
  DFF_X1 DFF_14( .CK(CK), .Q(g2920), .D(g26746) );
  DFF_X1 DFF_15( .CK(CK), .Q(g2984), .D(g19061) );
  DFF_X1 DFF_16( .CK(CK), .Q(g2985), .D(g19060) );
  DFF_X1 DFF_17( .CK(CK), .Q(g2930), .D(g19062) );
  DFF_X1 DFF_18( .CK(CK), .Q(g2929), .D(g2930) );
  DFF_X1 DFF_19( .CK(CK), .Q(g2879), .D(g16494) );
  DFF_X1 DFF_20( .CK(CK), .Q(g2934), .D(g16476) );
  DFF_X1 DFF_21( .CK(CK), .Q(g2935), .D(g16477) );
  DFF_X1 DFF_22( .CK(CK), .Q(g2938), .D(g16478) );
  DFF_X1 DFF_23( .CK(CK), .Q(g2941), .D(g16479) );
  DFF_X1 DFF_24( .CK(CK), .Q(g2944), .D(g16480) );
  DFF_X1 DFF_25( .CK(CK), .Q(g2947), .D(g16481) );
  DFF_X1 DFF_26( .CK(CK), .Q(g2953), .D(g16482) );
  DFF_X1 DFF_27( .CK(CK), .Q(g2956), .D(g16483) );
  DFF_X1 DFF_28( .CK(CK), .Q(g2959), .D(g16484) );
  DFF_X1 DFF_29( .CK(CK), .Q(g2962), .D(g16485) );
  DFF_X1 DFF_30( .CK(CK), .Q(g2963), .D(g16486) );
  DFF_X1 DFF_31( .CK(CK), .Q(g2966), .D(g16487) );
  DFF_X1 DFF_32( .CK(CK), .Q(g2969), .D(g16488) );
  DFF_X1 DFF_33( .CK(CK), .Q(g2972), .D(g16489) );
  DFF_X1 DFF_34( .CK(CK), .Q(g2975), .D(g16490) );
  DFF_X1 DFF_35( .CK(CK), .Q(g2978), .D(g16491) );
  DFF_X1 DFF_36( .CK(CK), .Q(g2981), .D(g16492) );
  DFF_X2 DFF_37( .CK(CK), .Q(g2874), .D(g16493) );
  DFF_X2 DFF_38( .CK(CK), .Q(g1506), .D(g20572) );
  DFF_X1 DFF_39( .CK(CK), .Q(g1501), .D(g20573) );
  DFF_X1 DFF_40( .CK(CK), .Q(g1496), .D(g20574) );
  DFF_X1 DFF_41( .CK(CK), .Q(g1491), .D(g20575) );
  DFF_X1 DFF_42( .CK(CK), .Q(g1486), .D(g20576) );
  DFF_X1 DFF_43( .CK(CK), .Q(g1481), .D(g20577) );
  DFF_X1 DFF_44( .CK(CK), .Q(g1476), .D(g20578) );
  DFF_X1 DFF_45( .CK(CK), .Q(g1471), .D(g20579) );
  DFF_X1 DFF_46( .CK(CK), .Q(g2877), .D(g23313) );
  DFF_X1 DFF_47( .CK(CK), .Q(g2861), .D(g21960) );
  DFF_X1 DFF_48( .CK(CK), .Q(g813), .D(g2861) );
  DFF_X1 DFF_49( .CK(CK), .Q(g2864), .D(g21961) );
  DFF_X1 DFF_50( .CK(CK), .Q(g809), .D(g2864) );
  DFF_X1 DFF_51( .CK(CK), .Q(g2867), .D(g21962) );
  DFF_X1 DFF_52( .CK(CK), .Q(g805), .D(g2867) );
  DFF_X1 DFF_53( .CK(CK), .Q(g2870), .D(g21963) );
  DFF_X1 DFF_54( .CK(CK), .Q(g801), .D(g2870) );
  DFF_X1 DFF_55( .CK(CK), .Q(g2818), .D(g21947) );
  DFF_X1 DFF_56( .CK(CK), .Q(g797), .D(g2818) );
  DFF_X1 DFF_57( .CK(CK), .Q(g2821), .D(g21948) );
  DFF_X1 DFF_58( .CK(CK), .Q(g793), .D(g2821) );
  DFF_X1 DFF_59( .CK(CK), .Q(g2824), .D(g21949) );
  DFF_X1 DFF_60( .CK(CK), .Q(g789), .D(g2824) );
  DFF_X1 DFF_61( .CK(CK), .Q(g2827), .D(g21950) );
  DFF_X1 DFF_62( .CK(CK), .Q(g785), .D(g2827) );
  DFF_X1 DFF_63( .CK(CK), .Q(g2830), .D(g23312) );
  DFF_X1 DFF_64( .CK(CK), .Q(g2873), .D(g2830) );
  DFF_X1 DFF_65( .CK(CK), .Q(g2833), .D(g21952) );
  DFF_X1 DFF_66( .CK(CK), .Q(g125), .D(g2833) );
  DFF_X1 DFF_67( .CK(CK), .Q(g2836), .D(g21953) );
  DFF_X1 DFF_68( .CK(CK), .Q(g121), .D(g2836) );
  DFF_X1 DFF_69( .CK(CK), .Q(g2839), .D(g21954) );
  DFF_X1 DFF_70( .CK(CK), .Q(g117), .D(g2839) );
  DFF_X1 DFF_71( .CK(CK), .Q(g2842), .D(g21955) );
  DFF_X1 DFF_72( .CK(CK), .Q(g113), .D(g2842) );
  DFF_X1 DFF_73( .CK(CK), .Q(g2845), .D(g21956) );
  DFF_X1 DFF_74( .CK(CK), .Q(g109), .D(g2845) );
  DFF_X1 DFF_75( .CK(CK), .Q(g2848), .D(g21957) );
  DFF_X1 DFF_76( .CK(CK), .Q(g105), .D(g2848) );
  DFF_X1 DFF_77( .CK(CK), .Q(g2851), .D(g21958) );
  DFF_X1 DFF_78( .CK(CK), .Q(g101), .D(g2851) );
  DFF_X1 DFF_79( .CK(CK), .Q(g2854), .D(g21959) );
  DFF_X1 DFF_80( .CK(CK), .Q(g97), .D(g2854) );
  DFF_X1 DFF_81( .CK(CK), .Q(g2858), .D(g23316) );
  DFF_X1 DFF_82( .CK(CK), .Q(g2857), .D(g2858) );
  DFF_X1 DFF_83( .CK(CK), .Q(g2200), .D(g20587) );
  DFF_X2 DFF_84( .CK(CK), .Q(g2195), .D(g20585) );
  DFF_X2 DFF_85( .CK(CK), .Q(g2190), .D(g20586) );
  DFF_X2 DFF_86( .CK(CK), .Q(g2185), .D(g20584) );
  DFF_X1 DFF_87( .CK(CK), .Q(g2180), .D(g20583) );
  DFF_X1 DFF_88( .CK(CK), .Q(g2175), .D(g20582) );
  DFF_X1 DFF_89( .CK(CK), .Q(g2170), .D(g20581) );
  DFF_X1 DFF_90( .CK(CK), .Q(g2165), .D(g20580) );
  DFF_X1 DFF_91( .CK(CK), .Q(g2878), .D(g23314) );
  DFF_X1 DFF_92( .CK(CK), .Q(g3129), .D(g13475) );
  DFF_X1 DFF_93( .CK(CK), .Q(g3117), .D(g3129) );
  DFF_X1 DFF_94( .CK(CK), .Q(g3109), .D(g3117) );
  DFF_X1 DFF_95( .CK(CK), .Q(g3210), .D(g20630) );
  DFF_X1 DFF_96( .CK(CK), .Q(g3211), .D(g20631) );
  DFF_X1 DFF_97( .CK(CK), .Q(g3084), .D(g20632) );
  DFF_X1 DFF_98( .CK(CK), .Q(g3085), .D(g20609) );
  DFF_X1 DFF_99( .CK(CK), .Q(g3086), .D(g20610) );
  DFF_X1 DFF_100( .CK(CK), .Q(g3087), .D(g20611) );
  DFF_X1 DFF_101( .CK(CK), .Q(g3091), .D(g20612) );
  DFF_X1 DFF_102( .CK(CK), .Q(g3092), .D(g20613) );
  DFF_X1 DFF_103( .CK(CK), .Q(g3093), .D(g20614) );
  DFF_X1 DFF_104( .CK(CK), .Q(g3094), .D(g20615) );
  DFF_X1 DFF_105( .CK(CK), .Q(g3095), .D(g20616) );
  DFF_X1 DFF_106( .CK(CK), .Q(g3096), .D(g20617) );
  DFF_X1 DFF_107( .CK(CK), .Q(g3097), .D(g26751) );
  DFF_X2 DFF_108( .CK(CK), .Q(g3098), .D(g26752) );
  DFF_X2 DFF_109( .CK(CK), .Q(g3099), .D(g26753) );
  DFF_X1 DFF_110( .CK(CK), .Q(g3100), .D(g29163) );
  DFF_X1 DFF_111( .CK(CK), .Q(g3101), .D(g29164) );
  DFF_X1 DFF_112( .CK(CK), .Q(g3102), .D(g29165) );
  DFF_X1 DFF_113( .CK(CK), .Q(g3103), .D(g30120) );
  DFF_X1 DFF_114( .CK(CK), .Q(g3104), .D(g30121) );
  DFF_X1 DFF_115( .CK(CK), .Q(g3105), .D(g30122) );
  DFF_X1 DFF_116( .CK(CK), .Q(g3106), .D(g30941) );
  DFF_X1 DFF_117( .CK(CK), .Q(g3107), .D(g30942) );
  DFF_X1 DFF_118( .CK(CK), .Q(g3108), .D(g30943) );
  DFF_X1 DFF_119( .CK(CK), .Q(g3155), .D(g20618) );
  DFF_X1 DFF_120( .CK(CK), .Q(g3158), .D(g20619) );
  DFF_X1 DFF_121( .CK(CK), .Q(g3161), .D(g20620) );
  DFF_X1 DFF_122( .CK(CK), .Q(g3164), .D(g20621) );
  DFF_X1 DFF_123( .CK(CK), .Q(g3167), .D(g20622) );
  DFF_X1 DFF_124( .CK(CK), .Q(g3170), .D(g20623) );
  DFF_X1 DFF_125( .CK(CK), .Q(g3173), .D(g20624) );
  DFF_X1 DFF_126( .CK(CK), .Q(g3176), .D(g20625) );
  DFF_X1 DFF_127( .CK(CK), .Q(g3179), .D(g20626) );
  DFF_X1 DFF_128( .CK(CK), .Q(g3182), .D(g20627) );
  DFF_X1 DFF_129( .CK(CK), .Q(g3185), .D(g20628) );
  DFF_X1 DFF_130( .CK(CK), .Q(g3088), .D(g20629) );
  DFF_X1 DFF_131( .CK(CK), .Q(g3191), .D(g27717) );
  DFF_X1 DFF_132( .CK(CK), .Q(g3194), .D(g28316) );
  DFF_X2 DFF_133( .CK(CK), .Q(g3197), .D(g28317) );
  DFF_X2 DFF_134( .CK(CK), .Q(g3198), .D(g28318) );
  DFF_X1 DFF_135( .CK(CK), .Q(g3201), .D(g28704) );
  DFF_X1 DFF_136( .CK(CK), .Q(g3204), .D(g28705) );
  DFF_X1 DFF_137( .CK(CK), .Q(g3207), .D(g28706) );
  DFF_X1 DFF_138( .CK(CK), .Q(g3188), .D(g29463) );
  DFF_X1 DFF_139( .CK(CK), .Q(g3133), .D(g29656) );
  DFF_X1 DFF_140( .CK(CK), .Q(g3132), .D(g28698) );
  DFF_X1 DFF_141( .CK(CK), .Q(g3128), .D(g29166) );
  DFF_X1 DFF_142( .CK(CK), .Q(g3127), .D(g28697) );
  DFF_X1 DFF_143( .CK(CK), .Q(g3126), .D(g28315) );
  DFF_X1 DFF_144( .CK(CK), .Q(g3125), .D(g28696) );
  DFF_X1 DFF_145( .CK(CK), .Q(g3124), .D(g28314) );
  DFF_X1 DFF_146( .CK(CK), .Q(g3123), .D(g28313) );
  DFF_X1 DFF_147( .CK(CK), .Q(g3120), .D(g28695) );
  DFF_X1 DFF_148( .CK(CK), .Q(g3114), .D(g28694) );
  DFF_X1 DFF_149( .CK(CK), .Q(g3113), .D(g28693) );
  DFF_X1 DFF_150( .CK(CK), .Q(g3112), .D(g28312) );
  DFF_X1 DFF_151( .CK(CK), .Q(g3110), .D(g28311) );
  DFF_X1 DFF_152( .CK(CK), .Q(g3111), .D(g28310) );
  DFF_X1 DFF_153( .CK(CK), .Q(g3139), .D(g29461) );
  DFF_X1 DFF_154( .CK(CK), .Q(g3136), .D(g28701) );
  DFF_X1 DFF_155( .CK(CK), .Q(g3134), .D(g28700) );
  DFF_X1 DFF_156( .CK(CK), .Q(g3135), .D(g28699) );
  DFF_X1 DFF_157( .CK(CK), .Q(g3151), .D(g29462) );
  DFF_X1 DFF_158( .CK(CK), .Q(g3142), .D(g28703) );
  DFF_X1 DFF_159( .CK(CK), .Q(g3147), .D(g28702) );
  DFF_X1 DFF_160( .CK(CK), .Q(g185), .D(g29657) );
  DFF_X2 DFF_161( .CK(CK), .Q(g138), .D(g13405) );
  DFF_X1 DFF_162( .CK(CK), .Q(g135), .D(g138) );
  DFF_X1 DFF_163( .CK(CK), .Q(g165), .D(g135) );
  DFF_X1 DFF_164( .CK(CK), .Q(g130), .D(g24259) );
  DFF_X1 DFF_165( .CK(CK), .Q(g131), .D(g24260) );
  DFF_X1 DFF_166( .CK(CK), .Q(g129), .D(g24261) );
  DFF_X1 DFF_167( .CK(CK), .Q(g133), .D(g24262) );
  DFF_X1 DFF_168( .CK(CK), .Q(g134), .D(g24263) );
  DFF_X1 DFF_169( .CK(CK), .Q(g132), .D(g24264) );
  DFF_X1 DFF_170( .CK(CK), .Q(g142), .D(g24265) );
  DFF_X1 DFF_171( .CK(CK), .Q(g143), .D(g24266) );
  DFF_X1 DFF_172( .CK(CK), .Q(g141), .D(g24267) );
  DFF_X1 DFF_173( .CK(CK), .Q(g145), .D(g24268) );
  DFF_X1 DFF_174( .CK(CK), .Q(g146), .D(g24269) );
  DFF_X1 DFF_175( .CK(CK), .Q(g144), .D(g24270) );
  DFF_X1 DFF_176( .CK(CK), .Q(g148), .D(g24271) );
  DFF_X1 DFF_177( .CK(CK), .Q(g149), .D(g24272) );
  DFF_X1 DFF_178( .CK(CK), .Q(g147), .D(g24273) );
  DFF_X1 DFF_179( .CK(CK), .Q(g151), .D(g24274) );
  DFF_X1 DFF_180( .CK(CK), .Q(g152), .D(g24275) );
  DFF_X1 DFF_181( .CK(CK), .Q(g150), .D(g24276) );
  DFF_X1 DFF_182( .CK(CK), .Q(g154), .D(g24277) );
  DFF_X1 DFF_183( .CK(CK), .Q(g155), .D(g24278) );
  DFF_X1 DFF_184( .CK(CK), .Q(g153), .D(g24279) );
  DFF_X1 DFF_185( .CK(CK), .Q(g157), .D(g24280) );
  DFF_X1 DFF_186( .CK(CK), .Q(g158), .D(g24281) );
  DFF_X1 DFF_187( .CK(CK), .Q(g156), .D(g24282) );
  DFF_X1 DFF_188( .CK(CK), .Q(g160), .D(g24283) );
  DFF_X1 DFF_189( .CK(CK), .Q(g161), .D(g24284) );
  DFF_X1 DFF_190( .CK(CK), .Q(g159), .D(g24285) );
  DFF_X2 DFF_191( .CK(CK), .Q(g163), .D(g24286) );
  DFF_X2 DFF_192( .CK(CK), .Q(g164), .D(g24287) );
  DFF_X1 DFF_193( .CK(CK), .Q(g162), .D(g24288) );
  DFF_X1 DFF_194( .CK(CK), .Q(g169), .D(g26679) );
  DFF_X1 DFF_195( .CK(CK), .Q(g170), .D(g26680) );
  DFF_X1 DFF_196( .CK(CK), .Q(g168), .D(g26681) );
  DFF_X1 DFF_197( .CK(CK), .Q(g172), .D(g26682) );
  DFF_X1 DFF_198( .CK(CK), .Q(g173), .D(g26683) );
  DFF_X1 DFF_199( .CK(CK), .Q(g171), .D(g26684) );
  DFF_X1 DFF_200( .CK(CK), .Q(g175), .D(g26685) );
  DFF_X1 DFF_201( .CK(CK), .Q(g176), .D(g26686) );
  DFF_X1 DFF_202( .CK(CK), .Q(g174), .D(g26687) );
  DFF_X1 DFF_203( .CK(CK), .Q(g178), .D(g26688) );
  DFF_X1 DFF_204( .CK(CK), .Q(g179), .D(g26689) );
  DFF_X1 DFF_205( .CK(CK), .Q(g177), .D(g26690) );
  DFF_X1 DFF_206( .CK(CK), .Q(g186), .D(g30506) );
  DFF_X1 DFF_207( .CK(CK), .Q(g189), .D(g30507) );
  DFF_X1 DFF_208( .CK(CK), .Q(g192), .D(g30508) );
  DFF_X1 DFF_209( .CK(CK), .Q(g231), .D(g30842) );
  DFF_X1 DFF_210( .CK(CK), .Q(g234), .D(g30843) );
  DFF_X1 DFF_211( .CK(CK), .Q(g237), .D(g30844) );
  DFF_X1 DFF_212( .CK(CK), .Q(g195), .D(g30836) );
  DFF_X1 DFF_213( .CK(CK), .Q(g198), .D(g30837) );
  DFF_X1 DFF_214( .CK(CK), .Q(g201), .D(g30838) );
  DFF_X1 DFF_215( .CK(CK), .Q(g240), .D(g30845) );
  DFF_X1 DFF_216( .CK(CK), .Q(g243), .D(g30846) );
  DFF_X1 DFF_217( .CK(CK), .Q(g246), .D(g30847) );
  DFF_X1 DFF_218( .CK(CK), .Q(g204), .D(g30509) );
  DFF_X1 DFF_219( .CK(CK), .Q(g207), .D(g30510) );
  DFF_X1 DFF_220( .CK(CK), .Q(g210), .D(g30511) );
  DFF_X1 DFF_221( .CK(CK), .Q(g249), .D(g30515) );
  DFF_X1 DFF_222( .CK(CK), .Q(g252), .D(g30516) );
  DFF_X1 DFF_223( .CK(CK), .Q(g255), .D(g30517) );
  DFF_X1 DFF_224( .CK(CK), .Q(g213), .D(g30512) );
  DFF_X1 DFF_225( .CK(CK), .Q(g216), .D(g30513) );
  DFF_X1 DFF_226( .CK(CK), .Q(g219), .D(g30514) );
  DFF_X2 DFF_227( .CK(CK), .Q(g258), .D(g30518) );
  DFF_X1 DFF_228( .CK(CK), .Q(g261), .D(g30519) );
  DFF_X1 DFF_229( .CK(CK), .Q(g264), .D(g30520) );
  DFF_X1 DFF_230( .CK(CK), .Q(g222), .D(g30839) );
  DFF_X1 DFF_231( .CK(CK), .Q(g225), .D(g30840) );
  DFF_X1 DFF_232( .CK(CK), .Q(g228), .D(g30841) );
  DFF_X1 DFF_233( .CK(CK), .Q(g267), .D(g30848) );
  DFF_X1 DFF_234( .CK(CK), .Q(g270), .D(g30849) );
  DFF_X1 DFF_235( .CK(CK), .Q(g273), .D(g30850) );
  DFF_X1 DFF_236( .CK(CK), .Q(g92), .D(g25983) );
  DFF_X1 DFF_237( .CK(CK), .Q(g88), .D(g26678) );
  DFF_X1 DFF_238( .CK(CK), .Q(g83), .D(g27189) );
  DFF_X1 DFF_239( .CK(CK), .Q(g79), .D(g27683) );
  DFF_X1 DFF_240( .CK(CK), .Q(g74), .D(g28206) );
  DFF_X1 DFF_241( .CK(CK), .Q(g70), .D(g28673) );
  DFF_X1 DFF_242( .CK(CK), .Q(g65), .D(g29131) );
  DFF_X1 DFF_243( .CK(CK), .Q(g61), .D(g29413) );
  DFF_X1 DFF_244( .CK(CK), .Q(g56), .D(g29627) );
  DFF_X1 DFF_245( .CK(CK), .Q(g52), .D(g29794) );
  DFF_X1 DFF_246( .CK(CK), .Q(g180), .D(g20555) );
  DFF_X1 DFF_247( .CK(CK), .Q(g182), .D(g180) );
  DFF_X1 DFF_248( .CK(CK), .Q(g181), .D(g182) );
  DFF_X1 DFF_249( .CK(CK), .Q(g276), .D(g13406) );
  DFF_X1 DFF_250( .CK(CK), .Q(g405), .D(g276) );
  DFF_X1 DFF_251( .CK(CK), .Q(g401), .D(g405) );
  DFF_X1 DFF_252( .CK(CK), .Q(g309), .D(g11496) );
  DFF_X1 DFF_253( .CK(CK), .Q(g354), .D(g28207) );
  DFF_X1 DFF_254( .CK(CK), .Q(g343), .D(g28208) );
  DFF_X1 DFF_255( .CK(CK), .Q(g346), .D(g28209) );
  DFF_X1 DFF_256( .CK(CK), .Q(g369), .D(g28210) );
  DFF_X1 DFF_257( .CK(CK), .Q(g358), .D(g28211) );
  DFF_X1 DFF_258( .CK(CK), .Q(g361), .D(g28212) );
  DFF_X1 DFF_259( .CK(CK), .Q(g384), .D(g28213) );
  DFF_X1 DFF_260( .CK(CK), .Q(g373), .D(g28214) );
  DFF_X2 DFF_261( .CK(CK), .Q(g376), .D(g28215) );
  DFF_X2 DFF_262( .CK(CK), .Q(g398), .D(g28216) );
  DFF_X1 DFF_263( .CK(CK), .Q(g388), .D(g28217) );
  DFF_X1 DFF_264( .CK(CK), .Q(g391), .D(g28218) );
  DFF_X1 DFF_265( .CK(CK), .Q(g408), .D(g29414) );
  DFF_X1 DFF_266( .CK(CK), .Q(g411), .D(g29415) );
  DFF_X1 DFF_267( .CK(CK), .Q(g414), .D(g29416) );
  DFF_X1 DFF_268( .CK(CK), .Q(g417), .D(g29631) );
  DFF_X1 DFF_269( .CK(CK), .Q(g420), .D(g29632) );
  DFF_X1 DFF_270( .CK(CK), .Q(g423), .D(g29633) );
  DFF_X1 DFF_271( .CK(CK), .Q(g427), .D(g29417) );
  DFF_X1 DFF_272( .CK(CK), .Q(g428), .D(g29418) );
  DFF_X1 DFF_273( .CK(CK), .Q(g426), .D(g29419) );
  DFF_X1 DFF_274( .CK(CK), .Q(g429), .D(g27684) );
  DFF_X1 DFF_275( .CK(CK), .Q(g432), .D(g27685) );
  DFF_X1 DFF_276( .CK(CK), .Q(g435), .D(g27686) );
  DFF_X1 DFF_277( .CK(CK), .Q(g438), .D(g27687) );
  DFF_X1 DFF_278( .CK(CK), .Q(g441), .D(g27688) );
  DFF_X1 DFF_279( .CK(CK), .Q(g444), .D(g27689) );
  DFF_X1 DFF_280( .CK(CK), .Q(g448), .D(g28674) );
  DFF_X1 DFF_281( .CK(CK), .Q(g449), .D(g28675) );
  DFF_X1 DFF_282( .CK(CK), .Q(g447), .D(g28676) );
  DFF_X1 DFF_283( .CK(CK), .Q(g312), .D(g29795) );
  DFF_X1 DFF_284( .CK(CK), .Q(g313), .D(g29796) );
  DFF_X1 DFF_285( .CK(CK), .Q(g314), .D(g29797) );
  DFF_X1 DFF_286( .CK(CK), .Q(g315), .D(g30851) );
  DFF_X1 DFF_287( .CK(CK), .Q(g316), .D(g30852) );
  DFF_X1 DFF_288( .CK(CK), .Q(g317), .D(g30853) );
  DFF_X1 DFF_289( .CK(CK), .Q(g318), .D(g30710) );
  DFF_X1 DFF_290( .CK(CK), .Q(g319), .D(g30711) );
  DFF_X1 DFF_291( .CK(CK), .Q(g320), .D(g30712) );
  DFF_X1 DFF_292( .CK(CK), .Q(g322), .D(g29628) );
  DFF_X1 DFF_293( .CK(CK), .Q(g323), .D(g29629) );
  DFF_X1 DFF_294( .CK(CK), .Q(g321), .D(g29630) );
  DFF_X1 DFF_295( .CK(CK), .Q(g403), .D(g27191) );
  DFF_X1 DFF_296( .CK(CK), .Q(g404), .D(g27192) );
  DFF_X1 DFF_297( .CK(CK), .Q(g402), .D(g27193) );
  DFF_X1 DFF_298( .CK(CK), .Q(g450), .D(g11509) );
  DFF_X1 DFF_299( .CK(CK), .Q(g451), .D(g450) );
  DFF_X1 DFF_300( .CK(CK), .Q(g452), .D(g11510) );
  DFF_X1 DFF_301( .CK(CK), .Q(g453), .D(g452) );
  DFF_X1 DFF_302( .CK(CK), .Q(g454), .D(g11511) );
  DFF_X1 DFF_303( .CK(CK), .Q(g279), .D(g454) );
  DFF_X1 DFF_304( .CK(CK), .Q(g280), .D(g11491) );
  DFF_X1 DFF_305( .CK(CK), .Q(g281), .D(g280) );
  DFF_X1 DFF_306( .CK(CK), .Q(g282), .D(g11492) );
  DFF_X1 DFF_307( .CK(CK), .Q(g283), .D(g282) );
  DFF_X1 DFF_308( .CK(CK), .Q(g284), .D(g11493) );
  DFF_X1 DFF_309( .CK(CK), .Q(g285), .D(g284) );
  DFF_X1 DFF_310( .CK(CK), .Q(g286), .D(g11494) );
  DFF_X1 DFF_311( .CK(CK), .Q(g287), .D(g286) );
  DFF_X1 DFF_312( .CK(CK), .Q(g288), .D(g11495) );
  DFF_X1 DFF_313( .CK(CK), .Q(g289), .D(g288) );
  DFF_X1 DFF_314( .CK(CK), .Q(g290), .D(g13407) );
  DFF_X1 DFF_315( .CK(CK), .Q(g291), .D(g290) );
  DFF_X1 DFF_316( .CK(CK), .Q(g299), .D(g19012) );
  DFF_X1 DFF_317( .CK(CK), .Q(g305), .D(g23148) );
  DFF_X1 DFF_318( .CK(CK), .Q(g308), .D(g23149) );
  DFF_X1 DFF_319( .CK(CK), .Q(g297), .D(g23150) );
  DFF_X1 DFF_320( .CK(CK), .Q(g296), .D(g23151) );
  DFF_X1 DFF_321( .CK(CK), .Q(g295), .D(g23152) );
  DFF_X1 DFF_322( .CK(CK), .Q(g294), .D(g23153) );
  DFF_X1 DFF_323( .CK(CK), .Q(g304), .D(g19016) );
  DFF_X1 DFF_324( .CK(CK), .Q(g303), .D(g19015) );
  DFF_X1 DFF_325( .CK(CK), .Q(g302), .D(g19014) );
  DFF_X1 DFF_326( .CK(CK), .Q(g301), .D(g19013) );
  DFF_X1 DFF_327( .CK(CK), .Q(g300), .D(g25130) );
  DFF_X1 DFF_328( .CK(CK), .Q(g298), .D(g27190) );
  DFF_X1 DFF_329( .CK(CK), .Q(g342), .D(g11497) );
  DFF_X1 DFF_330( .CK(CK), .Q(g349), .D(g342) );
  DFF_X1 DFF_331( .CK(CK), .Q(g350), .D(g11498) );
  DFF_X1 DFF_332( .CK(CK), .Q(g351), .D(g350) );
  DFF_X1 DFF_333( .CK(CK), .Q(g352), .D(g11499) );
  DFF_X1 DFF_334( .CK(CK), .Q(g353), .D(g352) );
  DFF_X1 DFF_335( .CK(CK), .Q(g357), .D(g11500) );
  DFF_X2 DFF_336( .CK(CK), .Q(g364), .D(g357) );
  DFF_X1 DFF_337( .CK(CK), .Q(g365), .D(g11501) );
  DFF_X1 DFF_338( .CK(CK), .Q(g366), .D(g365) );
  DFF_X1 DFF_339( .CK(CK), .Q(g367), .D(g11502) );
  DFF_X1 DFF_340( .CK(CK), .Q(g368), .D(g367) );
  DFF_X1 DFF_341( .CK(CK), .Q(g372), .D(g11503) );
  DFF_X1 DFF_342( .CK(CK), .Q(g379), .D(g372) );
  DFF_X2 DFF_343( .CK(CK), .Q(g380), .D(g11504) );
  DFF_X1 DFF_344( .CK(CK), .Q(g381), .D(g380) );
  DFF_X1 DFF_345( .CK(CK), .Q(g382), .D(g11505) );
  DFF_X1 DFF_346( .CK(CK), .Q(g383), .D(g382) );
  DFF_X1 DFF_347( .CK(CK), .Q(g387), .D(g11506) );
  DFF_X1 DFF_348( .CK(CK), .Q(g394), .D(g387) );
  DFF_X1 DFF_349( .CK(CK), .Q(g395), .D(g11507) );
  DFF_X1 DFF_350( .CK(CK), .Q(g396), .D(g395) );
  DFF_X1 DFF_351( .CK(CK), .Q(g397), .D(g11508) );
  DFF_X1 DFF_352( .CK(CK), .Q(g324), .D(g397) );
  DFF_X1 DFF_353( .CK(CK), .Q(g325), .D(g13408) );
  DFF_X1 DFF_354( .CK(CK), .Q(g331), .D(g325) );
  DFF_X1 DFF_355( .CK(CK), .Q(g337), .D(g331) );
  DFF_X1 DFF_356( .CK(CK), .Q(g545), .D(g13419) );
  DFF_X1 DFF_357( .CK(CK), .Q(g551), .D(g545) );
  DFF_X1 DFF_358( .CK(CK), .Q(g550), .D(g551) );
  DFF_X1 DFF_359( .CK(CK), .Q(g554), .D(g23160) );
  DFF_X1 DFF_360( .CK(CK), .Q(g557), .D(g20556) );
  DFF_X1 DFF_361( .CK(CK), .Q(g510), .D(g20557) );
  DFF_X1 DFF_362( .CK(CK), .Q(g513), .D(g16467) );
  DFF_X2 DFF_363( .CK(CK), .Q(g523), .D(g513) );
  DFF_X1 DFF_364( .CK(CK), .Q(g524), .D(g523) );
  DFF_X1 DFF_365( .CK(CK), .Q(g564), .D(g11512) );
  DFF_X1 DFF_366( .CK(CK), .Q(g569), .D(g564) );
  DFF_X1 DFF_367( .CK(CK), .Q(g570), .D(g11515) );
  DFF_X1 DFF_368( .CK(CK), .Q(g571), .D(g570) );
  DFF_X1 DFF_369( .CK(CK), .Q(g572), .D(g11516) );
  DFF_X1 DFF_370( .CK(CK), .Q(g573), .D(g572) );
  DFF_X1 DFF_371( .CK(CK), .Q(g574), .D(g11517) );
  DFF_X1 DFF_372( .CK(CK), .Q(g565), .D(g574) );
  DFF_X1 DFF_373( .CK(CK), .Q(g566), .D(g11513) );
  DFF_X1 DFF_374( .CK(CK), .Q(g567), .D(g566) );
  DFF_X1 DFF_375( .CK(CK), .Q(g568), .D(g11514) );
  DFF_X1 DFF_376( .CK(CK), .Q(g489), .D(g568) );
  DFF_X1 DFF_377( .CK(CK), .Q(g474), .D(g13409) );
  DFF_X1 DFF_378( .CK(CK), .Q(g481), .D(g474) );
  DFF_X1 DFF_379( .CK(CK), .Q(g485), .D(g481) );
  DFF_X1 DFF_380( .CK(CK), .Q(g486), .D(g24292) );
  DFF_X1 DFF_381( .CK(CK), .Q(g487), .D(g24293) );
  DFF_X1 DFF_382( .CK(CK), .Q(g488), .D(g24294) );
  DFF_X1 DFF_383( .CK(CK), .Q(g455), .D(g25139) );
  DFF_X1 DFF_384( .CK(CK), .Q(g458), .D(g25131) );
  DFF_X1 DFF_385( .CK(CK), .Q(g461), .D(g25132) );
  DFF_X1 DFF_386( .CK(CK), .Q(g477), .D(g25136) );
  DFF_X1 DFF_387( .CK(CK), .Q(g478), .D(g25137) );
  DFF_X1 DFF_388( .CK(CK), .Q(g479), .D(g25138) );
  DFF_X1 DFF_389( .CK(CK), .Q(g480), .D(g24289) );
  DFF_X1 DFF_390( .CK(CK), .Q(g484), .D(g24290) );
  DFF_X1 DFF_391( .CK(CK), .Q(g464), .D(g24291) );
  DFF_X1 DFF_392( .CK(CK), .Q(g465), .D(g25133) );
  DFF_X1 DFF_393( .CK(CK), .Q(g468), .D(g25134) );
  DFF_X1 DFF_394( .CK(CK), .Q(g471), .D(g25135) );
  DFF_X1 DFF_395( .CK(CK), .Q(g528), .D(g16468) );
  DFF_X1 DFF_396( .CK(CK), .Q(g535), .D(g528) );
  DFF_X1 DFF_397( .CK(CK), .Q(g542), .D(g535) );
  DFF_X1 DFF_398( .CK(CK), .Q(g543), .D(g19021) );
  DFF_X1 DFF_399( .CK(CK), .Q(g544), .D(g543) );
  DFF_X1 DFF_400( .CK(CK), .Q(g548), .D(g23159) );
  DFF_X1 DFF_401( .CK(CK), .Q(g549), .D(g19022) );
  DFF_X1 DFF_402( .CK(CK), .Q(g499), .D(g549) );
  DFF_X2 DFF_403( .CK(CK), .Q(g558), .D(g19023) );
  DFF_X1 DFF_404( .CK(CK), .Q(g559), .D(g558) );
  DFF_X1 DFF_405( .CK(CK), .Q(g576), .D(g28219) );
  DFF_X1 DFF_406( .CK(CK), .Q(g577), .D(g28220) );
  DFF_X1 DFF_407( .CK(CK), .Q(g575), .D(g28221) );
  DFF_X1 DFF_408( .CK(CK), .Q(g579), .D(g28222) );
  DFF_X1 DFF_409( .CK(CK), .Q(g580), .D(g28223) );
  DFF_X1 DFF_410( .CK(CK), .Q(g578), .D(g28224) );
  DFF_X1 DFF_411( .CK(CK), .Q(g582), .D(g28225) );
  DFF_X1 DFF_412( .CK(CK), .Q(g583), .D(g28226) );
  DFF_X1 DFF_413( .CK(CK), .Q(g581), .D(g28227) );
  DFF_X1 DFF_414( .CK(CK), .Q(g585), .D(g28228) );
  DFF_X1 DFF_415( .CK(CK), .Q(g586), .D(g28229) );
  DFF_X1 DFF_416( .CK(CK), .Q(g584), .D(g28230) );
  DFF_X1 DFF_417( .CK(CK), .Q(g587), .D(g25985) );
  DFF_X1 DFF_418( .CK(CK), .Q(g590), .D(g25986) );
  DFF_X1 DFF_419( .CK(CK), .Q(g593), .D(g25987) );
  DFF_X1 DFF_420( .CK(CK), .Q(g596), .D(g25988) );
  DFF_X1 DFF_421( .CK(CK), .Q(g599), .D(g25989) );
  DFF_X1 DFF_422( .CK(CK), .Q(g602), .D(g25990) );
  DFF_X1 DFF_423( .CK(CK), .Q(g614), .D(g29135) );
  DFF_X2 DFF_424( .CK(CK), .Q(g617), .D(g29136) );
  DFF_X2 DFF_425( .CK(CK), .Q(g620), .D(g29137) );
  DFF_X2 DFF_426( .CK(CK), .Q(g605), .D(g29132) );
  DFF_X2 DFF_427( .CK(CK), .Q(g608), .D(g29133) );
  DFF_X2 DFF_428( .CK(CK), .Q(g611), .D(g29134) );
  DFF_X2 DFF_429( .CK(CK), .Q(g490), .D(g27194) );
  DFF_X2 DFF_430( .CK(CK), .Q(g493), .D(g27195) );
  DFF_X1 DFF_431( .CK(CK), .Q(g496), .D(g27196) );
  DFF_X1 DFF_432( .CK(CK), .Q(g506), .D(g8284) );
  DFF_X1 DFF_433( .CK(CK), .Q(g507), .D(g24295) );
  DFF_X1 DFF_434( .CK(CK), .Q(g508), .D(g19017) );
  DFF_X1 DFF_435( .CK(CK), .Q(g509), .D(g19018) );
  DFF_X1 DFF_436( .CK(CK), .Q(g514), .D(g19019) );
  DFF_X1 DFF_437( .CK(CK), .Q(g515), .D(g19020) );
  DFF_X1 DFF_438( .CK(CK), .Q(g516), .D(g23158) );
  DFF_X1 DFF_439( .CK(CK), .Q(g517), .D(g23157) );
  DFF_X1 DFF_440( .CK(CK), .Q(g518), .D(g23156) );
  DFF_X1 DFF_441( .CK(CK), .Q(g519), .D(g23155) );
  DFF_X1 DFF_442( .CK(CK), .Q(g520), .D(g23154) );
  DFF_X1 DFF_443( .CK(CK), .Q(g525), .D(g520) );
  DFF_X1 DFF_444( .CK(CK), .Q(g529), .D(g13410) );
  DFF_X1 DFF_445( .CK(CK), .Q(g530), .D(g13411) );
  DFF_X1 DFF_446( .CK(CK), .Q(g531), .D(g13412) );
  DFF_X1 DFF_447( .CK(CK), .Q(g532), .D(g13413) );
  DFF_X1 DFF_448( .CK(CK), .Q(g533), .D(g13414) );
  DFF_X1 DFF_449( .CK(CK), .Q(g534), .D(g13415) );
  DFF_X1 DFF_450( .CK(CK), .Q(g536), .D(g13416) );
  DFF_X1 DFF_451( .CK(CK), .Q(g537), .D(g13417) );
  DFF_X1 DFF_452( .CK(CK), .Q(g538), .D(g25984) );
  DFF_X1 DFF_453( .CK(CK), .Q(g541), .D(g13418) );
  DFF_X1 DFF_454( .CK(CK), .Q(g623), .D(g13420) );
  DFF_X1 DFF_455( .CK(CK), .Q(g626), .D(g623) );
  DFF_X1 DFF_456( .CK(CK), .Q(g629), .D(g626) );
  DFF_X1 DFF_457( .CK(CK), .Q(g630), .D(g20558) );
  DFF_X1 DFF_458( .CK(CK), .Q(g659), .D(g21943) );
  DFF_X1 DFF_459( .CK(CK), .Q(g640), .D(g23161) );
  DFF_X1 DFF_460( .CK(CK), .Q(g633), .D(g24296) );
  DFF_X1 DFF_461( .CK(CK), .Q(g653), .D(g25140) );
  DFF_X1 DFF_462( .CK(CK), .Q(g646), .D(g25991) );
  DFF_X1 DFF_463( .CK(CK), .Q(g660), .D(g26691) );
  DFF_X1 DFF_464( .CK(CK), .Q(g672), .D(g27197) );
  DFF_X1 DFF_465( .CK(CK), .Q(g666), .D(g27690) );
  DFF_X1 DFF_466( .CK(CK), .Q(g679), .D(g28231) );
  DFF_X1 DFF_467( .CK(CK), .Q(g686), .D(g28677) );
  DFF_X1 DFF_468( .CK(CK), .Q(g692), .D(g29138) );
  DFF_X1 DFF_469( .CK(CK), .Q(g699), .D(g23162) );
  DFF_X1 DFF_470( .CK(CK), .Q(g700), .D(g23163) );
  DFF_X1 DFF_471( .CK(CK), .Q(g698), .D(g23164) );
  DFF_X1 DFF_472( .CK(CK), .Q(g702), .D(g23165) );
  DFF_X1 DFF_473( .CK(CK), .Q(g703), .D(g23166) );
  DFF_X1 DFF_474( .CK(CK), .Q(g701), .D(g23167) );
  DFF_X1 DFF_475( .CK(CK), .Q(g705), .D(g23168) );
  DFF_X1 DFF_476( .CK(CK), .Q(g706), .D(g23169) );
  DFF_X1 DFF_477( .CK(CK), .Q(g704), .D(g23170) );
  DFF_X1 DFF_478( .CK(CK), .Q(g708), .D(g23171) );
  DFF_X1 DFF_479( .CK(CK), .Q(g709), .D(g23172) );
  DFF_X1 DFF_480( .CK(CK), .Q(g707), .D(g23173) );
  DFF_X1 DFF_481( .CK(CK), .Q(g711), .D(g23174) );
  DFF_X1 DFF_482( .CK(CK), .Q(g712), .D(g23175) );
  DFF_X1 DFF_483( .CK(CK), .Q(g710), .D(g23176) );
  DFF_X1 DFF_484( .CK(CK), .Q(g714), .D(g23177) );
  DFF_X1 DFF_485( .CK(CK), .Q(g715), .D(g23178) );
  DFF_X1 DFF_486( .CK(CK), .Q(g713), .D(g23179) );
  DFF_X2 DFF_487( .CK(CK), .Q(g717), .D(g23180) );
  DFF_X2 DFF_488( .CK(CK), .Q(g718), .D(g23181) );
  DFF_X2 DFF_489( .CK(CK), .Q(g716), .D(g23182) );
  DFF_X2 DFF_490( .CK(CK), .Q(g720), .D(g23183) );
  DFF_X2 DFF_491( .CK(CK), .Q(g721), .D(g23184) );
  DFF_X1 DFF_492( .CK(CK), .Q(g719), .D(g23185) );
  DFF_X1 DFF_493( .CK(CK), .Q(g723), .D(g23186) );
  DFF_X1 DFF_494( .CK(CK), .Q(g724), .D(g23187) );
  DFF_X1 DFF_495( .CK(CK), .Q(g722), .D(g23188) );
  DFF_X1 DFF_496( .CK(CK), .Q(g726), .D(g23189) );
  DFF_X1 DFF_497( .CK(CK), .Q(g727), .D(g23190) );
  DFF_X1 DFF_498( .CK(CK), .Q(g725), .D(g23191) );
  DFF_X1 DFF_499( .CK(CK), .Q(g729), .D(g23192) );
  DFF_X1 DFF_500( .CK(CK), .Q(g730), .D(g23193) );
  DFF_X1 DFF_501( .CK(CK), .Q(g728), .D(g23194) );
  DFF_X1 DFF_502( .CK(CK), .Q(g732), .D(g23195) );
  DFF_X1 DFF_503( .CK(CK), .Q(g733), .D(g23196) );
  DFF_X1 DFF_504( .CK(CK), .Q(g731), .D(g23197) );
  DFF_X1 DFF_505( .CK(CK), .Q(g735), .D(g26692) );
  DFF_X1 DFF_506( .CK(CK), .Q(g736), .D(g26693) );
  DFF_X1 DFF_507( .CK(CK), .Q(g734), .D(g26694) );
  DFF_X1 DFF_508( .CK(CK), .Q(g738), .D(g24297) );
  DFF_X1 DFF_509( .CK(CK), .Q(g739), .D(g24298) );
  DFF_X1 DFF_510( .CK(CK), .Q(g737), .D(g24299) );
  DFF_X1 DFF_511( .CK(CK), .Q(g826), .D(g13421) );
  DFF_X1 DFF_512( .CK(CK), .Q(g823), .D(g826) );
  DFF_X2 DFF_513( .CK(CK), .Q(g853), .D(g823) );
  DFF_X1 DFF_514( .CK(CK), .Q(g818), .D(g24300) );
  DFF_X1 DFF_515( .CK(CK), .Q(g819), .D(g24301) );
  DFF_X1 DFF_516( .CK(CK), .Q(g817), .D(g24302) );
  DFF_X1 DFF_517( .CK(CK), .Q(g821), .D(g24303) );
  DFF_X1 DFF_518( .CK(CK), .Q(g822), .D(g24304) );
  DFF_X1 DFF_519( .CK(CK), .Q(g820), .D(g24305) );
  DFF_X1 DFF_520( .CK(CK), .Q(g830), .D(g24306) );
  DFF_X1 DFF_521( .CK(CK), .Q(g831), .D(g24307) );
  DFF_X1 DFF_522( .CK(CK), .Q(g829), .D(g24308) );
  DFF_X1 DFF_523( .CK(CK), .Q(g833), .D(g24309) );
  DFF_X1 DFF_524( .CK(CK), .Q(g834), .D(g24310) );
  DFF_X1 DFF_525( .CK(CK), .Q(g832), .D(g24311) );
  DFF_X1 DFF_526( .CK(CK), .Q(g836), .D(g24312) );
  DFF_X1 DFF_527( .CK(CK), .Q(g837), .D(g24313) );
  DFF_X1 DFF_528( .CK(CK), .Q(g835), .D(g24314) );
  DFF_X1 DFF_529( .CK(CK), .Q(g839), .D(g24315) );
  DFF_X1 DFF_530( .CK(CK), .Q(g840), .D(g24316) );
  DFF_X1 DFF_531( .CK(CK), .Q(g838), .D(g24317) );
  DFF_X1 DFF_532( .CK(CK), .Q(g842), .D(g24318) );
  DFF_X1 DFF_533( .CK(CK), .Q(g843), .D(g24319) );
  DFF_X1 DFF_534( .CK(CK), .Q(g841), .D(g24320) );
  DFF_X1 DFF_535( .CK(CK), .Q(g845), .D(g24321) );
  DFF_X1 DFF_536( .CK(CK), .Q(g846), .D(g24322) );
  DFF_X1 DFF_537( .CK(CK), .Q(g844), .D(g24323) );
  DFF_X2 DFF_538( .CK(CK), .Q(g848), .D(g24324) );
  DFF_X2 DFF_539( .CK(CK), .Q(g849), .D(g24325) );
  DFF_X1 DFF_540( .CK(CK), .Q(g847), .D(g24326) );
  DFF_X1 DFF_541( .CK(CK), .Q(g851), .D(g24327) );
  DFF_X1 DFF_542( .CK(CK), .Q(g852), .D(g24328) );
  DFF_X1 DFF_543( .CK(CK), .Q(g850), .D(g24329) );
  DFF_X1 DFF_544( .CK(CK), .Q(g857), .D(g26696) );
  DFF_X1 DFF_545( .CK(CK), .Q(g858), .D(g26697) );
  DFF_X1 DFF_546( .CK(CK), .Q(g856), .D(g26698) );
  DFF_X1 DFF_547( .CK(CK), .Q(g860), .D(g26699) );
  DFF_X1 DFF_548( .CK(CK), .Q(g861), .D(g26700) );
  DFF_X1 DFF_549( .CK(CK), .Q(g859), .D(g26701) );
  DFF_X1 DFF_550( .CK(CK), .Q(g863), .D(g26702) );
  DFF_X1 DFF_551( .CK(CK), .Q(g864), .D(g26703) );
  DFF_X1 DFF_552( .CK(CK), .Q(g862), .D(g26704) );
  DFF_X1 DFF_553( .CK(CK), .Q(g866), .D(g26705) );
  DFF_X1 DFF_554( .CK(CK), .Q(g867), .D(g26706) );
  DFF_X1 DFF_555( .CK(CK), .Q(g865), .D(g26707) );
  DFF_X1 DFF_556( .CK(CK), .Q(g873), .D(g30521) );
  DFF_X1 DFF_557( .CK(CK), .Q(g876), .D(g30522) );
  DFF_X1 DFF_558( .CK(CK), .Q(g879), .D(g30523) );
  DFF_X1 DFF_559( .CK(CK), .Q(g918), .D(g30860) );
  DFF_X1 DFF_560( .CK(CK), .Q(g921), .D(g30861) );
  DFF_X1 DFF_561( .CK(CK), .Q(g924), .D(g30862) );
  DFF_X1 DFF_562( .CK(CK), .Q(g882), .D(g30854) );
  DFF_X1 DFF_563( .CK(CK), .Q(g885), .D(g30855) );
  DFF_X1 DFF_564( .CK(CK), .Q(g888), .D(g30856) );
  DFF_X1 DFF_565( .CK(CK), .Q(g927), .D(g30863) );
  DFF_X1 DFF_566( .CK(CK), .Q(g930), .D(g30864) );
  DFF_X1 DFF_567( .CK(CK), .Q(g933), .D(g30865) );
  DFF_X1 DFF_568( .CK(CK), .Q(g891), .D(g30524) );
  DFF_X1 DFF_569( .CK(CK), .Q(g894), .D(g30525) );
  DFF_X1 DFF_570( .CK(CK), .Q(g897), .D(g30526) );
  DFF_X1 DFF_571( .CK(CK), .Q(g936), .D(g30530) );
  DFF_X1 DFF_572( .CK(CK), .Q(g939), .D(g30531) );
  DFF_X1 DFF_573( .CK(CK), .Q(g942), .D(g30532) );
  DFF_X2 DFF_574( .CK(CK), .Q(g900), .D(g30527) );
  DFF_X1 DFF_575( .CK(CK), .Q(g903), .D(g30528) );
  DFF_X1 DFF_576( .CK(CK), .Q(g906), .D(g30529) );
  DFF_X1 DFF_577( .CK(CK), .Q(g945), .D(g30533) );
  DFF_X1 DFF_578( .CK(CK), .Q(g948), .D(g30534) );
  DFF_X1 DFF_579( .CK(CK), .Q(g951), .D(g30535) );
  DFF_X1 DFF_580( .CK(CK), .Q(g909), .D(g30857) );
  DFF_X1 DFF_581( .CK(CK), .Q(g912), .D(g30858) );
  DFF_X1 DFF_582( .CK(CK), .Q(g915), .D(g30859) );
  DFF_X1 DFF_583( .CK(CK), .Q(g954), .D(g30866) );
  DFF_X1 DFF_584( .CK(CK), .Q(g957), .D(g30867) );
  DFF_X1 DFF_585( .CK(CK), .Q(g960), .D(g30868) );
  DFF_X1 DFF_586( .CK(CK), .Q(g780), .D(g25992) );
  DFF_X1 DFF_587( .CK(CK), .Q(g776), .D(g26695) );
  DFF_X1 DFF_588( .CK(CK), .Q(g771), .D(g27198) );
  DFF_X1 DFF_589( .CK(CK), .Q(g767), .D(g27691) );
  DFF_X1 DFF_590( .CK(CK), .Q(g762), .D(g28232) );
  DFF_X1 DFF_591( .CK(CK), .Q(g758), .D(g28678) );
  DFF_X1 DFF_592( .CK(CK), .Q(g753), .D(g29139) );
  DFF_X1 DFF_593( .CK(CK), .Q(g749), .D(g29420) );
  DFF_X1 DFF_594( .CK(CK), .Q(g744), .D(g29634) );
  DFF_X1 DFF_595( .CK(CK), .Q(g740), .D(g29798) );
  DFF_X1 DFF_596( .CK(CK), .Q(g868), .D(g20559) );
  DFF_X1 DFF_597( .CK(CK), .Q(g870), .D(g868) );
  DFF_X1 DFF_598( .CK(CK), .Q(g869), .D(g870) );
  DFF_X1 DFF_599( .CK(CK), .Q(g963), .D(g13422) );
  DFF_X1 DFF_600( .CK(CK), .Q(g1092), .D(g963) );
  DFF_X1 DFF_601( .CK(CK), .Q(g1088), .D(g1092) );
  DFF_X1 DFF_602( .CK(CK), .Q(g996), .D(g11523) );
  DFF_X1 DFF_603( .CK(CK), .Q(g1041), .D(g28233) );
  DFF_X1 DFF_604( .CK(CK), .Q(g1030), .D(g28234) );
  DFF_X1 DFF_605( .CK(CK), .Q(g1033), .D(g28235) );
  DFF_X1 DFF_606( .CK(CK), .Q(g1056), .D(g28236) );
  DFF_X1 DFF_607( .CK(CK), .Q(g1045), .D(g28237) );
  DFF_X2 DFF_608( .CK(CK), .Q(g1048), .D(g28238) );
  DFF_X1 DFF_609( .CK(CK), .Q(g1071), .D(g28239) );
  DFF_X1 DFF_610( .CK(CK), .Q(g1060), .D(g28240) );
  DFF_X1 DFF_611( .CK(CK), .Q(g1063), .D(g28241) );
  DFF_X1 DFF_612( .CK(CK), .Q(g1085), .D(g28242) );
  DFF_X1 DFF_613( .CK(CK), .Q(g1075), .D(g28243) );
  DFF_X1 DFF_614( .CK(CK), .Q(g1078), .D(g28244) );
  DFF_X1 DFF_615( .CK(CK), .Q(g1095), .D(g29421) );
  DFF_X1 DFF_616( .CK(CK), .Q(g1098), .D(g29422) );
  DFF_X1 DFF_617( .CK(CK), .Q(g1101), .D(g29423) );
  DFF_X1 DFF_618( .CK(CK), .Q(g1104), .D(g29638) );
  DFF_X1 DFF_619( .CK(CK), .Q(g1107), .D(g29639) );
  DFF_X1 DFF_620( .CK(CK), .Q(g1110), .D(g29640) );
  DFF_X1 DFF_621( .CK(CK), .Q(g1114), .D(g29424) );
  DFF_X1 DFF_622( .CK(CK), .Q(g1115), .D(g29425) );
  DFF_X1 DFF_623( .CK(CK), .Q(g1113), .D(g29426) );
  DFF_X1 DFF_624( .CK(CK), .Q(g1116), .D(g27692) );
  DFF_X1 DFF_625( .CK(CK), .Q(g1119), .D(g27693) );
  DFF_X1 DFF_626( .CK(CK), .Q(g1122), .D(g27694) );
  DFF_X1 DFF_627( .CK(CK), .Q(g1125), .D(g27695) );
  DFF_X1 DFF_628( .CK(CK), .Q(g1128), .D(g27696) );
  DFF_X1 DFF_629( .CK(CK), .Q(g1131), .D(g27697) );
  DFF_X1 DFF_630( .CK(CK), .Q(g1135), .D(g28679) );
  DFF_X1 DFF_631( .CK(CK), .Q(g1136), .D(g28680) );
  DFF_X1 DFF_632( .CK(CK), .Q(g1134), .D(g28681) );
  DFF_X1 DFF_633( .CK(CK), .Q(g999), .D(g29799) );
  DFF_X1 DFF_634( .CK(CK), .Q(g1000), .D(g29800) );
  DFF_X1 DFF_635( .CK(CK), .Q(g1001), .D(g29801) );
  DFF_X1 DFF_636( .CK(CK), .Q(g1002), .D(g30869) );
  DFF_X1 DFF_637( .CK(CK), .Q(g1003), .D(g30870) );
  DFF_X1 DFF_638( .CK(CK), .Q(g1004), .D(g30871) );
  DFF_X1 DFF_639( .CK(CK), .Q(g1005), .D(g30713) );
  DFF_X1 DFF_640( .CK(CK), .Q(g1006), .D(g30714) );
  DFF_X1 DFF_641( .CK(CK), .Q(g1007), .D(g30715) );
  DFF_X1 DFF_642( .CK(CK), .Q(g1009), .D(g29635) );
  DFF_X1 DFF_643( .CK(CK), .Q(g1010), .D(g29636) );
  DFF_X1 DFF_644( .CK(CK), .Q(g1008), .D(g29637) );
  DFF_X1 DFF_645( .CK(CK), .Q(g1090), .D(g27206) );
  DFF_X1 DFF_646( .CK(CK), .Q(g1091), .D(g27207) );
  DFF_X1 DFF_647( .CK(CK), .Q(g1089), .D(g27208) );
  DFF_X1 DFF_648( .CK(CK), .Q(g1137), .D(g11536) );
  DFF_X1 DFF_649( .CK(CK), .Q(g1138), .D(g1137) );
  DFF_X1 DFF_650( .CK(CK), .Q(g1139), .D(g11537) );
  DFF_X1 DFF_651( .CK(CK), .Q(g1140), .D(g1139) );
  DFF_X1 DFF_652( .CK(CK), .Q(g1141), .D(g11538) );
  DFF_X1 DFF_653( .CK(CK), .Q(g966), .D(g1141) );
  DFF_X1 DFF_654( .CK(CK), .Q(g967), .D(g11518) );
  DFF_X1 DFF_655( .CK(CK), .Q(g968), .D(g967) );
  DFF_X1 DFF_656( .CK(CK), .Q(g969), .D(g11519) );
  DFF_X1 DFF_657( .CK(CK), .Q(g970), .D(g969) );
  DFF_X1 DFF_658( .CK(CK), .Q(g971), .D(g11520) );
  DFF_X1 DFF_659( .CK(CK), .Q(g972), .D(g971) );
  DFF_X1 DFF_660( .CK(CK), .Q(g973), .D(g11521) );
  DFF_X1 DFF_661( .CK(CK), .Q(g974), .D(g973) );
  DFF_X1 DFF_662( .CK(CK), .Q(g975), .D(g11522) );
  DFF_X1 DFF_663( .CK(CK), .Q(g976), .D(g975) );
  DFF_X1 DFF_664( .CK(CK), .Q(g977), .D(g13423) );
  DFF_X1 DFF_665( .CK(CK), .Q(g978), .D(g977) );
  DFF_X1 DFF_666( .CK(CK), .Q(g986), .D(g19024) );
  DFF_X1 DFF_667( .CK(CK), .Q(g992), .D(g27200) );
  DFF_X1 DFF_668( .CK(CK), .Q(g995), .D(g27201) );
  DFF_X1 DFF_669( .CK(CK), .Q(g984), .D(g27202) );
  DFF_X1 DFF_670( .CK(CK), .Q(g983), .D(g27203) );
  DFF_X1 DFF_671( .CK(CK), .Q(g982), .D(g27204) );
  DFF_X1 DFF_672( .CK(CK), .Q(g981), .D(g27205) );
  DFF_X1 DFF_673( .CK(CK), .Q(g991), .D(g19028) );
  DFF_X1 DFF_674( .CK(CK), .Q(g990), .D(g19027) );
  DFF_X1 DFF_675( .CK(CK), .Q(g989), .D(g19026) );
  DFF_X1 DFF_676( .CK(CK), .Q(g988), .D(g19025) );
  DFF_X1 DFF_677( .CK(CK), .Q(g987), .D(g25141) );
  DFF_X1 DFF_678( .CK(CK), .Q(g985), .D(g27199) );
  DFF_X1 DFF_679( .CK(CK), .Q(g1029), .D(g11524) );
  DFF_X1 DFF_680( .CK(CK), .Q(g1036), .D(g1029) );
  DFF_X2 DFF_681( .CK(CK), .Q(g1037), .D(g11525) );
  DFF_X1 DFF_682( .CK(CK), .Q(g1038), .D(g1037) );
  DFF_X1 DFF_683( .CK(CK), .Q(g1039), .D(g11526) );
  DFF_X1 DFF_684( .CK(CK), .Q(g1040), .D(g1039) );
  DFF_X1 DFF_685( .CK(CK), .Q(g1044), .D(g11527) );
  DFF_X1 DFF_686( .CK(CK), .Q(g1051), .D(g1044) );
  DFF_X1 DFF_687( .CK(CK), .Q(g1052), .D(g11528) );
  DFF_X1 DFF_688( .CK(CK), .Q(g1053), .D(g1052) );
  DFF_X1 DFF_689( .CK(CK), .Q(g1054), .D(g11529) );
  DFF_X1 DFF_690( .CK(CK), .Q(g1055), .D(g1054) );
  DFF_X1 DFF_691( .CK(CK), .Q(g1059), .D(g11530) );
  DFF_X1 DFF_692( .CK(CK), .Q(g1066), .D(g1059) );
  DFF_X1 DFF_693( .CK(CK), .Q(g1067), .D(g11531) );
  DFF_X1 DFF_694( .CK(CK), .Q(g1068), .D(g1067) );
  DFF_X1 DFF_695( .CK(CK), .Q(g1069), .D(g11532) );
  DFF_X1 DFF_696( .CK(CK), .Q(g1070), .D(g1069) );
  DFF_X1 DFF_697( .CK(CK), .Q(g1074), .D(g11533) );
  DFF_X1 DFF_698( .CK(CK), .Q(g1081), .D(g1074) );
  DFF_X1 DFF_699( .CK(CK), .Q(g1082), .D(g11534) );
  DFF_X1 DFF_700( .CK(CK), .Q(g1083), .D(g1082) );
  DFF_X1 DFF_701( .CK(CK), .Q(g1084), .D(g11535) );
  DFF_X1 DFF_702( .CK(CK), .Q(g1011), .D(g1084) );
  DFF_X1 DFF_703( .CK(CK), .Q(g1012), .D(g13424) );
  DFF_X1 DFF_704( .CK(CK), .Q(g1018), .D(g1012) );
  DFF_X1 DFF_705( .CK(CK), .Q(g1024), .D(g1018) );
  DFF_X1 DFF_706( .CK(CK), .Q(g1231), .D(g13435) );
  DFF_X1 DFF_707( .CK(CK), .Q(g1237), .D(g1231) );
  DFF_X1 DFF_708( .CK(CK), .Q(g1236), .D(g1237) );
  DFF_X1 DFF_709( .CK(CK), .Q(g1240), .D(g23198) );
  DFF_X1 DFF_710( .CK(CK), .Q(g1243), .D(g20560) );
  DFF_X1 DFF_711( .CK(CK), .Q(g1196), .D(g20561) );
  DFF_X1 DFF_712( .CK(CK), .Q(g1199), .D(g16469) );
  DFF_X1 DFF_713( .CK(CK), .Q(g1209), .D(g1199) );
  DFF_X1 DFF_714( .CK(CK), .Q(g1210), .D(g1209) );
  DFF_X1 DFF_715( .CK(CK), .Q(g1250), .D(g11539) );
  DFF_X1 DFF_716( .CK(CK), .Q(g1255), .D(g1250) );
  DFF_X1 DFF_717( .CK(CK), .Q(g1256), .D(g11542) );
  DFF_X1 DFF_718( .CK(CK), .Q(g1257), .D(g1256) );
  DFF_X1 DFF_719( .CK(CK), .Q(g1258), .D(g11543) );
  DFF_X1 DFF_720( .CK(CK), .Q(g1259), .D(g1258) );
  DFF_X1 DFF_721( .CK(CK), .Q(g1260), .D(g11544) );
  DFF_X1 DFF_722( .CK(CK), .Q(g1251), .D(g1260) );
  DFF_X1 DFF_723( .CK(CK), .Q(g1252), .D(g11540) );
  DFF_X1 DFF_724( .CK(CK), .Q(g1253), .D(g1252) );
  DFF_X1 DFF_725( .CK(CK), .Q(g1254), .D(g11541) );
  DFF_X1 DFF_726( .CK(CK), .Q(g1176), .D(g1254) );
  DFF_X1 DFF_727( .CK(CK), .Q(g1161), .D(g13425) );
  DFF_X1 DFF_728( .CK(CK), .Q(g1168), .D(g1161) );
  DFF_X2 DFF_729( .CK(CK), .Q(g1172), .D(g1168) );
  DFF_X1 DFF_730( .CK(CK), .Q(g1173), .D(g24333) );
  DFF_X1 DFF_731( .CK(CK), .Q(g1174), .D(g24334) );
  DFF_X1 DFF_732( .CK(CK), .Q(g1175), .D(g24335) );
  DFF_X1 DFF_733( .CK(CK), .Q(g1142), .D(g25150) );
  DFF_X1 DFF_734( .CK(CK), .Q(g1145), .D(g25142) );
  DFF_X1 DFF_735( .CK(CK), .Q(g1148), .D(g25143) );
  DFF_X1 DFF_736( .CK(CK), .Q(g1164), .D(g25147) );
  DFF_X1 DFF_737( .CK(CK), .Q(g1165), .D(g25148) );
  DFF_X1 DFF_738( .CK(CK), .Q(g1166), .D(g25149) );
  DFF_X1 DFF_739( .CK(CK), .Q(g1167), .D(g24330) );
  DFF_X1 DFF_740( .CK(CK), .Q(g1171), .D(g24331) );
  DFF_X1 DFF_741( .CK(CK), .Q(g1151), .D(g24332) );
  DFF_X1 DFF_742( .CK(CK), .Q(g1152), .D(g25144) );
  DFF_X1 DFF_743( .CK(CK), .Q(g1155), .D(g25145) );
  DFF_X1 DFF_744( .CK(CK), .Q(g1158), .D(g25146) );
  DFF_X1 DFF_745( .CK(CK), .Q(g1214), .D(g16470) );
  DFF_X1 DFF_746( .CK(CK), .Q(g1221), .D(g1214) );
  DFF_X1 DFF_747( .CK(CK), .Q(g1228), .D(g1221) );
  DFF_X1 DFF_748( .CK(CK), .Q(g1229), .D(g19033) );
  DFF_X1 DFF_749( .CK(CK), .Q(g1230), .D(g1229) );
  DFF_X1 DFF_750( .CK(CK), .Q(g1234), .D(g27217) );
  DFF_X1 DFF_751( .CK(CK), .Q(g1235), .D(g19034) );
  DFF_X1 DFF_752( .CK(CK), .Q(g1186), .D(g1235) );
  DFF_X1 DFF_753( .CK(CK), .Q(g1244), .D(g19035) );
  DFF_X1 DFF_754( .CK(CK), .Q(g1245), .D(g1244) );
  DFF_X1 DFF_755( .CK(CK), .Q(g1262), .D(g28245) );
  DFF_X1 DFF_756( .CK(CK), .Q(g1263), .D(g28246) );
  DFF_X1 DFF_757( .CK(CK), .Q(g1261), .D(g28247) );
  DFF_X1 DFF_758( .CK(CK), .Q(g1265), .D(g28248) );
  DFF_X1 DFF_759( .CK(CK), .Q(g1266), .D(g28249) );
  DFF_X1 DFF_760( .CK(CK), .Q(g1264), .D(g28250) );
  DFF_X1 DFF_761( .CK(CK), .Q(g1268), .D(g28251) );
  DFF_X1 DFF_762( .CK(CK), .Q(g1269), .D(g28252) );
  DFF_X1 DFF_763( .CK(CK), .Q(g1267), .D(g28253) );
  DFF_X1 DFF_764( .CK(CK), .Q(g1271), .D(g28254) );
  DFF_X1 DFF_765( .CK(CK), .Q(g1272), .D(g28255) );
  DFF_X1 DFF_766( .CK(CK), .Q(g1270), .D(g28256) );
  DFF_X1 DFF_767( .CK(CK), .Q(g1273), .D(g25994) );
  DFF_X1 DFF_768( .CK(CK), .Q(g1276), .D(g25995) );
  DFF_X1 DFF_769( .CK(CK), .Q(g1279), .D(g25996) );
  DFF_X1 DFF_770( .CK(CK), .Q(g1282), .D(g25997) );
  DFF_X1 DFF_771( .CK(CK), .Q(g1285), .D(g25998) );
  DFF_X1 DFF_772( .CK(CK), .Q(g1288), .D(g25999) );
  DFF_X1 DFF_773( .CK(CK), .Q(g1300), .D(g29143) );
  DFF_X1 DFF_774( .CK(CK), .Q(g1303), .D(g29144) );
  DFF_X1 DFF_775( .CK(CK), .Q(g1306), .D(g29145) );
  DFF_X1 DFF_776( .CK(CK), .Q(g1291), .D(g29140) );
  DFF_X1 DFF_777( .CK(CK), .Q(g1294), .D(g29141) );
  DFF_X1 DFF_778( .CK(CK), .Q(g1297), .D(g29142) );
  DFF_X1 DFF_779( .CK(CK), .Q(g1177), .D(g27209) );
  DFF_X1 DFF_780( .CK(CK), .Q(g1180), .D(g27210) );
  DFF_X1 DFF_781( .CK(CK), .Q(g1183), .D(g27211) );
  DFF_X1 DFF_782( .CK(CK), .Q(g1192), .D(g8293) );
  DFF_X1 DFF_783( .CK(CK), .Q(g1193), .D(g24336) );
  DFF_X1 DFF_784( .CK(CK), .Q(g1194), .D(g19029) );
  DFF_X1 DFF_785( .CK(CK), .Q(g1195), .D(g19030) );
  DFF_X1 DFF_786( .CK(CK), .Q(g1200), .D(g19031) );
  DFF_X1 DFF_787( .CK(CK), .Q(g1201), .D(g19032) );
  DFF_X1 DFF_788( .CK(CK), .Q(g1202), .D(g27216) );
  DFF_X1 DFF_789( .CK(CK), .Q(g1203), .D(g27215) );
  DFF_X1 DFF_790( .CK(CK), .Q(g1204), .D(g27214) );
  DFF_X1 DFF_791( .CK(CK), .Q(g1205), .D(g27213) );
  DFF_X1 DFF_792( .CK(CK), .Q(g1206), .D(g27212) );
  DFF_X1 DFF_793( .CK(CK), .Q(g1211), .D(g1206) );
  DFF_X1 DFF_794( .CK(CK), .Q(g1215), .D(g13426) );
  DFF_X1 DFF_795( .CK(CK), .Q(g1216), .D(g13427) );
  DFF_X1 DFF_796( .CK(CK), .Q(g1217), .D(g13428) );
  DFF_X1 DFF_797( .CK(CK), .Q(g1218), .D(g13429) );
  DFF_X1 DFF_798( .CK(CK), .Q(g1219), .D(g13430) );
  DFF_X2 DFF_799( .CK(CK), .Q(g1220), .D(g13431) );
  DFF_X1 DFF_800( .CK(CK), .Q(g1222), .D(g13432) );
  DFF_X1 DFF_801( .CK(CK), .Q(g1223), .D(g13433) );
  DFF_X1 DFF_802( .CK(CK), .Q(g1224), .D(g25993) );
  DFF_X1 DFF_803( .CK(CK), .Q(g1227), .D(g13434) );
  DFF_X1 DFF_804( .CK(CK), .Q(g1309), .D(g13436) );
  DFF_X1 DFF_805( .CK(CK), .Q(g1312), .D(g1309) );
  DFF_X1 DFF_806( .CK(CK), .Q(g1315), .D(g1312) );
  DFF_X1 DFF_807( .CK(CK), .Q(g1316), .D(g20562) );
  DFF_X1 DFF_808( .CK(CK), .Q(g1345), .D(g21944) );
  DFF_X1 DFF_809( .CK(CK), .Q(g1326), .D(g23199) );
  DFF_X1 DFF_810( .CK(CK), .Q(g1319), .D(g24337) );
  DFF_X1 DFF_811( .CK(CK), .Q(g1339), .D(g25151) );
  DFF_X1 DFF_812( .CK(CK), .Q(g1332), .D(g26000) );
  DFF_X1 DFF_813( .CK(CK), .Q(g1346), .D(g26708) );
  DFF_X1 DFF_814( .CK(CK), .Q(g1358), .D(g27218) );
  DFF_X1 DFF_815( .CK(CK), .Q(g1352), .D(g27698) );
  DFF_X1 DFF_816( .CK(CK), .Q(g1365), .D(g28257) );
  DFF_X1 DFF_817( .CK(CK), .Q(g1372), .D(g28682) );
  DFF_X1 DFF_818( .CK(CK), .Q(g1378), .D(g29146) );
  DFF_X1 DFF_819( .CK(CK), .Q(g1385), .D(g23200) );
  DFF_X1 DFF_820( .CK(CK), .Q(g1386), .D(g23201) );
  DFF_X1 DFF_821( .CK(CK), .Q(g1384), .D(g23202) );
  DFF_X1 DFF_822( .CK(CK), .Q(g1388), .D(g23203) );
  DFF_X1 DFF_823( .CK(CK), .Q(g1389), .D(g23204) );
  DFF_X1 DFF_824( .CK(CK), .Q(g1387), .D(g23205) );
  DFF_X1 DFF_825( .CK(CK), .Q(g1391), .D(g23206) );
  DFF_X1 DFF_826( .CK(CK), .Q(g1392), .D(g23207) );
  DFF_X1 DFF_827( .CK(CK), .Q(g1390), .D(g23208) );
  DFF_X1 DFF_828( .CK(CK), .Q(g1394), .D(g23209) );
  DFF_X1 DFF_829( .CK(CK), .Q(g1395), .D(g23210) );
  DFF_X1 DFF_830( .CK(CK), .Q(g1393), .D(g23211) );
  DFF_X1 DFF_831( .CK(CK), .Q(g1397), .D(g23212) );
  DFF_X1 DFF_832( .CK(CK), .Q(g1398), .D(g23213) );
  DFF_X2 DFF_833( .CK(CK), .Q(g1396), .D(g23214) );
  DFF_X1 DFF_834( .CK(CK), .Q(g1400), .D(g23215) );
  DFF_X1 DFF_835( .CK(CK), .Q(g1401), .D(g23216) );
  DFF_X1 DFF_836( .CK(CK), .Q(g1399), .D(g23217) );
  DFF_X1 DFF_837( .CK(CK), .Q(g1403), .D(g23218) );
  DFF_X1 DFF_838( .CK(CK), .Q(g1404), .D(g23219) );
  DFF_X1 DFF_839( .CK(CK), .Q(g1402), .D(g23220) );
  DFF_X1 DFF_840( .CK(CK), .Q(g1406), .D(g23221) );
  DFF_X1 DFF_841( .CK(CK), .Q(g1407), .D(g23222) );
  DFF_X1 DFF_842( .CK(CK), .Q(g1405), .D(g23223) );
  DFF_X1 DFF_843( .CK(CK), .Q(g1409), .D(g23224) );
  DFF_X1 DFF_844( .CK(CK), .Q(g1410), .D(g23225) );
  DFF_X1 DFF_845( .CK(CK), .Q(g1408), .D(g23226) );
  DFF_X1 DFF_846( .CK(CK), .Q(g1412), .D(g23227) );
  DFF_X1 DFF_847( .CK(CK), .Q(g1413), .D(g23228) );
  DFF_X1 DFF_848( .CK(CK), .Q(g1411), .D(g23229) );
  DFF_X1 DFF_849( .CK(CK), .Q(g1415), .D(g23230) );
  DFF_X1 DFF_850( .CK(CK), .Q(g1416), .D(g23231) );
  DFF_X1 DFF_851( .CK(CK), .Q(g1414), .D(g23232) );
  DFF_X1 DFF_852( .CK(CK), .Q(g1418), .D(g23233) );
  DFF_X1 DFF_853( .CK(CK), .Q(g1419), .D(g23234) );
  DFF_X1 DFF_854( .CK(CK), .Q(g1417), .D(g23235) );
  DFF_X1 DFF_855( .CK(CK), .Q(g1421), .D(g26709) );
  DFF_X1 DFF_856( .CK(CK), .Q(g1422), .D(g26710) );
  DFF_X1 DFF_857( .CK(CK), .Q(g1420), .D(g26711) );
  DFF_X1 DFF_858( .CK(CK), .Q(g1424), .D(g24338) );
  DFF_X1 DFF_859( .CK(CK), .Q(g1425), .D(g24339) );
  DFF_X1 DFF_860( .CK(CK), .Q(g1423), .D(g24340) );
  DFF_X1 DFF_861( .CK(CK), .Q(g1520), .D(g13437) );
  DFF_X1 DFF_862( .CK(CK), .Q(g1517), .D(g1520) );
  DFF_X1 DFF_863( .CK(CK), .Q(g1547), .D(g1517) );
  DFF_X1 DFF_864( .CK(CK), .Q(g1512), .D(g24341) );
  DFF_X1 DFF_865( .CK(CK), .Q(g1513), .D(g24342) );
  DFF_X1 DFF_866( .CK(CK), .Q(g1511), .D(g24343) );
  DFF_X1 DFF_867( .CK(CK), .Q(g1515), .D(g24344) );
  DFF_X1 DFF_868( .CK(CK), .Q(g1516), .D(g24345) );
  DFF_X1 DFF_869( .CK(CK), .Q(g1514), .D(g24346) );
  DFF_X1 DFF_870( .CK(CK), .Q(g1524), .D(g24347) );
  DFF_X1 DFF_871( .CK(CK), .Q(g1525), .D(g24348) );
  DFF_X1 DFF_872( .CK(CK), .Q(g1523), .D(g24349) );
  DFF_X1 DFF_873( .CK(CK), .Q(g1527), .D(g24350) );
  DFF_X1 DFF_874( .CK(CK), .Q(g1528), .D(g24351) );
  DFF_X1 DFF_875( .CK(CK), .Q(g1526), .D(g24352) );
  DFF_X1 DFF_876( .CK(CK), .Q(g1530), .D(g24353) );
  DFF_X1 DFF_877( .CK(CK), .Q(g1531), .D(g24354) );
  DFF_X1 DFF_878( .CK(CK), .Q(g1529), .D(g24355) );
  DFF_X1 DFF_879( .CK(CK), .Q(g1533), .D(g24356) );
  DFF_X1 DFF_880( .CK(CK), .Q(g1534), .D(g24357) );
  DFF_X1 DFF_881( .CK(CK), .Q(g1532), .D(g24358) );
  DFF_X1 DFF_882( .CK(CK), .Q(g1536), .D(g24359) );
  DFF_X1 DFF_883( .CK(CK), .Q(g1537), .D(g24360) );
  DFF_X1 DFF_884( .CK(CK), .Q(g1535), .D(g24361) );
  DFF_X1 DFF_885( .CK(CK), .Q(g1539), .D(g24362) );
  DFF_X1 DFF_886( .CK(CK), .Q(g1540), .D(g24363) );
  DFF_X1 DFF_887( .CK(CK), .Q(g1538), .D(g24364) );
  DFF_X1 DFF_888( .CK(CK), .Q(g1542), .D(g24365) );
  DFF_X1 DFF_889( .CK(CK), .Q(g1543), .D(g24366) );
  DFF_X1 DFF_890( .CK(CK), .Q(g1541), .D(g24367) );
  DFF_X1 DFF_891( .CK(CK), .Q(g1545), .D(g24368) );
  DFF_X1 DFF_892( .CK(CK), .Q(g1546), .D(g24369) );
  DFF_X1 DFF_893( .CK(CK), .Q(g1544), .D(g24370) );
  DFF_X1 DFF_894( .CK(CK), .Q(g1551), .D(g26713) );
  DFF_X1 DFF_895( .CK(CK), .Q(g1552), .D(g26714) );
  DFF_X1 DFF_896( .CK(CK), .Q(g1550), .D(g26715) );
  DFF_X1 DFF_897( .CK(CK), .Q(g1554), .D(g26716) );
  DFF_X1 DFF_898( .CK(CK), .Q(g1555), .D(g26717) );
  DFF_X1 DFF_899( .CK(CK), .Q(g1553), .D(g26718) );
  DFF_X1 DFF_900( .CK(CK), .Q(g1557), .D(g26719) );
  DFF_X1 DFF_901( .CK(CK), .Q(g1558), .D(g26720) );
  DFF_X1 DFF_902( .CK(CK), .Q(g1556), .D(g26721) );
  DFF_X1 DFF_903( .CK(CK), .Q(g1560), .D(g26722) );
  DFF_X1 DFF_904( .CK(CK), .Q(g1561), .D(g26723) );
  DFF_X1 DFF_905( .CK(CK), .Q(g1559), .D(g26724) );
  DFF_X1 DFF_906( .CK(CK), .Q(g1567), .D(g30536) );
  DFF_X1 DFF_907( .CK(CK), .Q(g1570), .D(g30537) );
  DFF_X2 DFF_908( .CK(CK), .Q(g1573), .D(g30538) );
  DFF_X1 DFF_909( .CK(CK), .Q(g1612), .D(g30878) );
  DFF_X1 DFF_910( .CK(CK), .Q(g1615), .D(g30879) );
  DFF_X1 DFF_911( .CK(CK), .Q(g1618), .D(g30880) );
  DFF_X1 DFF_912( .CK(CK), .Q(g1576), .D(g30872) );
  DFF_X1 DFF_913( .CK(CK), .Q(g1579), .D(g30873) );
  DFF_X1 DFF_914( .CK(CK), .Q(g1582), .D(g30874) );
  DFF_X1 DFF_915( .CK(CK), .Q(g1621), .D(g30881) );
  DFF_X1 DFF_916( .CK(CK), .Q(g1624), .D(g30882) );
  DFF_X1 DFF_917( .CK(CK), .Q(g1627), .D(g30883) );
  DFF_X1 DFF_918( .CK(CK), .Q(g1585), .D(g30539) );
  DFF_X1 DFF_919( .CK(CK), .Q(g1588), .D(g30540) );
  DFF_X1 DFF_920( .CK(CK), .Q(g1591), .D(g30541) );
  DFF_X1 DFF_921( .CK(CK), .Q(g1630), .D(g30545) );
  DFF_X1 DFF_922( .CK(CK), .Q(g1633), .D(g30546) );
  DFF_X1 DFF_923( .CK(CK), .Q(g1636), .D(g30547) );
  DFF_X1 DFF_924( .CK(CK), .Q(g1594), .D(g30542) );
  DFF_X1 DFF_925( .CK(CK), .Q(g1597), .D(g30543) );
  DFF_X1 DFF_926( .CK(CK), .Q(g1600), .D(g30544) );
  DFF_X1 DFF_927( .CK(CK), .Q(g1639), .D(g30548) );
  DFF_X1 DFF_928( .CK(CK), .Q(g1642), .D(g30549) );
  DFF_X1 DFF_929( .CK(CK), .Q(g1645), .D(g30550) );
  DFF_X1 DFF_930( .CK(CK), .Q(g1603), .D(g30875) );
  DFF_X1 DFF_931( .CK(CK), .Q(g1606), .D(g30876) );
  DFF_X1 DFF_932( .CK(CK), .Q(g1609), .D(g30877) );
  DFF_X1 DFF_933( .CK(CK), .Q(g1648), .D(g30884) );
  DFF_X1 DFF_934( .CK(CK), .Q(g1651), .D(g30885) );
  DFF_X1 DFF_935( .CK(CK), .Q(g1654), .D(g30886) );
  DFF_X1 DFF_936( .CK(CK), .Q(g1466), .D(g26001) );
  DFF_X1 DFF_937( .CK(CK), .Q(g1462), .D(g26712) );
  DFF_X1 DFF_938( .CK(CK), .Q(g1457), .D(g27219) );
  DFF_X1 DFF_939( .CK(CK), .Q(g1453), .D(g27699) );
  DFF_X1 DFF_940( .CK(CK), .Q(g1448), .D(g28258) );
  DFF_X1 DFF_941( .CK(CK), .Q(g1444), .D(g28683) );
  DFF_X1 DFF_942( .CK(CK), .Q(g1439), .D(g29147) );
  DFF_X1 DFF_943( .CK(CK), .Q(g1435), .D(g29427) );
  DFF_X1 DFF_944( .CK(CK), .Q(g1430), .D(g29641) );
  DFF_X1 DFF_945( .CK(CK), .Q(g1426), .D(g29802) );
  DFF_X1 DFF_946( .CK(CK), .Q(g1562), .D(g20563) );
  DFF_X1 DFF_947( .CK(CK), .Q(g1564), .D(g1562) );
  DFF_X1 DFF_948( .CK(CK), .Q(g1563), .D(g1564) );
  DFF_X1 DFF_949( .CK(CK), .Q(g1657), .D(g13438) );
  DFF_X1 DFF_950( .CK(CK), .Q(g1786), .D(g1657) );
  DFF_X1 DFF_951( .CK(CK), .Q(g1782), .D(g1786) );
  DFF_X1 DFF_952( .CK(CK), .Q(g1690), .D(g11550) );
  DFF_X2 DFF_953( .CK(CK), .Q(g1735), .D(g28259) );
  DFF_X1 DFF_954( .CK(CK), .Q(g1724), .D(g28260) );
  DFF_X1 DFF_955( .CK(CK), .Q(g1727), .D(g28261) );
  DFF_X1 DFF_956( .CK(CK), .Q(g1750), .D(g28262) );
  DFF_X1 DFF_957( .CK(CK), .Q(g1739), .D(g28263) );
  DFF_X1 DFF_958( .CK(CK), .Q(g1742), .D(g28264) );
  DFF_X1 DFF_959( .CK(CK), .Q(g1765), .D(g28265) );
  DFF_X1 DFF_960( .CK(CK), .Q(g1754), .D(g28266) );
  DFF_X1 DFF_961( .CK(CK), .Q(g1757), .D(g28267) );
  DFF_X1 DFF_962( .CK(CK), .Q(g1779), .D(g28268) );
  DFF_X1 DFF_963( .CK(CK), .Q(g1769), .D(g28269) );
  DFF_X1 DFF_964( .CK(CK), .Q(g1772), .D(g28270) );
  DFF_X1 DFF_965( .CK(CK), .Q(g1789), .D(g29434) );
  DFF_X1 DFF_966( .CK(CK), .Q(g1792), .D(g29435) );
  DFF_X1 DFF_967( .CK(CK), .Q(g1795), .D(g29436) );
  DFF_X1 DFF_968( .CK(CK), .Q(g1798), .D(g29645) );
  DFF_X1 DFF_969( .CK(CK), .Q(g1801), .D(g29646) );
  DFF_X1 DFF_970( .CK(CK), .Q(g1804), .D(g29647) );
  DFF_X1 DFF_971( .CK(CK), .Q(g1808), .D(g29437) );
  DFF_X1 DFF_972( .CK(CK), .Q(g1809), .D(g29438) );
  DFF_X1 DFF_973( .CK(CK), .Q(g1807), .D(g29439) );
  DFF_X1 DFF_974( .CK(CK), .Q(g1810), .D(g27700) );
  DFF_X1 DFF_975( .CK(CK), .Q(g1813), .D(g27701) );
  DFF_X2 DFF_976( .CK(CK), .Q(g1816), .D(g27702) );
  DFF_X2 DFF_977( .CK(CK), .Q(g1819), .D(g27703) );
  DFF_X1 DFF_978( .CK(CK), .Q(g1822), .D(g27704) );
  DFF_X1 DFF_979( .CK(CK), .Q(g1825), .D(g27705) );
  DFF_X1 DFF_980( .CK(CK), .Q(g1829), .D(g28684) );
  DFF_X1 DFF_981( .CK(CK), .Q(g1830), .D(g28685) );
  DFF_X1 DFF_982( .CK(CK), .Q(g1828), .D(g28686) );
  DFF_X1 DFF_983( .CK(CK), .Q(g1693), .D(g29803) );
  DFF_X1 DFF_984( .CK(CK), .Q(g1694), .D(g29804) );
  DFF_X1 DFF_985( .CK(CK), .Q(g1695), .D(g29805) );
  DFF_X1 DFF_986( .CK(CK), .Q(g1696), .D(g30887) );
  DFF_X1 DFF_987( .CK(CK), .Q(g1697), .D(g30888) );
  DFF_X1 DFF_988( .CK(CK), .Q(g1698), .D(g30889) );
  DFF_X1 DFF_989( .CK(CK), .Q(g1699), .D(g30716) );
  DFF_X1 DFF_990( .CK(CK), .Q(g1700), .D(g30717) );
  DFF_X1 DFF_991( .CK(CK), .Q(g1701), .D(g30718) );
  DFF_X1 DFF_992( .CK(CK), .Q(g1703), .D(g29642) );
  DFF_X1 DFF_993( .CK(CK), .Q(g1704), .D(g29643) );
  DFF_X1 DFF_994( .CK(CK), .Q(g1702), .D(g29644) );
  DFF_X1 DFF_995( .CK(CK), .Q(g1784), .D(g27221) );
  DFF_X1 DFF_996( .CK(CK), .Q(g1785), .D(g27222) );
  DFF_X1 DFF_997( .CK(CK), .Q(g1783), .D(g27223) );
  DFF_X1 DFF_998( .CK(CK), .Q(g1831), .D(g11563) );
  DFF_X1 DFF_999( .CK(CK), .Q(g1832), .D(g1831) );
  DFF_X1 DFF_1000( .CK(CK), .Q(g1833), .D(g11564) );
  DFF_X1 DFF_1001( .CK(CK), .Q(g1834), .D(g1833) );
  DFF_X1 DFF_1002( .CK(CK), .Q(g1835), .D(g11565) );
  DFF_X1 DFF_1003( .CK(CK), .Q(g1660), .D(g1835) );
  DFF_X1 DFF_1004( .CK(CK), .Q(g1661), .D(g11545) );
  DFF_X1 DFF_1005( .CK(CK), .Q(g1662), .D(g1661) );
  DFF_X1 DFF_1006( .CK(CK), .Q(g1663), .D(g11546) );
  DFF_X1 DFF_1007( .CK(CK), .Q(g1664), .D(g1663) );
  DFF_X1 DFF_1008( .CK(CK), .Q(g1665), .D(g11547) );
  DFF_X1 DFF_1009( .CK(CK), .Q(g1666), .D(g1665) );
  DFF_X1 DFF_1010( .CK(CK), .Q(g1667), .D(g11548) );
  DFF_X2 DFF_1011( .CK(CK), .Q(g1668), .D(g1667) );
  DFF_X1 DFF_1012( .CK(CK), .Q(g1669), .D(g11549) );
  DFF_X1 DFF_1013( .CK(CK), .Q(g1670), .D(g1669) );
  DFF_X1 DFF_1014( .CK(CK), .Q(g1671), .D(g13439) );
  DFF_X1 DFF_1015( .CK(CK), .Q(g1672), .D(g1671) );
  DFF_X1 DFF_1016( .CK(CK), .Q(g1680), .D(g19036) );
  DFF_X1 DFF_1017( .CK(CK), .Q(g1686), .D(g29428) );
  DFF_X1 DFF_1018( .CK(CK), .Q(g1689), .D(g29429) );
  DFF_X1 DFF_1019( .CK(CK), .Q(g1678), .D(g29430) );
  DFF_X1 DFF_1020( .CK(CK), .Q(g1677), .D(g29431) );
  DFF_X1 DFF_1021( .CK(CK), .Q(g1676), .D(g29432) );
  DFF_X1 DFF_1022( .CK(CK), .Q(g1675), .D(g29433) );
  DFF_X1 DFF_1023( .CK(CK), .Q(g1685), .D(g19040) );
  DFF_X1 DFF_1024( .CK(CK), .Q(g1684), .D(g19039) );
  DFF_X1 DFF_1025( .CK(CK), .Q(g1683), .D(g19038) );
  DFF_X1 DFF_1026( .CK(CK), .Q(g1682), .D(g19037) );
  DFF_X1 DFF_1027( .CK(CK), .Q(g1681), .D(g25152) );
  DFF_X1 DFF_1028( .CK(CK), .Q(g1679), .D(g27220) );
  DFF_X1 DFF_1029( .CK(CK), .Q(g1723), .D(g11551) );
  DFF_X1 DFF_1030( .CK(CK), .Q(g1730), .D(g1723) );
  DFF_X2 DFF_1031( .CK(CK), .Q(g1731), .D(g11552) );
  DFF_X1 DFF_1032( .CK(CK), .Q(g1732), .D(g1731) );
  DFF_X1 DFF_1033( .CK(CK), .Q(g1733), .D(g11553) );
  DFF_X1 DFF_1034( .CK(CK), .Q(g1734), .D(g1733) );
  DFF_X1 DFF_1035( .CK(CK), .Q(g1738), .D(g11554) );
  DFF_X1 DFF_1036( .CK(CK), .Q(g1745), .D(g1738) );
  DFF_X1 DFF_1037( .CK(CK), .Q(g1746), .D(g11555) );
  DFF_X1 DFF_1038( .CK(CK), .Q(g1747), .D(g1746) );
  DFF_X1 DFF_1039( .CK(CK), .Q(g1748), .D(g11556) );
  DFF_X1 DFF_1040( .CK(CK), .Q(g1749), .D(g1748) );
  DFF_X1 DFF_1041( .CK(CK), .Q(g1753), .D(g11557) );
  DFF_X1 DFF_1042( .CK(CK), .Q(g1760), .D(g1753) );
  DFF_X1 DFF_1043( .CK(CK), .Q(g1761), .D(g11558) );
  DFF_X1 DFF_1044( .CK(CK), .Q(g1762), .D(g1761) );
  DFF_X1 DFF_1045( .CK(CK), .Q(g1763), .D(g11559) );
  DFF_X1 DFF_1046( .CK(CK), .Q(g1764), .D(g1763) );
  DFF_X1 DFF_1047( .CK(CK), .Q(g1768), .D(g11560) );
  DFF_X1 DFF_1048( .CK(CK), .Q(g1775), .D(g1768) );
  DFF_X1 DFF_1049( .CK(CK), .Q(g1776), .D(g11561) );
  DFF_X1 DFF_1050( .CK(CK), .Q(g1777), .D(g1776) );
  DFF_X1 DFF_1051( .CK(CK), .Q(g1778), .D(g11562) );
  DFF_X1 DFF_1052( .CK(CK), .Q(g1705), .D(g1778) );
  DFF_X1 DFF_1053( .CK(CK), .Q(g1706), .D(g13440) );
  DFF_X1 DFF_1054( .CK(CK), .Q(g1712), .D(g1706) );
  DFF_X1 DFF_1055( .CK(CK), .Q(g1718), .D(g1712) );
  DFF_X1 DFF_1056( .CK(CK), .Q(g1925), .D(g13451) );
  DFF_X1 DFF_1057( .CK(CK), .Q(g1931), .D(g1925) );
  DFF_X1 DFF_1058( .CK(CK), .Q(g1930), .D(g1931) );
  DFF_X1 DFF_1059( .CK(CK), .Q(g1934), .D(g23236) );
  DFF_X1 DFF_1060( .CK(CK), .Q(g1937), .D(g20564) );
  DFF_X1 DFF_1061( .CK(CK), .Q(g1890), .D(g20565) );
  DFF_X1 DFF_1062( .CK(CK), .Q(g1893), .D(g16471) );
  DFF_X1 DFF_1063( .CK(CK), .Q(g1903), .D(g1893) );
  DFF_X1 DFF_1064( .CK(CK), .Q(g1904), .D(g1903) );
  DFF_X1 DFF_1065( .CK(CK), .Q(g1944), .D(g11566) );
  DFF_X1 DFF_1066( .CK(CK), .Q(g1949), .D(g1944) );
  DFF_X1 DFF_1067( .CK(CK), .Q(g1950), .D(g11569) );
  DFF_X1 DFF_1068( .CK(CK), .Q(g1951), .D(g1950) );
  DFF_X1 DFF_1069( .CK(CK), .Q(g1952), .D(g11570) );
  DFF_X1 DFF_1070( .CK(CK), .Q(g1953), .D(g1952) );
  DFF_X1 DFF_1071( .CK(CK), .Q(g1954), .D(g11571) );
  DFF_X1 DFF_1072( .CK(CK), .Q(g1945), .D(g1954) );
  DFF_X1 DFF_1073( .CK(CK), .Q(g1946), .D(g11567) );
  DFF_X1 DFF_1074( .CK(CK), .Q(g1947), .D(g1946) );
  DFF_X2 DFF_1075( .CK(CK), .Q(g1948), .D(g11568) );
  DFF_X1 DFF_1076( .CK(CK), .Q(g1870), .D(g1948) );
  DFF_X1 DFF_1077( .CK(CK), .Q(g1855), .D(g13441) );
  DFF_X1 DFF_1078( .CK(CK), .Q(g1862), .D(g1855) );
  DFF_X1 DFF_1079( .CK(CK), .Q(g1866), .D(g1862) );
  DFF_X1 DFF_1080( .CK(CK), .Q(g1867), .D(g24374) );
  DFF_X1 DFF_1081( .CK(CK), .Q(g1868), .D(g24375) );
  DFF_X1 DFF_1082( .CK(CK), .Q(g1869), .D(g24376) );
  DFF_X1 DFF_1083( .CK(CK), .Q(g1836), .D(g25161) );
  DFF_X1 DFF_1084( .CK(CK), .Q(g1839), .D(g25153) );
  DFF_X1 DFF_1085( .CK(CK), .Q(g1842), .D(g25154) );
  DFF_X1 DFF_1086( .CK(CK), .Q(g1858), .D(g25158) );
  DFF_X1 DFF_1087( .CK(CK), .Q(g1859), .D(g25159) );
  DFF_X1 DFF_1088( .CK(CK), .Q(g1860), .D(g25160) );
  DFF_X1 DFF_1089( .CK(CK), .Q(g1861), .D(g24371) );
  DFF_X1 DFF_1090( .CK(CK), .Q(g1865), .D(g24372) );
  DFF_X1 DFF_1091( .CK(CK), .Q(g1845), .D(g24373) );
  DFF_X1 DFF_1092( .CK(CK), .Q(g1846), .D(g25155) );
  DFF_X2 DFF_1093( .CK(CK), .Q(g1849), .D(g25156) );
  DFF_X1 DFF_1094( .CK(CK), .Q(g1852), .D(g25157) );
  DFF_X1 DFF_1095( .CK(CK), .Q(g1908), .D(g16472) );
  DFF_X1 DFF_1096( .CK(CK), .Q(g1915), .D(g1908) );
  DFF_X1 DFF_1097( .CK(CK), .Q(g1922), .D(g1915) );
  DFF_X1 DFF_1098( .CK(CK), .Q(g1923), .D(g19045) );
  DFF_X1 DFF_1099( .CK(CK), .Q(g1924), .D(g1923) );
  DFF_X1 DFF_1100( .CK(CK), .Q(g1928), .D(g29445) );
  DFF_X1 DFF_1101( .CK(CK), .Q(g1929), .D(g19046) );
  DFF_X1 DFF_1102( .CK(CK), .Q(g1880), .D(g1929) );
  DFF_X1 DFF_1103( .CK(CK), .Q(g1938), .D(g19047) );
  DFF_X1 DFF_1104( .CK(CK), .Q(g1939), .D(g1938) );
  DFF_X1 DFF_1105( .CK(CK), .Q(g1956), .D(g28271) );
  DFF_X1 DFF_1106( .CK(CK), .Q(g1957), .D(g28272) );
  DFF_X1 DFF_1107( .CK(CK), .Q(g1955), .D(g28273) );
  DFF_X1 DFF_1108( .CK(CK), .Q(g1959), .D(g28274) );
  DFF_X1 DFF_1109( .CK(CK), .Q(g1960), .D(g28275) );
  DFF_X1 DFF_1110( .CK(CK), .Q(g1958), .D(g28276) );
  DFF_X1 DFF_1111( .CK(CK), .Q(g1962), .D(g28277) );
  DFF_X1 DFF_1112( .CK(CK), .Q(g1963), .D(g28278) );
  DFF_X1 DFF_1113( .CK(CK), .Q(g1961), .D(g28279) );
  DFF_X1 DFF_1114( .CK(CK), .Q(g1965), .D(g28280) );
  DFF_X1 DFF_1115( .CK(CK), .Q(g1966), .D(g28281) );
  DFF_X1 DFF_1116( .CK(CK), .Q(g1964), .D(g28282) );
  DFF_X2 DFF_1117( .CK(CK), .Q(g1967), .D(g26003) );
  DFF_X2 DFF_1118( .CK(CK), .Q(g1970), .D(g26004) );
  DFF_X1 DFF_1119( .CK(CK), .Q(g1973), .D(g26005) );
  DFF_X1 DFF_1120( .CK(CK), .Q(g1976), .D(g26006) );
  DFF_X1 DFF_1121( .CK(CK), .Q(g1979), .D(g26007) );
  DFF_X1 DFF_1122( .CK(CK), .Q(g1982), .D(g26008) );
  DFF_X1 DFF_1123( .CK(CK), .Q(g1994), .D(g29151) );
  DFF_X1 DFF_1124( .CK(CK), .Q(g1997), .D(g29152) );
  DFF_X1 DFF_1125( .CK(CK), .Q(g2000), .D(g29153) );
  DFF_X1 DFF_1126( .CK(CK), .Q(g1985), .D(g29148) );
  DFF_X1 DFF_1127( .CK(CK), .Q(g1988), .D(g29149) );
  DFF_X1 DFF_1128( .CK(CK), .Q(g1991), .D(g29150) );
  DFF_X1 DFF_1129( .CK(CK), .Q(g1871), .D(g27224) );
  DFF_X1 DFF_1130( .CK(CK), .Q(g1874), .D(g27225) );
  DFF_X1 DFF_1131( .CK(CK), .Q(g1877), .D(g27226) );
  DFF_X1 DFF_1132( .CK(CK), .Q(g1886), .D(g8302) );
  DFF_X1 DFF_1133( .CK(CK), .Q(g1887), .D(g24377) );
  DFF_X1 DFF_1134( .CK(CK), .Q(g1888), .D(g19041) );
  DFF_X1 DFF_1135( .CK(CK), .Q(g1889), .D(g19042) );
  DFF_X1 DFF_1136( .CK(CK), .Q(g1894), .D(g19043) );
  DFF_X1 DFF_1137( .CK(CK), .Q(g1895), .D(g19044) );
  DFF_X1 DFF_1138( .CK(CK), .Q(g1896), .D(g29444) );
  DFF_X1 DFF_1139( .CK(CK), .Q(g1897), .D(g29443) );
  DFF_X1 DFF_1140( .CK(CK), .Q(g1898), .D(g29442) );
  DFF_X1 DFF_1141( .CK(CK), .Q(g1899), .D(g29441) );
  DFF_X1 DFF_1142( .CK(CK), .Q(g1900), .D(g29440) );
  DFF_X1 DFF_1143( .CK(CK), .Q(g1905), .D(g1900) );
  DFF_X1 DFF_1144( .CK(CK), .Q(g1909), .D(g13442) );
  DFF_X1 DFF_1145( .CK(CK), .Q(g1910), .D(g13443) );
  DFF_X1 DFF_1146( .CK(CK), .Q(g1911), .D(g13444) );
  DFF_X1 DFF_1147( .CK(CK), .Q(g1912), .D(g13445) );
  DFF_X1 DFF_1148( .CK(CK), .Q(g1913), .D(g13446) );
  DFF_X1 DFF_1149( .CK(CK), .Q(g1914), .D(g13447) );
  DFF_X1 DFF_1150( .CK(CK), .Q(g1916), .D(g13448) );
  DFF_X1 DFF_1151( .CK(CK), .Q(g1917), .D(g13449) );
  DFF_X1 DFF_1152( .CK(CK), .Q(g1918), .D(g26002) );
  DFF_X1 DFF_1153( .CK(CK), .Q(g1921), .D(g13450) );
  DFF_X1 DFF_1154( .CK(CK), .Q(g2003), .D(g13452) );
  DFF_X1 DFF_1155( .CK(CK), .Q(g2006), .D(g2003) );
  DFF_X1 DFF_1156( .CK(CK), .Q(g2009), .D(g2006) );
  DFF_X1 DFF_1157( .CK(CK), .Q(g2010), .D(g20566) );
  DFF_X1 DFF_1158( .CK(CK), .Q(g2039), .D(g21945) );
  DFF_X1 DFF_1159( .CK(CK), .Q(g2020), .D(g23237) );
  DFF_X1 DFF_1160( .CK(CK), .Q(g2013), .D(g24378) );
  DFF_X1 DFF_1161( .CK(CK), .Q(g2033), .D(g25162) );
  DFF_X1 DFF_1162( .CK(CK), .Q(g2026), .D(g26009) );
  DFF_X1 DFF_1163( .CK(CK), .Q(g2040), .D(g26725) );
  DFF_X1 DFF_1164( .CK(CK), .Q(g2052), .D(g27227) );
  DFF_X1 DFF_1165( .CK(CK), .Q(g2046), .D(g27706) );
  DFF_X1 DFF_1166( .CK(CK), .Q(g2059), .D(g28283) );
  DFF_X1 DFF_1167( .CK(CK), .Q(g2066), .D(g28687) );
  DFF_X1 DFF_1168( .CK(CK), .Q(g2072), .D(g29154) );
  DFF_X1 DFF_1169( .CK(CK), .Q(g2079), .D(g23238) );
  DFF_X1 DFF_1170( .CK(CK), .Q(g2080), .D(g23239) );
  DFF_X1 DFF_1171( .CK(CK), .Q(g2078), .D(g23240) );
  DFF_X1 DFF_1172( .CK(CK), .Q(g2082), .D(g23241) );
  DFF_X1 DFF_1173( .CK(CK), .Q(g2083), .D(g23242) );
  DFF_X1 DFF_1174( .CK(CK), .Q(g2081), .D(g23243) );
  DFF_X1 DFF_1175( .CK(CK), .Q(g2085), .D(g23244) );
  DFF_X1 DFF_1176( .CK(CK), .Q(g2086), .D(g23245) );
  DFF_X1 DFF_1177( .CK(CK), .Q(g2084), .D(g23246) );
  DFF_X1 DFF_1178( .CK(CK), .Q(g2088), .D(g23247) );
  DFF_X1 DFF_1179( .CK(CK), .Q(g2089), .D(g23248) );
  DFF_X1 DFF_1180( .CK(CK), .Q(g2087), .D(g23249) );
  DFF_X1 DFF_1181( .CK(CK), .Q(g2091), .D(g23250) );
  DFF_X1 DFF_1182( .CK(CK), .Q(g2092), .D(g23251) );
  DFF_X1 DFF_1183( .CK(CK), .Q(g2090), .D(g23252) );
  DFF_X1 DFF_1184( .CK(CK), .Q(g2094), .D(g23253) );
  DFF_X1 DFF_1185( .CK(CK), .Q(g2095), .D(g23254) );
  DFF_X1 DFF_1186( .CK(CK), .Q(g2093), .D(g23255) );
  DFF_X1 DFF_1187( .CK(CK), .Q(g2097), .D(g23256) );
  DFF_X1 DFF_1188( .CK(CK), .Q(g2098), .D(g23257) );
  DFF_X1 DFF_1189( .CK(CK), .Q(g2096), .D(g23258) );
  DFF_X1 DFF_1190( .CK(CK), .Q(g2100), .D(g23259) );
  DFF_X1 DFF_1191( .CK(CK), .Q(g2101), .D(g23260) );
  DFF_X1 DFF_1192( .CK(CK), .Q(g2099), .D(g23261) );
  DFF_X1 DFF_1193( .CK(CK), .Q(g2103), .D(g23262) );
  DFF_X1 DFF_1194( .CK(CK), .Q(g2104), .D(g23263) );
  DFF_X2 DFF_1195( .CK(CK), .Q(g2102), .D(g23264) );
  DFF_X2 DFF_1196( .CK(CK), .Q(g2106), .D(g23265) );
  DFF_X1 DFF_1197( .CK(CK), .Q(g2107), .D(g23266) );
  DFF_X1 DFF_1198( .CK(CK), .Q(g2105), .D(g23267) );
  DFF_X1 DFF_1199( .CK(CK), .Q(g2109), .D(g23268) );
  DFF_X1 DFF_1200( .CK(CK), .Q(g2110), .D(g23269) );
  DFF_X1 DFF_1201( .CK(CK), .Q(g2108), .D(g23270) );
  DFF_X1 DFF_1202( .CK(CK), .Q(g2112), .D(g23271) );
  DFF_X1 DFF_1203( .CK(CK), .Q(g2113), .D(g23272) );
  DFF_X1 DFF_1204( .CK(CK), .Q(g2111), .D(g23273) );
  DFF_X1 DFF_1205( .CK(CK), .Q(g2115), .D(g26726) );
  DFF_X1 DFF_1206( .CK(CK), .Q(g2116), .D(g26727) );
  DFF_X1 DFF_1207( .CK(CK), .Q(g2114), .D(g26728) );
  DFF_X1 DFF_1208( .CK(CK), .Q(g2118), .D(g24379) );
  DFF_X1 DFF_1209( .CK(CK), .Q(g2119), .D(g24380) );
  DFF_X1 DFF_1210( .CK(CK), .Q(g2117), .D(g24381) );
  DFF_X1 DFF_1211( .CK(CK), .Q(g2214), .D(g13453) );
  DFF_X1 DFF_1212( .CK(CK), .Q(g2211), .D(g2214) );
  DFF_X1 DFF_1213( .CK(CK), .Q(g2241), .D(g2211) );
  DFF_X1 DFF_1214( .CK(CK), .Q(g2206), .D(g24382) );
  DFF_X1 DFF_1215( .CK(CK), .Q(g2207), .D(g24383) );
  DFF_X1 DFF_1216( .CK(CK), .Q(g2205), .D(g24384) );
  DFF_X1 DFF_1217( .CK(CK), .Q(g2209), .D(g24385) );
  DFF_X1 DFF_1218( .CK(CK), .Q(g2210), .D(g24386) );
  DFF_X1 DFF_1219( .CK(CK), .Q(g2208), .D(g24387) );
  DFF_X1 DFF_1220( .CK(CK), .Q(g2218), .D(g24388) );
  DFF_X1 DFF_1221( .CK(CK), .Q(g2219), .D(g24389) );
  DFF_X1 DFF_1222( .CK(CK), .Q(g2217), .D(g24390) );
  DFF_X1 DFF_1223( .CK(CK), .Q(g2221), .D(g24391) );
  DFF_X1 DFF_1224( .CK(CK), .Q(g2222), .D(g24392) );
  DFF_X1 DFF_1225( .CK(CK), .Q(g2220), .D(g24393) );
  DFF_X1 DFF_1226( .CK(CK), .Q(g2224), .D(g24394) );
  DFF_X1 DFF_1227( .CK(CK), .Q(g2225), .D(g24395) );
  DFF_X1 DFF_1228( .CK(CK), .Q(g2223), .D(g24396) );
  DFF_X1 DFF_1229( .CK(CK), .Q(g2227), .D(g24397) );
  DFF_X1 DFF_1230( .CK(CK), .Q(g2228), .D(g24398) );
  DFF_X1 DFF_1231( .CK(CK), .Q(g2226), .D(g24399) );
  DFF_X1 DFF_1232( .CK(CK), .Q(g2230), .D(g24400) );
  DFF_X1 DFF_1233( .CK(CK), .Q(g2231), .D(g24401) );
  DFF_X1 DFF_1234( .CK(CK), .Q(g2229), .D(g24402) );
  DFF_X1 DFF_1235( .CK(CK), .Q(g2233), .D(g24403) );
  DFF_X2 DFF_1236( .CK(CK), .Q(g2234), .D(g24404) );
  DFF_X1 DFF_1237( .CK(CK), .Q(g2232), .D(g24405) );
  DFF_X1 DFF_1238( .CK(CK), .Q(g2236), .D(g24406) );
  DFF_X1 DFF_1239( .CK(CK), .Q(g2237), .D(g24407) );
  DFF_X1 DFF_1240( .CK(CK), .Q(g2235), .D(g24408) );
  DFF_X1 DFF_1241( .CK(CK), .Q(g2239), .D(g24409) );
  DFF_X1 DFF_1242( .CK(CK), .Q(g2240), .D(g24410) );
  DFF_X1 DFF_1243( .CK(CK), .Q(g2238), .D(g24411) );
  DFF_X1 DFF_1244( .CK(CK), .Q(g2245), .D(g26730) );
  DFF_X1 DFF_1245( .CK(CK), .Q(g2246), .D(g26731) );
  DFF_X1 DFF_1246( .CK(CK), .Q(g2244), .D(g26732) );
  DFF_X1 DFF_1247( .CK(CK), .Q(g2248), .D(g26733) );
  DFF_X1 DFF_1248( .CK(CK), .Q(g2249), .D(g26734) );
  DFF_X2 DFF_1249( .CK(CK), .Q(g2247), .D(g26735) );
  DFF_X1 DFF_1250( .CK(CK), .Q(g2251), .D(g26736) );
  DFF_X1 DFF_1251( .CK(CK), .Q(g2252), .D(g26737) );
  DFF_X1 DFF_1252( .CK(CK), .Q(g2250), .D(g26738) );
  DFF_X1 DFF_1253( .CK(CK), .Q(g2254), .D(g26739) );
  DFF_X1 DFF_1254( .CK(CK), .Q(g2255), .D(g26740) );
  DFF_X1 DFF_1255( .CK(CK), .Q(g2253), .D(g26741) );
  DFF_X1 DFF_1256( .CK(CK), .Q(g2261), .D(g30551) );
  DFF_X1 DFF_1257( .CK(CK), .Q(g2264), .D(g30552) );
  DFF_X1 DFF_1258( .CK(CK), .Q(g2267), .D(g30553) );
  DFF_X1 DFF_1259( .CK(CK), .Q(g2306), .D(g30896) );
  DFF_X1 DFF_1260( .CK(CK), .Q(g2309), .D(g30897) );
  DFF_X1 DFF_1261( .CK(CK), .Q(g2312), .D(g30898) );
  DFF_X1 DFF_1262( .CK(CK), .Q(g2270), .D(g30890) );
  DFF_X1 DFF_1263( .CK(CK), .Q(g2273), .D(g30891) );
  DFF_X1 DFF_1264( .CK(CK), .Q(g2276), .D(g30892) );
  DFF_X1 DFF_1265( .CK(CK), .Q(g2315), .D(g30899) );
  DFF_X1 DFF_1266( .CK(CK), .Q(g2318), .D(g30900) );
  DFF_X1 DFF_1267( .CK(CK), .Q(g2321), .D(g30901) );
  DFF_X1 DFF_1268( .CK(CK), .Q(g2279), .D(g30554) );
  DFF_X1 DFF_1269( .CK(CK), .Q(g2282), .D(g30555) );
  DFF_X1 DFF_1270( .CK(CK), .Q(g2285), .D(g30556) );
  DFF_X1 DFF_1271( .CK(CK), .Q(g2324), .D(g30560) );
  DFF_X1 DFF_1272( .CK(CK), .Q(g2327), .D(g30561) );
  DFF_X1 DFF_1273( .CK(CK), .Q(g2330), .D(g30562) );
  DFF_X1 DFF_1274( .CK(CK), .Q(g2288), .D(g30557) );
  DFF_X1 DFF_1275( .CK(CK), .Q(g2291), .D(g30558) );
  DFF_X1 DFF_1276( .CK(CK), .Q(g2294), .D(g30559) );
  DFF_X1 DFF_1277( .CK(CK), .Q(g2333), .D(g30563) );
  DFF_X1 DFF_1278( .CK(CK), .Q(g2336), .D(g30564) );
  DFF_X1 DFF_1279( .CK(CK), .Q(g2339), .D(g30565) );
  DFF_X1 DFF_1280( .CK(CK), .Q(g2297), .D(g30893) );
  DFF_X1 DFF_1281( .CK(CK), .Q(g2300), .D(g30894) );
  DFF_X1 DFF_1282( .CK(CK), .Q(g2303), .D(g30895) );
  DFF_X1 DFF_1283( .CK(CK), .Q(g2342), .D(g30902) );
  DFF_X1 DFF_1284( .CK(CK), .Q(g2345), .D(g30903) );
  DFF_X1 DFF_1285( .CK(CK), .Q(g2348), .D(g30904) );
  DFF_X1 DFF_1286( .CK(CK), .Q(g2160), .D(g26010) );
  DFF_X1 DFF_1287( .CK(CK), .Q(g2156), .D(g26729) );
  DFF_X1 DFF_1288( .CK(CK), .Q(g2151), .D(g27228) );
  DFF_X1 DFF_1289( .CK(CK), .Q(g2147), .D(g27707) );
  DFF_X1 DFF_1290( .CK(CK), .Q(g2142), .D(g28284) );
  DFF_X1 DFF_1291( .CK(CK), .Q(g2138), .D(g28688) );
  DFF_X1 DFF_1292( .CK(CK), .Q(g2133), .D(g29155) );
  DFF_X1 DFF_1293( .CK(CK), .Q(g2129), .D(g29446) );
  DFF_X1 DFF_1294( .CK(CK), .Q(g2124), .D(g29648) );
  DFF_X1 DFF_1295( .CK(CK), .Q(g2120), .D(g29806) );
  DFF_X1 DFF_1296( .CK(CK), .Q(g2256), .D(g20567) );
  DFF_X1 DFF_1297( .CK(CK), .Q(g2258), .D(g2256) );
  DFF_X1 DFF_1298( .CK(CK), .Q(g2257), .D(g2258) );
  DFF_X1 DFF_1299( .CK(CK), .Q(g2351), .D(g13454) );
  DFF_X1 DFF_1300( .CK(CK), .Q(g2480), .D(g2351) );
  DFF_X2 DFF_1301( .CK(CK), .Q(g2476), .D(g2480) );
  DFF_X2 DFF_1302( .CK(CK), .Q(g2384), .D(g11577) );
  DFF_X2 DFF_1303( .CK(CK), .Q(g2429), .D(g28285) );
  DFF_X1 DFF_1304( .CK(CK), .Q(g2418), .D(g28286) );
  DFF_X1 DFF_1305( .CK(CK), .Q(g2421), .D(g28287) );
  DFF_X1 DFF_1306( .CK(CK), .Q(g2444), .D(g28288) );
  DFF_X1 DFF_1307( .CK(CK), .Q(g2433), .D(g28289) );
  DFF_X1 DFF_1308( .CK(CK), .Q(g2436), .D(g28290) );
  DFF_X1 DFF_1309( .CK(CK), .Q(g2459), .D(g28291) );
  DFF_X1 DFF_1310( .CK(CK), .Q(g2448), .D(g28292) );
  DFF_X1 DFF_1311( .CK(CK), .Q(g2451), .D(g28293) );
  DFF_X1 DFF_1312( .CK(CK), .Q(g2473), .D(g28294) );
  DFF_X1 DFF_1313( .CK(CK), .Q(g2463), .D(g28295) );
  DFF_X1 DFF_1314( .CK(CK), .Q(g2466), .D(g28296) );
  DFF_X1 DFF_1315( .CK(CK), .Q(g2483), .D(g29447) );
  DFF_X1 DFF_1316( .CK(CK), .Q(g2486), .D(g29448) );
  DFF_X1 DFF_1317( .CK(CK), .Q(g2489), .D(g29449) );
  DFF_X1 DFF_1318( .CK(CK), .Q(g2492), .D(g29652) );
  DFF_X1 DFF_1319( .CK(CK), .Q(g2495), .D(g29653) );
  DFF_X1 DFF_1320( .CK(CK), .Q(g2498), .D(g29654) );
  DFF_X1 DFF_1321( .CK(CK), .Q(g2502), .D(g29450) );
  DFF_X1 DFF_1322( .CK(CK), .Q(g2503), .D(g29451) );
  DFF_X1 DFF_1323( .CK(CK), .Q(g2501), .D(g29452) );
  DFF_X1 DFF_1324( .CK(CK), .Q(g2504), .D(g27708) );
  DFF_X1 DFF_1325( .CK(CK), .Q(g2507), .D(g27709) );
  DFF_X1 DFF_1326( .CK(CK), .Q(g2510), .D(g27710) );
  DFF_X1 DFF_1327( .CK(CK), .Q(g2513), .D(g27711) );
  DFF_X1 DFF_1328( .CK(CK), .Q(g2516), .D(g27712) );
  DFF_X1 DFF_1329( .CK(CK), .Q(g2519), .D(g27713) );
  DFF_X1 DFF_1330( .CK(CK), .Q(g2523), .D(g28689) );
  DFF_X1 DFF_1331( .CK(CK), .Q(g2524), .D(g28690) );
  DFF_X1 DFF_1332( .CK(CK), .Q(g2522), .D(g28691) );
  DFF_X1 DFF_1333( .CK(CK), .Q(g2387), .D(g29807) );
  DFF_X1 DFF_1334( .CK(CK), .Q(g2388), .D(g29808) );
  DFF_X1 DFF_1335( .CK(CK), .Q(g2389), .D(g29809) );
  DFF_X1 DFF_1336( .CK(CK), .Q(g2390), .D(g30905) );
  DFF_X1 DFF_1337( .CK(CK), .Q(g2391), .D(g30906) );
  DFF_X1 DFF_1338( .CK(CK), .Q(g2392), .D(g30907) );
  DFF_X1 DFF_1339( .CK(CK), .Q(g2393), .D(g30719) );
  DFF_X1 DFF_1340( .CK(CK), .Q(g2394), .D(g30720) );
  DFF_X1 DFF_1341( .CK(CK), .Q(g2395), .D(g30721) );
  DFF_X1 DFF_1342( .CK(CK), .Q(g2397), .D(g29649) );
  DFF_X1 DFF_1343( .CK(CK), .Q(g2398), .D(g29650) );
  DFF_X1 DFF_1344( .CK(CK), .Q(g2396), .D(g29651) );
  DFF_X1 DFF_1345( .CK(CK), .Q(g2478), .D(g27230) );
  DFF_X1 DFF_1346( .CK(CK), .Q(g2479), .D(g27231) );
  DFF_X1 DFF_1347( .CK(CK), .Q(g2477), .D(g27232) );
  DFF_X1 DFF_1348( .CK(CK), .Q(g2525), .D(g11590) );
  DFF_X1 DFF_1349( .CK(CK), .Q(g2526), .D(g2525) );
  DFF_X1 DFF_1350( .CK(CK), .Q(g2527), .D(g11591) );
  DFF_X1 DFF_1351( .CK(CK), .Q(g2528), .D(g2527) );
  DFF_X1 DFF_1352( .CK(CK), .Q(g2529), .D(g11592) );
  DFF_X1 DFF_1353( .CK(CK), .Q(g2354), .D(g2529) );
  DFF_X1 DFF_1354( .CK(CK), .Q(g2355), .D(g11572) );
  DFF_X1 DFF_1355( .CK(CK), .Q(g2356), .D(g2355) );
  DFF_X1 DFF_1356( .CK(CK), .Q(g2357), .D(g11573) );
  DFF_X1 DFF_1357( .CK(CK), .Q(g2358), .D(g2357) );
  DFF_X1 DFF_1358( .CK(CK), .Q(g2359), .D(g11574) );
  DFF_X1 DFF_1359( .CK(CK), .Q(g2360), .D(g2359) );
  DFF_X1 DFF_1360( .CK(CK), .Q(g2361), .D(g11575) );
  DFF_X1 DFF_1361( .CK(CK), .Q(g2362), .D(g2361) );
  DFF_X1 DFF_1362( .CK(CK), .Q(g2363), .D(g11576) );
  DFF_X1 DFF_1363( .CK(CK), .Q(g2364), .D(g2363) );
  DFF_X1 DFF_1364( .CK(CK), .Q(g2365), .D(g13455) );
  DFF_X1 DFF_1365( .CK(CK), .Q(g2366), .D(g2365) );
  DFF_X1 DFF_1366( .CK(CK), .Q(g2374), .D(g19048) );
  DFF_X1 DFF_1367( .CK(CK), .Q(g2380), .D(g30314) );
  DFF_X1 DFF_1368( .CK(CK), .Q(g2383), .D(g30315) );
  DFF_X1 DFF_1369( .CK(CK), .Q(g2372), .D(g30316) );
  DFF_X1 DFF_1370( .CK(CK), .Q(g2371), .D(g30317) );
  DFF_X1 DFF_1371( .CK(CK), .Q(g2370), .D(g30318) );
  DFF_X2 DFF_1372( .CK(CK), .Q(g2369), .D(g30319) );
  DFF_X2 DFF_1373( .CK(CK), .Q(g2379), .D(g19052) );
  DFF_X2 DFF_1374( .CK(CK), .Q(g2378), .D(g19051) );
  DFF_X1 DFF_1375( .CK(CK), .Q(g2377), .D(g19050) );
  DFF_X1 DFF_1376( .CK(CK), .Q(g2376), .D(g19049) );
  DFF_X1 DFF_1377( .CK(CK), .Q(g2375), .D(g25163) );
  DFF_X1 DFF_1378( .CK(CK), .Q(g2373), .D(g27229) );
  DFF_X1 DFF_1379( .CK(CK), .Q(g2417), .D(g11578) );
  DFF_X1 DFF_1380( .CK(CK), .Q(g2424), .D(g2417) );
  DFF_X1 DFF_1381( .CK(CK), .Q(g2425), .D(g11579) );
  DFF_X1 DFF_1382( .CK(CK), .Q(g2426), .D(g2425) );
  DFF_X1 DFF_1383( .CK(CK), .Q(g2427), .D(g11580) );
  DFF_X1 DFF_1384( .CK(CK), .Q(g2428), .D(g2427) );
  DFF_X1 DFF_1385( .CK(CK), .Q(g2432), .D(g11581) );
  DFF_X1 DFF_1386( .CK(CK), .Q(g2439), .D(g2432) );
  DFF_X1 DFF_1387( .CK(CK), .Q(g2440), .D(g11582) );
  DFF_X1 DFF_1388( .CK(CK), .Q(g2441), .D(g2440) );
  DFF_X1 DFF_1389( .CK(CK), .Q(g2442), .D(g11583) );
  DFF_X1 DFF_1390( .CK(CK), .Q(g2443), .D(g2442) );
  DFF_X1 DFF_1391( .CK(CK), .Q(g2447), .D(g11584) );
  DFF_X1 DFF_1392( .CK(CK), .Q(g2454), .D(g2447) );
  DFF_X1 DFF_1393( .CK(CK), .Q(g2455), .D(g11585) );
  DFF_X1 DFF_1394( .CK(CK), .Q(g2456), .D(g2455) );
  DFF_X1 DFF_1395( .CK(CK), .Q(g2457), .D(g11586) );
  DFF_X1 DFF_1396( .CK(CK), .Q(g2458), .D(g2457) );
  DFF_X1 DFF_1397( .CK(CK), .Q(g2462), .D(g11587) );
  DFF_X1 DFF_1398( .CK(CK), .Q(g2469), .D(g2462) );
  DFF_X1 DFF_1399( .CK(CK), .Q(g2470), .D(g11588) );
  DFF_X1 DFF_1400( .CK(CK), .Q(g2471), .D(g2470) );
  DFF_X1 DFF_1401( .CK(CK), .Q(g2472), .D(g11589) );
  DFF_X1 DFF_1402( .CK(CK), .Q(g2399), .D(g2472) );
  DFF_X1 DFF_1403( .CK(CK), .Q(g2400), .D(g13456) );
  DFF_X1 DFF_1404( .CK(CK), .Q(g2406), .D(g2400) );
  DFF_X1 DFF_1405( .CK(CK), .Q(g2412), .D(g2406) );
  DFF_X1 DFF_1406( .CK(CK), .Q(g2619), .D(g13467) );
  DFF_X1 DFF_1407( .CK(CK), .Q(g2625), .D(g2619) );
  DFF_X1 DFF_1408( .CK(CK), .Q(g2624), .D(g2625) );
  DFF_X1 DFF_1409( .CK(CK), .Q(g2628), .D(g23274) );
  DFF_X1 DFF_1410( .CK(CK), .Q(g2631), .D(g20568) );
  DFF_X1 DFF_1411( .CK(CK), .Q(g2584), .D(g20569) );
  DFF_X1 DFF_1412( .CK(CK), .Q(g2587), .D(g16473) );
  DFF_X1 DFF_1413( .CK(CK), .Q(g2597), .D(g2587) );
  DFF_X1 DFF_1414( .CK(CK), .Q(g2598), .D(g2597) );
  DFF_X1 DFF_1415( .CK(CK), .Q(g2638), .D(g11593) );
  DFF_X1 DFF_1416( .CK(CK), .Q(g2643), .D(g2638) );
  DFF_X1 DFF_1417( .CK(CK), .Q(g2644), .D(g11596) );
  DFF_X1 DFF_1418( .CK(CK), .Q(g2645), .D(g2644) );
  DFF_X1 DFF_1419( .CK(CK), .Q(g2646), .D(g11597) );
  DFF_X1 DFF_1420( .CK(CK), .Q(g2647), .D(g2646) );
  DFF_X1 DFF_1421( .CK(CK), .Q(g2648), .D(g11598) );
  DFF_X1 DFF_1422( .CK(CK), .Q(g2639), .D(g2648) );
  DFF_X1 DFF_1423( .CK(CK), .Q(g2640), .D(g11594) );
  DFF_X1 DFF_1424( .CK(CK), .Q(g2641), .D(g2640) );
  DFF_X1 DFF_1425( .CK(CK), .Q(g2642), .D(g11595) );
  DFF_X1 DFF_1426( .CK(CK), .Q(g2564), .D(g2642) );
  DFF_X1 DFF_1427( .CK(CK), .Q(g2549), .D(g13457) );
  DFF_X1 DFF_1428( .CK(CK), .Q(g2556), .D(g2549) );
  DFF_X1 DFF_1429( .CK(CK), .Q(g2560), .D(g2556) );
  DFF_X1 DFF_1430( .CK(CK), .Q(g2561), .D(g24415) );
  DFF_X1 DFF_1431( .CK(CK), .Q(g2562), .D(g24416) );
  DFF_X1 DFF_1432( .CK(CK), .Q(g2563), .D(g24417) );
  DFF_X1 DFF_1433( .CK(CK), .Q(g2530), .D(g25172) );
  DFF_X1 DFF_1434( .CK(CK), .Q(g2533), .D(g25164) );
  DFF_X1 DFF_1435( .CK(CK), .Q(g2536), .D(g25165) );
  DFF_X1 DFF_1436( .CK(CK), .Q(g2552), .D(g25169) );
  DFF_X1 DFF_1437( .CK(CK), .Q(g2553), .D(g25170) );
  DFF_X1 DFF_1438( .CK(CK), .Q(g2554), .D(g25171) );
  DFF_X1 DFF_1439( .CK(CK), .Q(g2555), .D(g24412) );
  DFF_X1 DFF_1440( .CK(CK), .Q(g2559), .D(g24413) );
  DFF_X1 DFF_1441( .CK(CK), .Q(g2539), .D(g24414) );
  DFF_X1 DFF_1442( .CK(CK), .Q(g2540), .D(g25166) );
  DFF_X1 DFF_1443( .CK(CK), .Q(g2543), .D(g25167) );
  DFF_X1 DFF_1444( .CK(CK), .Q(g2546), .D(g25168) );
  DFF_X1 DFF_1445( .CK(CK), .Q(g2602), .D(g16474) );
  DFF_X1 DFF_1446( .CK(CK), .Q(g2609), .D(g2602) );
  DFF_X1 DFF_1447( .CK(CK), .Q(g2616), .D(g2609) );
  DFF_X1 DFF_1448( .CK(CK), .Q(g2617), .D(g19057) );
  DFF_X1 DFF_1449( .CK(CK), .Q(g2618), .D(g2617) );
  DFF_X1 DFF_1450( .CK(CK), .Q(g2622), .D(g30325) );
  DFF_X1 DFF_1451( .CK(CK), .Q(g2623), .D(g19058) );
  DFF_X1 DFF_1452( .CK(CK), .Q(g2574), .D(g2623) );
  DFF_X1 DFF_1453( .CK(CK), .Q(g2632), .D(g19059) );
  DFF_X1 DFF_1454( .CK(CK), .Q(g2633), .D(g2632) );
  DFF_X1 DFF_1455( .CK(CK), .Q(g2650), .D(g28297) );
  DFF_X1 DFF_1456( .CK(CK), .Q(g2651), .D(g28298) );
  DFF_X1 DFF_1457( .CK(CK), .Q(g2649), .D(g28299) );
  DFF_X1 DFF_1458( .CK(CK), .Q(g2653), .D(g28300) );
  DFF_X1 DFF_1459( .CK(CK), .Q(g2654), .D(g28301) );
  DFF_X1 DFF_1460( .CK(CK), .Q(g2652), .D(g28302) );
  DFF_X1 DFF_1461( .CK(CK), .Q(g2656), .D(g28303) );
  DFF_X1 DFF_1462( .CK(CK), .Q(g2657), .D(g28304) );
  DFF_X1 DFF_1463( .CK(CK), .Q(g2655), .D(g28305) );
  DFF_X1 DFF_1464( .CK(CK), .Q(g2659), .D(g28306) );
  DFF_X1 DFF_1465( .CK(CK), .Q(g2660), .D(g28307) );
  DFF_X1 DFF_1466( .CK(CK), .Q(g2658), .D(g28308) );
  DFF_X1 DFF_1467( .CK(CK), .Q(g2661), .D(g26012) );
  DFF_X1 DFF_1468( .CK(CK), .Q(g2664), .D(g26013) );
  DFF_X1 DFF_1469( .CK(CK), .Q(g2667), .D(g26014) );
  DFF_X1 DFF_1470( .CK(CK), .Q(g2670), .D(g26015) );
  DFF_X1 DFF_1471( .CK(CK), .Q(g2673), .D(g26016) );
  DFF_X1 DFF_1472( .CK(CK), .Q(g2676), .D(g26017) );
  DFF_X1 DFF_1473( .CK(CK), .Q(g2688), .D(g29159) );
  DFF_X2 DFF_1474( .CK(CK), .Q(g2691), .D(g29160) );
  DFF_X2 DFF_1475( .CK(CK), .Q(g2694), .D(g29161) );
  DFF_X1 DFF_1476( .CK(CK), .Q(g2679), .D(g29156) );
  DFF_X1 DFF_1477( .CK(CK), .Q(g2682), .D(g29157) );
  DFF_X1 DFF_1478( .CK(CK), .Q(g2685), .D(g29158) );
  DFF_X1 DFF_1479( .CK(CK), .Q(g2565), .D(g27233) );
  DFF_X1 DFF_1480( .CK(CK), .Q(g2568), .D(g27234) );
  DFF_X1 DFF_1481( .CK(CK), .Q(g2571), .D(g27235) );
  DFF_X1 DFF_1482( .CK(CK), .Q(g2580), .D(g8311) );
  DFF_X1 DFF_1483( .CK(CK), .Q(g2581), .D(g24418) );
  DFF_X1 DFF_1484( .CK(CK), .Q(g2582), .D(g19053) );
  DFF_X1 DFF_1485( .CK(CK), .Q(g2583), .D(g19054) );
  DFF_X1 DFF_1486( .CK(CK), .Q(g2588), .D(g19055) );
  DFF_X1 DFF_1487( .CK(CK), .Q(g2589), .D(g19056) );
  DFF_X1 DFF_1488( .CK(CK), .Q(g2590), .D(g30324) );
  DFF_X1 DFF_1489( .CK(CK), .Q(g2591), .D(g30323) );
  DFF_X1 DFF_1490( .CK(CK), .Q(g2592), .D(g30322) );
  DFF_X1 DFF_1491( .CK(CK), .Q(g2593), .D(g30321) );
  DFF_X1 DFF_1492( .CK(CK), .Q(g2594), .D(g30320) );
  DFF_X1 DFF_1493( .CK(CK), .Q(g2599), .D(g2594) );
  DFF_X1 DFF_1494( .CK(CK), .Q(g2603), .D(g13458) );
  DFF_X1 DFF_1495( .CK(CK), .Q(g2604), .D(g13459) );
  DFF_X1 DFF_1496( .CK(CK), .Q(g2605), .D(g13460) );
  DFF_X1 DFF_1497( .CK(CK), .Q(g2606), .D(g13461) );
  DFF_X1 DFF_1498( .CK(CK), .Q(g2607), .D(g13462) );
  DFF_X1 DFF_1499( .CK(CK), .Q(g2608), .D(g13463) );
  DFF_X1 DFF_1500( .CK(CK), .Q(g2610), .D(g13464) );
  DFF_X1 DFF_1501( .CK(CK), .Q(g2611), .D(g13465) );
  DFF_X1 DFF_1502( .CK(CK), .Q(g2612), .D(g26011) );
  DFF_X1 DFF_1503( .CK(CK), .Q(g2615), .D(g13466) );
  DFF_X1 DFF_1504( .CK(CK), .Q(g2697), .D(g13468) );
  DFF_X1 DFF_1505( .CK(CK), .Q(g2700), .D(g2697) );
  DFF_X1 DFF_1506( .CK(CK), .Q(g2703), .D(g2700) );
  DFF_X1 DFF_1507( .CK(CK), .Q(g2704), .D(g20570) );
  DFF_X1 DFF_1508( .CK(CK), .Q(g2733), .D(g21946) );
  DFF_X1 DFF_1509( .CK(CK), .Q(g2714), .D(g23275) );
  DFF_X1 DFF_1510( .CK(CK), .Q(g2707), .D(g24419) );
  DFF_X1 DFF_1511( .CK(CK), .Q(g2727), .D(g25173) );
  DFF_X1 DFF_1512( .CK(CK), .Q(g2720), .D(g26018) );
  DFF_X1 DFF_1513( .CK(CK), .Q(g2734), .D(g26742) );
  DFF_X1 DFF_1514( .CK(CK), .Q(g2746), .D(g27236) );
  DFF_X1 DFF_1515( .CK(CK), .Q(g2740), .D(g27714) );
  DFF_X1 DFF_1516( .CK(CK), .Q(g2753), .D(g28309) );
  DFF_X1 DFF_1517( .CK(CK), .Q(g2760), .D(g28692) );
  DFF_X1 DFF_1518( .CK(CK), .Q(g2766), .D(g29162) );
  DFF_X1 DFF_1519( .CK(CK), .Q(g2773), .D(g23276) );
  DFF_X1 DFF_1520( .CK(CK), .Q(g2774), .D(g23277) );
  DFF_X1 DFF_1521( .CK(CK), .Q(g2772), .D(g23278) );
  DFF_X1 DFF_1522( .CK(CK), .Q(g2776), .D(g23279) );
  DFF_X1 DFF_1523( .CK(CK), .Q(g2777), .D(g23280) );
  DFF_X1 DFF_1524( .CK(CK), .Q(g2775), .D(g23281) );
  DFF_X1 DFF_1525( .CK(CK), .Q(g2779), .D(g23282) );
  DFF_X1 DFF_1526( .CK(CK), .Q(g2780), .D(g23283) );
  DFF_X1 DFF_1527( .CK(CK), .Q(g2778), .D(g23284) );
  DFF_X1 DFF_1528( .CK(CK), .Q(g2782), .D(g23285) );
  DFF_X1 DFF_1529( .CK(CK), .Q(g2783), .D(g23286) );
  DFF_X1 DFF_1530( .CK(CK), .Q(g2781), .D(g23287) );
  DFF_X1 DFF_1531( .CK(CK), .Q(g2785), .D(g23288) );
  DFF_X1 DFF_1532( .CK(CK), .Q(g2786), .D(g23289) );
  DFF_X1 DFF_1533( .CK(CK), .Q(g2784), .D(g23290) );
  DFF_X1 DFF_1534( .CK(CK), .Q(g2788), .D(g23291) );
  DFF_X1 DFF_1535( .CK(CK), .Q(g2789), .D(g23292) );
  DFF_X1 DFF_1536( .CK(CK), .Q(g2787), .D(g23293) );
  DFF_X2 DFF_1537( .CK(CK), .Q(g2791), .D(g23294) );
  DFF_X2 DFF_1538( .CK(CK), .Q(g2792), .D(g23295) );
  DFF_X2 DFF_1539( .CK(CK), .Q(g2790), .D(g23296) );
  DFF_X2 DFF_1540( .CK(CK), .Q(g2794), .D(g23297) );
  DFF_X1 DFF_1541( .CK(CK), .Q(g2795), .D(g23298) );
  DFF_X1 DFF_1542( .CK(CK), .Q(g2793), .D(g23299) );
  DFF_X1 DFF_1543( .CK(CK), .Q(g2797), .D(g23300) );
  DFF_X1 DFF_1544( .CK(CK), .Q(g2798), .D(g23301) );
  DFF_X1 DFF_1545( .CK(CK), .Q(g2796), .D(g23302) );
  DFF_X1 DFF_1546( .CK(CK), .Q(g2800), .D(g23303) );
  DFF_X1 DFF_1547( .CK(CK), .Q(g2801), .D(g23304) );
  DFF_X1 DFF_1548( .CK(CK), .Q(g2799), .D(g23305) );
  DFF_X1 DFF_1549( .CK(CK), .Q(g2803), .D(g23306) );
  DFF_X1 DFF_1550( .CK(CK), .Q(g2804), .D(g23307) );
  DFF_X1 DFF_1551( .CK(CK), .Q(g2802), .D(g23308) );
  DFF_X1 DFF_1552( .CK(CK), .Q(g2806), .D(g23309) );
  DFF_X1 DFF_1553( .CK(CK), .Q(g2807), .D(g23310) );
  DFF_X1 DFF_1554( .CK(CK), .Q(g2805), .D(g23311) );
  DFF_X1 DFF_1555( .CK(CK), .Q(g2809), .D(g26743) );
  DFF_X1 DFF_1556( .CK(CK), .Q(g2810), .D(g26744) );
  DFF_X1 DFF_1557( .CK(CK), .Q(g2808), .D(g26745) );
  DFF_X1 DFF_1558( .CK(CK), .Q(g2812), .D(g24420) );
  DFF_X1 DFF_1559( .CK(CK), .Q(g2813), .D(g24421) );
  DFF_X1 DFF_1560( .CK(CK), .Q(g2811), .D(g24422) );
  DFF_X1 DFF_1561( .CK(CK), .Q(g3054), .D(g23317) );
  DFF_X1 DFF_1562( .CK(CK), .Q(g3079), .D(g23318) );
  DFF_X1 DFF_1563( .CK(CK), .Q(g3080), .D(g21965) );
  DFF_X1 DFF_1564( .CK(CK), .Q(g3043), .D(g29453) );
  DFF_X1 DFF_1565( .CK(CK), .Q(g3044), .D(g29454) );
  DFF_X1 DFF_1566( .CK(CK), .Q(g3045), .D(g29455) );
  DFF_X1 DFF_1567( .CK(CK), .Q(g3046), .D(g29456) );
  DFF_X1 DFF_1568( .CK(CK), .Q(g3047), .D(g29457) );
  DFF_X1 DFF_1569( .CK(CK), .Q(g3048), .D(g29458) );
  DFF_X1 DFF_1570( .CK(CK), .Q(g3049), .D(g29459) );
  DFF_X1 DFF_1571( .CK(CK), .Q(g3050), .D(g29460) );
  DFF_X1 DFF_1572( .CK(CK), .Q(g3051), .D(g29655) );
  DFF_X1 DFF_1573( .CK(CK), .Q(g3052), .D(g29972) );
  DFF_X1 DFF_1574( .CK(CK), .Q(g3053), .D(g29973) );
  DFF_X1 DFF_1575( .CK(CK), .Q(g3055), .D(g29974) );
  DFF_X1 DFF_1576( .CK(CK), .Q(g3056), .D(g29975) );
  DFF_X1 DFF_1577( .CK(CK), .Q(g3057), .D(g29976) );
  DFF_X1 DFF_1578( .CK(CK), .Q(g3058), .D(g29977) );
  DFF_X1 DFF_1579( .CK(CK), .Q(g3059), .D(g29978) );
  DFF_X1 DFF_1580( .CK(CK), .Q(g3060), .D(g29979) );
  DFF_X1 DFF_1581( .CK(CK), .Q(g3061), .D(g30119) );
  DFF_X1 DFF_1582( .CK(CK), .Q(g3062), .D(g30908) );
  DFF_X1 DFF_1583( .CK(CK), .Q(g3063), .D(g30909) );
  DFF_X1 DFF_1584( .CK(CK), .Q(g3064), .D(g30910) );
  DFF_X1 DFF_1585( .CK(CK), .Q(g3065), .D(g30911) );
  DFF_X1 DFF_1586( .CK(CK), .Q(g3066), .D(g30912) );
  DFF_X1 DFF_1587( .CK(CK), .Q(g3067), .D(g30913) );
  DFF_X1 DFF_1588( .CK(CK), .Q(g3068), .D(g30914) );
  DFF_X1 DFF_1589( .CK(CK), .Q(g3069), .D(g30915) );
  DFF_X1 DFF_1590( .CK(CK), .Q(g3070), .D(g30940) );
  DFF_X1 DFF_1591( .CK(CK), .Q(g3071), .D(g30980) );
  DFF_X2 DFF_1592( .CK(CK), .Q(g3072), .D(g30981) );
  DFF_X2 DFF_1593( .CK(CK), .Q(g3073), .D(g30982) );
  DFF_X1 DFF_1594( .CK(CK), .Q(g3074), .D(g30983) );
  DFF_X1 DFF_1595( .CK(CK), .Q(g3075), .D(g30984) );
  DFF_X1 DFF_1596( .CK(CK), .Q(g3076), .D(g30985) );
  DFF_X1 DFF_1597( .CK(CK), .Q(g3077), .D(g30986) );
  DFF_X1 DFF_1598( .CK(CK), .Q(g3078), .D(g30987) );
  DFF_X1 DFF_1599( .CK(CK), .Q(g2997), .D(g30989) );
  DFF_X1 DFF_1600( .CK(CK), .Q(g2993), .D(g26748) );
  DFF_X1 DFF_1601( .CK(CK), .Q(g2998), .D(g27238) );
  DFF_X1 DFF_1602( .CK(CK), .Q(g3006), .D(g25177) );
  DFF_X1 DFF_1603( .CK(CK), .Q(g3002), .D(g26021) );
  DFF_X1 DFF_1604( .CK(CK), .Q(g3013), .D(g26750) );
  DFF_X1 DFF_1605( .CK(CK), .Q(g3010), .D(g27239) );
  DFF_X1 DFF_1606( .CK(CK), .Q(g3024), .D(g27716) );
  DFF_X1 DFF_1607( .CK(CK), .Q(g3018), .D(g24425) );
  DFF_X1 DFF_1608( .CK(CK), .Q(g3028), .D(g25176) );
  DFF_X1 DFF_1609( .CK(CK), .Q(g3036), .D(g26022) );
  DFF_X1 DFF_1610( .CK(CK), .Q(g3032), .D(g26749) );
  DFF_X1 DFF_1611( .CK(CK), .Q(g3040), .D(g16497) );
  DFF_X1 DFF_1612( .CK(CK), .Q(g2986), .D(g3040) );
  DFF_X1 DFF_1613( .CK(CK), .Q(g2987), .D(g16495) );
  DFF_X1 DFF_1614( .CK(CK), .Q(g48), .D(g20595) );
  DFF_X1 DFF_1615( .CK(CK), .Q(g45), .D(g20596) );
  DFF_X1 DFF_1616( .CK(CK), .Q(g42), .D(g20597) );
  DFF_X1 DFF_1617( .CK(CK), .Q(g39), .D(g20598) );
  DFF_X1 DFF_1618( .CK(CK), .Q(g27), .D(g20599) );
  DFF_X1 DFF_1619( .CK(CK), .Q(g30), .D(g20600) );
  DFF_X1 DFF_1620( .CK(CK), .Q(g33), .D(g20601) );
  DFF_X1 DFF_1621( .CK(CK), .Q(g36), .D(g20602) );
  DFF_X1 DFF_1622( .CK(CK), .Q(g3083), .D(g20603) );
  DFF_X1 DFF_1623( .CK(CK), .Q(g26), .D(g20604) );
  DFF_X1 DFF_1624( .CK(CK), .Q(g2992), .D(g21966) );
  DFF_X1 DFF_1625( .CK(CK), .Q(g23), .D(g20605) );
  DFF_X1 DFF_1626( .CK(CK), .Q(g20), .D(g20606) );
  DFF_X1 DFF_1627( .CK(CK), .Q(g17), .D(g20607) );
  DFF_X1 DFF_1628( .CK(CK), .Q(g11), .D(g20608) );
  DFF_X2 DFF_1629( .CK(CK), .Q(g14), .D(g20589) );
  DFF_X1 DFF_1630( .CK(CK), .Q(g5), .D(g20590) );
  DFF_X1 DFF_1631( .CK(CK), .Q(g8), .D(g20591) );
  DFF_X1 DFF_1632( .CK(CK), .Q(g2), .D(g20592) );
  DFF_X1 DFF_1633( .CK(CK), .Q(g2990), .D(g20593) );
  DFF_X1 DFF_1634( .CK(CK), .Q(g2991), .D(g21964) );
  DFF_X1 DFF_1635( .CK(CK), .Q(g1), .D(g20594) );
  INV_X1 NOT_0( .ZN(II13089), .A(g563) );
  INV_X1 NOT_1( .ZN(g562), .A(II13089) );
  INV_X1 NOT_2( .ZN(II13092), .A(g1249) );
  INV_X1 NOT_3( .ZN(g1248), .A(II13092) );
  INV_X1 NOT_4( .ZN(II13095), .A(g1943) );
  INV_X1 NOT_5( .ZN(g1942), .A(II13095) );
  INV_X1 NOT_6( .ZN(II13098), .A(g2637) );
  INV_X1 NOT_7( .ZN(g2636), .A(II13098) );
  INV_X1 NOT_8( .ZN(II13101), .A(g1) );
  INV_X1 NOT_9( .ZN(g3235), .A(II13101) );
  INV_X1 NOT_10( .ZN(II13104), .A(g2) );
  INV_X1 NOT_11( .ZN(g3236), .A(II13104) );
  INV_X1 NOT_12( .ZN(II13107), .A(g5) );
  INV_X1 NOT_13( .ZN(g3237), .A(II13107) );
  INV_X1 NOT_14( .ZN(II13110), .A(g8) );
  INV_X1 NOT_15( .ZN(g3238), .A(II13110) );
  INV_X1 NOT_16( .ZN(II13113), .A(g11) );
  INV_X1 NOT_17( .ZN(g3239), .A(II13113) );
  INV_X1 NOT_18( .ZN(II13116), .A(g14) );
  INV_X1 NOT_19( .ZN(g3240), .A(II13116) );
  INV_X1 NOT_20( .ZN(II13119), .A(g17) );
  INV_X1 NOT_21( .ZN(g3241), .A(II13119) );
  INV_X1 NOT_22( .ZN(II13122), .A(g20) );
  INV_X1 NOT_23( .ZN(g3242), .A(II13122) );
  INV_X1 NOT_24( .ZN(II13125), .A(g23) );
  INV_X1 NOT_25( .ZN(g3243), .A(II13125) );
  INV_X1 NOT_26( .ZN(II13128), .A(g26) );
  INV_X2 NOT_27( .ZN(g3244), .A(II13128) );
  INV_X2 NOT_28( .ZN(II13131), .A(g27) );
  INV_X1 NOT_29( .ZN(g3245), .A(II13131) );
  INV_X1 NOT_30( .ZN(II13134), .A(g30) );
  INV_X1 NOT_31( .ZN(g3246), .A(II13134) );
  INV_X1 NOT_32( .ZN(II13137), .A(g33) );
  INV_X1 NOT_33( .ZN(g3247), .A(II13137) );
  INV_X1 NOT_34( .ZN(II13140), .A(g36) );
  INV_X1 NOT_35( .ZN(g3248), .A(II13140) );
  INV_X1 NOT_36( .ZN(II13143), .A(g39) );
  INV_X1 NOT_37( .ZN(g3249), .A(II13143) );
  INV_X1 NOT_38( .ZN(II13146), .A(g42) );
  INV_X1 NOT_39( .ZN(g3250), .A(II13146) );
  INV_X1 NOT_40( .ZN(II13149), .A(g45) );
  INV_X1 NOT_41( .ZN(g3251), .A(II13149) );
  INV_X1 NOT_42( .ZN(II13152), .A(g48) );
  INV_X1 NOT_43( .ZN(g3252), .A(II13152) );
  INV_X1 NOT_44( .ZN(II13155), .A(g51) );
  INV_X1 NOT_45( .ZN(g3253), .A(II13155) );
  INV_X1 NOT_46( .ZN(II13158), .A(g165) );
  INV_X1 NOT_47( .ZN(g3254), .A(II13158) );
  INV_X1 NOT_48( .ZN(II13161), .A(g308) );
  INV_X1 NOT_49( .ZN(g3304), .A(II13161) );
  INV_X1 NOT_50( .ZN(g3305), .A(g305) );
  INV_X1 NOT_51( .ZN(II13165), .A(g401) );
  INV_X1 NOT_52( .ZN(g3306), .A(II13165) );
  INV_X1 NOT_53( .ZN(g3337), .A(g309) );
  INV_X1 NOT_54( .ZN(II13169), .A(g550) );
  INV_X1 NOT_55( .ZN(g3338), .A(II13169) );
  INV_X1 NOT_56( .ZN(g3365), .A(g499) );
  INV_X1 NOT_57( .ZN(II13173), .A(g629) );
  INV_X1 NOT_58( .ZN(g3366), .A(II13173) );
  INV_X1 NOT_59( .ZN(II13176), .A(g630) );
  INV_X1 NOT_60( .ZN(g3398), .A(II13176) );
  INV_X1 NOT_61( .ZN(II13179), .A(g853) );
  INV_X1 NOT_62( .ZN(g3410), .A(II13179) );
  INV_X1 NOT_63( .ZN(II13182), .A(g995) );
  INV_X1 NOT_64( .ZN(g3460), .A(II13182) );
  INV_X1 NOT_65( .ZN(g3461), .A(g992) );
  INV_X1 NOT_66( .ZN(II13186), .A(g1088) );
  INV_X1 NOT_67( .ZN(g3462), .A(II13186) );
  INV_X1 NOT_68( .ZN(g3493), .A(g996) );
  INV_X1 NOT_69( .ZN(II13190), .A(g1236) );
  INV_X1 NOT_70( .ZN(g3494), .A(II13190) );
  INV_X2 NOT_71( .ZN(g3521), .A(g1186) );
  INV_X2 NOT_72( .ZN(II13194), .A(g1315) );
  INV_X2 NOT_73( .ZN(g3522), .A(II13194) );
  INV_X1 NOT_74( .ZN(II13197), .A(g1316) );
  INV_X1 NOT_75( .ZN(g3554), .A(II13197) );
  INV_X1 NOT_76( .ZN(II13200), .A(g1547) );
  INV_X1 NOT_77( .ZN(g3566), .A(II13200) );
  INV_X1 NOT_78( .ZN(II13203), .A(g1689) );
  INV_X1 NOT_79( .ZN(g3616), .A(II13203) );
  INV_X1 NOT_80( .ZN(g3617), .A(g1686) );
  INV_X1 NOT_81( .ZN(II13207), .A(g1782) );
  INV_X1 NOT_82( .ZN(g3618), .A(II13207) );
  INV_X1 NOT_83( .ZN(g3649), .A(g1690) );
  INV_X1 NOT_84( .ZN(II13211), .A(g1930) );
  INV_X1 NOT_85( .ZN(g3650), .A(II13211) );
  INV_X1 NOT_86( .ZN(g3677), .A(g1880) );
  INV_X1 NOT_87( .ZN(II13215), .A(g2009) );
  INV_X1 NOT_88( .ZN(g3678), .A(II13215) );
  INV_X1 NOT_89( .ZN(II13218), .A(g2010) );
  INV_X1 NOT_90( .ZN(g3710), .A(II13218) );
  INV_X1 NOT_91( .ZN(II13221), .A(g2241) );
  INV_X1 NOT_92( .ZN(g3722), .A(II13221) );
  INV_X1 NOT_93( .ZN(II13224), .A(g2383) );
  INV_X1 NOT_94( .ZN(g3772), .A(II13224) );
  INV_X1 NOT_95( .ZN(g3773), .A(g2380) );
  INV_X1 NOT_96( .ZN(II13228), .A(g2476) );
  INV_X1 NOT_97( .ZN(g3774), .A(II13228) );
  INV_X1 NOT_98( .ZN(g3805), .A(g2384) );
  INV_X1 NOT_99( .ZN(II13232), .A(g2624) );
  INV_X1 NOT_100( .ZN(g3806), .A(II13232) );
  INV_X1 NOT_101( .ZN(g3833), .A(g2574) );
  INV_X1 NOT_102( .ZN(II13236), .A(g2703) );
  INV_X1 NOT_103( .ZN(g3834), .A(II13236) );
  INV_X1 NOT_104( .ZN(II13239), .A(g2704) );
  INV_X1 NOT_105( .ZN(g3866), .A(II13239) );
  INV_X1 NOT_106( .ZN(II13242), .A(g2879) );
  INV_X1 NOT_107( .ZN(g3878), .A(II13242) );
  INV_X1 NOT_108( .ZN(g3897), .A(g2950) );
  INV_X1 NOT_109( .ZN(II13246), .A(g2987) );
  INV_X1 NOT_110( .ZN(g3900), .A(II13246) );
  INV_X1 NOT_111( .ZN(g3919), .A(g3080) );
  INV_X1 NOT_112( .ZN(g3922), .A(g150) );
  INV_X1 NOT_113( .ZN(g3925), .A(g155) );
  INV_X1 NOT_114( .ZN(g3928), .A(g157) );
  INV_X1 NOT_115( .ZN(g3931), .A(g171) );
  INV_X1 NOT_116( .ZN(g3934), .A(g176) );
  INV_X1 NOT_117( .ZN(g3937), .A(g178) );
  INV_X1 NOT_118( .ZN(g3940), .A(g408) );
  INV_X1 NOT_119( .ZN(g3941), .A(g455) );
  INV_X1 NOT_120( .ZN(g3942), .A(g699) );
  INV_X1 NOT_121( .ZN(g3945), .A(g726) );
  INV_X1 NOT_122( .ZN(g3948), .A(g835) );
  INV_X1 NOT_123( .ZN(g3951), .A(g840) );
  INV_X1 NOT_124( .ZN(g3954), .A(g842) );
  INV_X1 NOT_125( .ZN(g3957), .A(g856) );
  INV_X1 NOT_126( .ZN(g3960), .A(g861) );
  INV_X1 NOT_127( .ZN(g3963), .A(g863) );
  INV_X1 NOT_128( .ZN(g3966), .A(g1526) );
  INV_X1 NOT_129( .ZN(g3969), .A(g1531) );
  INV_X1 NOT_130( .ZN(g3972), .A(g1533) );
  INV_X1 NOT_131( .ZN(g3975), .A(g1552) );
  INV_X1 NOT_132( .ZN(g3978), .A(g1554) );
  INV_X1 NOT_133( .ZN(g3981), .A(g2217) );
  INV_X1 NOT_134( .ZN(g3984), .A(g2222) );
  INV_X2 NOT_135( .ZN(g3987), .A(g2224) );
  INV_X2 NOT_136( .ZN(g3990), .A(g2245) );
  INV_X2 NOT_137( .ZN(II13275), .A(g2848) );
  INV_X1 NOT_138( .ZN(g3993), .A(II13275) );
  INV_X1 NOT_139( .ZN(g3994), .A(g2848) );
  INV_X1 NOT_140( .ZN(g3995), .A(g3064) );
  INV_X1 NOT_141( .ZN(g3996), .A(g3073) );
  INV_X1 NOT_142( .ZN(g3997), .A(g45) );
  INV_X1 NOT_143( .ZN(g3998), .A(g23) );
  INV_X1 NOT_144( .ZN(g3999), .A(g3204) );
  INV_X1 NOT_145( .ZN(g4000), .A(g153) );
  INV_X1 NOT_146( .ZN(g4003), .A(g158) );
  INV_X1 NOT_147( .ZN(g4006), .A(g160) );
  INV_X1 NOT_148( .ZN(g4009), .A(g174) );
  INV_X1 NOT_149( .ZN(g4012), .A(g179) );
  INV_X1 NOT_150( .ZN(g4015), .A(g411) );
  INV_X1 NOT_151( .ZN(g4016), .A(g417) );
  INV_X1 NOT_152( .ZN(g4017), .A(g427) );
  INV_X1 NOT_153( .ZN(g4020), .A(g700) );
  INV_X1 NOT_154( .ZN(g4023), .A(g702) );
  INV_X1 NOT_155( .ZN(g4026), .A(g727) );
  INV_X1 NOT_156( .ZN(g4029), .A(g838) );
  INV_X1 NOT_157( .ZN(g4032), .A(g843) );
  INV_X1 NOT_158( .ZN(g4035), .A(g845) );
  INV_X1 NOT_159( .ZN(g4038), .A(g859) );
  INV_X1 NOT_160( .ZN(g4041), .A(g864) );
  INV_X1 NOT_161( .ZN(g4044), .A(g866) );
  INV_X1 NOT_162( .ZN(g4047), .A(g1095) );
  INV_X1 NOT_163( .ZN(g4048), .A(g1142) );
  INV_X1 NOT_164( .ZN(g4049), .A(g1385) );
  INV_X1 NOT_165( .ZN(g4052), .A(g1412) );
  INV_X1 NOT_166( .ZN(g4055), .A(g1529) );
  INV_X1 NOT_167( .ZN(g4058), .A(g1534) );
  INV_X1 NOT_168( .ZN(g4061), .A(g1536) );
  INV_X1 NOT_169( .ZN(g4064), .A(g1550) );
  INV_X1 NOT_170( .ZN(g4067), .A(g1555) );
  INV_X1 NOT_171( .ZN(g4070), .A(g1557) );
  INV_X1 NOT_172( .ZN(g4073), .A(g2220) );
  INV_X1 NOT_173( .ZN(g4076), .A(g2225) );
  INV_X1 NOT_174( .ZN(g4079), .A(g2227) );
  INV_X1 NOT_175( .ZN(g4082), .A(g2246) );
  INV_X1 NOT_176( .ZN(g4085), .A(g2248) );
  INV_X1 NOT_177( .ZN(II13316), .A(g2836) );
  INV_X1 NOT_178( .ZN(g4088), .A(II13316) );
  INV_X1 NOT_179( .ZN(g4089), .A(g2836) );
  INV_X1 NOT_180( .ZN(II13320), .A(g2864) );
  INV_X1 NOT_181( .ZN(g4090), .A(II13320) );
  INV_X1 NOT_182( .ZN(g4091), .A(g2864) );
  INV_X1 NOT_183( .ZN(g4092), .A(g3074) );
  INV_X1 NOT_184( .ZN(g4093), .A(g33) );
  INV_X4 NOT_185( .ZN(g4094), .A(g3207) );
  INV_X4 NOT_186( .ZN(g4095), .A(g130) );
  INV_X4 NOT_187( .ZN(g4098), .A(g156) );
  INV_X1 NOT_188( .ZN(g4101), .A(g161) );
  INV_X1 NOT_189( .ZN(g4104), .A(g163) );
  INV_X1 NOT_190( .ZN(g4107), .A(g177) );
  INV_X1 NOT_191( .ZN(g4110), .A(g414) );
  INV_X1 NOT_192( .ZN(g4111), .A(g420) );
  INV_X1 NOT_193( .ZN(g4112), .A(g428) );
  INV_X1 NOT_194( .ZN(g4115), .A(g698) );
  INV_X1 NOT_195( .ZN(g4118), .A(g703) );
  INV_X1 NOT_196( .ZN(g4121), .A(g705) );
  INV_X1 NOT_197( .ZN(g4124), .A(g725) );
  INV_X1 NOT_198( .ZN(g4127), .A(g841) );
  INV_X1 NOT_199( .ZN(g4130), .A(g846) );
  INV_X1 NOT_200( .ZN(g4133), .A(g848) );
  INV_X1 NOT_201( .ZN(g4136), .A(g862) );
  INV_X1 NOT_202( .ZN(g4139), .A(g867) );
  INV_X1 NOT_203( .ZN(g4142), .A(g1098) );
  INV_X1 NOT_204( .ZN(g4143), .A(g1104) );
  INV_X1 NOT_205( .ZN(g4144), .A(g1114) );
  INV_X1 NOT_206( .ZN(g4147), .A(g1386) );
  INV_X1 NOT_207( .ZN(g4150), .A(g1388) );
  INV_X1 NOT_208( .ZN(g4153), .A(g1413) );
  INV_X1 NOT_209( .ZN(g4156), .A(g1532) );
  INV_X1 NOT_210( .ZN(g4159), .A(g1537) );
  INV_X1 NOT_211( .ZN(g4162), .A(g1539) );
  INV_X1 NOT_212( .ZN(g4165), .A(g1553) );
  INV_X1 NOT_213( .ZN(g4168), .A(g1558) );
  INV_X1 NOT_214( .ZN(g4171), .A(g1560) );
  INV_X1 NOT_215( .ZN(g4174), .A(g1789) );
  INV_X1 NOT_216( .ZN(g4175), .A(g1836) );
  INV_X1 NOT_217( .ZN(g4176), .A(g2079) );
  INV_X1 NOT_218( .ZN(g4179), .A(g2106) );
  INV_X1 NOT_219( .ZN(g4182), .A(g2223) );
  INV_X1 NOT_220( .ZN(g4185), .A(g2228) );
  INV_X1 NOT_221( .ZN(g4188), .A(g2230) );
  INV_X1 NOT_222( .ZN(g4191), .A(g2244) );
  INV_X1 NOT_223( .ZN(g4194), .A(g2249) );
  INV_X1 NOT_224( .ZN(g4197), .A(g2251) );
  INV_X1 NOT_225( .ZN(II13366), .A(g2851) );
  INV_X1 NOT_226( .ZN(g4200), .A(II13366) );
  INV_X1 NOT_227( .ZN(g4201), .A(g2851) );
  INV_X1 NOT_228( .ZN(g4202), .A(g42) );
  INV_X1 NOT_229( .ZN(g4203), .A(g20) );
  INV_X1 NOT_230( .ZN(g4204), .A(g3188) );
  INV_X1 NOT_231( .ZN(g4205), .A(g131) );
  INV_X1 NOT_232( .ZN(g4208), .A(g133) );
  INV_X1 NOT_233( .ZN(g4211), .A(g159) );
  INV_X1 NOT_234( .ZN(g4214), .A(g164) );
  INV_X1 NOT_235( .ZN(g4217), .A(g354) );
  INV_X1 NOT_236( .ZN(g4220), .A(g423) );
  INV_X1 NOT_237( .ZN(g4221), .A(g426) );
  INV_X1 NOT_238( .ZN(g4224), .A(g429) );
  INV_X1 NOT_239( .ZN(g4225), .A(g701) );
  INV_X1 NOT_240( .ZN(g4228), .A(g706) );
  INV_X1 NOT_241( .ZN(g4231), .A(g708) );
  INV_X1 NOT_242( .ZN(g4234), .A(g818) );
  INV_X1 NOT_243( .ZN(g4237), .A(g844) );
  INV_X1 NOT_244( .ZN(g4240), .A(g849) );
  INV_X1 NOT_245( .ZN(g4243), .A(g851) );
  INV_X1 NOT_246( .ZN(g4246), .A(g865) );
  INV_X1 NOT_247( .ZN(g4249), .A(g1101) );
  INV_X1 NOT_248( .ZN(g4250), .A(g1107) );
  INV_X1 NOT_249( .ZN(g4251), .A(g1115) );
  INV_X1 NOT_250( .ZN(g4254), .A(g1384) );
  INV_X1 NOT_251( .ZN(g4257), .A(g1389) );
  INV_X1 NOT_252( .ZN(g4260), .A(g1391) );
  INV_X1 NOT_253( .ZN(g4263), .A(g1411) );
  INV_X4 NOT_254( .ZN(g4266), .A(g1535) );
  INV_X4 NOT_255( .ZN(g4269), .A(g1540) );
  INV_X4 NOT_256( .ZN(g4272), .A(g1542) );
  INV_X1 NOT_257( .ZN(g4275), .A(g1556) );
  INV_X1 NOT_258( .ZN(g4278), .A(g1561) );
  INV_X1 NOT_259( .ZN(g4281), .A(g1792) );
  INV_X1 NOT_260( .ZN(g4282), .A(g1798) );
  INV_X1 NOT_261( .ZN(g4283), .A(g1808) );
  INV_X1 NOT_262( .ZN(g4286), .A(g2080) );
  INV_X1 NOT_263( .ZN(g4289), .A(g2082) );
  INV_X1 NOT_264( .ZN(g4292), .A(g2107) );
  INV_X1 NOT_265( .ZN(g4295), .A(g2226) );
  INV_X1 NOT_266( .ZN(g4298), .A(g2231) );
  INV_X1 NOT_267( .ZN(g4301), .A(g2233) );
  INV_X1 NOT_268( .ZN(g4304), .A(g2247) );
  INV_X1 NOT_269( .ZN(g4307), .A(g2252) );
  INV_X1 NOT_270( .ZN(g4310), .A(g2254) );
  INV_X1 NOT_271( .ZN(g4313), .A(g2483) );
  INV_X1 NOT_272( .ZN(g4314), .A(g2530) );
  INV_X1 NOT_273( .ZN(g4315), .A(g2773) );
  INV_X1 NOT_274( .ZN(g4318), .A(g2800) );
  INV_X1 NOT_275( .ZN(II13417), .A(g2839) );
  INV_X1 NOT_276( .ZN(g4321), .A(II13417) );
  INV_X1 NOT_277( .ZN(g4322), .A(g2839) );
  INV_X1 NOT_278( .ZN(II13421), .A(g2867) );
  INV_X1 NOT_279( .ZN(g4323), .A(II13421) );
  INV_X1 NOT_280( .ZN(g4324), .A(g2867) );
  INV_X1 NOT_281( .ZN(g4325), .A(g36) );
  INV_X1 NOT_282( .ZN(g4326), .A(g181) );
  INV_X1 NOT_283( .ZN(g4329), .A(g129) );
  INV_X1 NOT_284( .ZN(g4332), .A(g134) );
  INV_X1 NOT_285( .ZN(g4335), .A(g162) );
  INV_X1 NOT_286( .ZN(II13430), .A(g101) );
  INV_X1 NOT_287( .ZN(g4338), .A(II13430) );
  INV_X1 NOT_288( .ZN(II13433), .A(g105) );
  INV_X1 NOT_289( .ZN(g4339), .A(II13433) );
  INV_X1 NOT_290( .ZN(g4340), .A(g343) );
  INV_X1 NOT_291( .ZN(g4343), .A(g369) );
  INV_X1 NOT_292( .ZN(g4346), .A(g432) );
  INV_X1 NOT_293( .ZN(g4347), .A(g438) );
  INV_X1 NOT_294( .ZN(g4348), .A(g704) );
  INV_X1 NOT_295( .ZN(g4351), .A(g709) );
  INV_X1 NOT_296( .ZN(g4354), .A(g711) );
  INV_X1 NOT_297( .ZN(g4357), .A(g729) );
  INV_X1 NOT_298( .ZN(g4360), .A(g819) );
  INV_X1 NOT_299( .ZN(g4363), .A(g821) );
  INV_X1 NOT_300( .ZN(g4366), .A(g847) );
  INV_X1 NOT_301( .ZN(g4369), .A(g852) );
  INV_X1 NOT_302( .ZN(g4372), .A(g1041) );
  INV_X1 NOT_303( .ZN(g4375), .A(g1110) );
  INV_X1 NOT_304( .ZN(g4376), .A(g1113) );
  INV_X1 NOT_305( .ZN(g4379), .A(g1116) );
  INV_X1 NOT_306( .ZN(g4380), .A(g1387) );
  INV_X8 NOT_307( .ZN(g4383), .A(g1392) );
  INV_X8 NOT_308( .ZN(g4386), .A(g1394) );
  INV_X1 NOT_309( .ZN(g4389), .A(g1512) );
  INV_X1 NOT_310( .ZN(g4392), .A(g1538) );
  INV_X1 NOT_311( .ZN(g4395), .A(g1543) );
  INV_X1 NOT_312( .ZN(g4398), .A(g1545) );
  INV_X1 NOT_313( .ZN(g4401), .A(g1559) );
  INV_X1 NOT_314( .ZN(g4404), .A(g1795) );
  INV_X1 NOT_315( .ZN(g4405), .A(g1801) );
  INV_X1 NOT_316( .ZN(g4406), .A(g1809) );
  INV_X1 NOT_317( .ZN(g4409), .A(g2078) );
  INV_X1 NOT_318( .ZN(g4412), .A(g2083) );
  INV_X1 NOT_319( .ZN(g4415), .A(g2085) );
  INV_X1 NOT_320( .ZN(g4418), .A(g2105) );
  INV_X1 NOT_321( .ZN(g4421), .A(g2229) );
  INV_X1 NOT_322( .ZN(g4424), .A(g2234) );
  INV_X1 NOT_323( .ZN(g4427), .A(g2236) );
  INV_X1 NOT_324( .ZN(g4430), .A(g2250) );
  INV_X1 NOT_325( .ZN(g4433), .A(g2255) );
  INV_X1 NOT_326( .ZN(g4436), .A(g2486) );
  INV_X1 NOT_327( .ZN(g4437), .A(g2492) );
  INV_X1 NOT_328( .ZN(g4438), .A(g2502) );
  INV_X1 NOT_329( .ZN(g4441), .A(g2774) );
  INV_X1 NOT_330( .ZN(g4444), .A(g2776) );
  INV_X1 NOT_331( .ZN(g4447), .A(g2801) );
  INV_X1 NOT_332( .ZN(II13478), .A(g2854) );
  INV_X1 NOT_333( .ZN(g4450), .A(II13478) );
  INV_X1 NOT_334( .ZN(g4451), .A(g2854) );
  INV_X1 NOT_335( .ZN(g4452), .A(g17) );
  INV_X1 NOT_336( .ZN(g4453), .A(g132) );
  INV_X1 NOT_337( .ZN(g4456), .A(g309) );
  INV_X1 NOT_338( .ZN(g4465), .A(g346) );
  INV_X1 NOT_339( .ZN(g4468), .A(g358) );
  INV_X1 NOT_340( .ZN(g4471), .A(g384) );
  INV_X1 NOT_341( .ZN(g4474), .A(g435) );
  INV_X1 NOT_342( .ZN(g4475), .A(g441) );
  INV_X1 NOT_343( .ZN(g4476), .A(g576) );
  INV_X1 NOT_344( .ZN(g4479), .A(g587) );
  INV_X1 NOT_345( .ZN(g4480), .A(g707) );
  INV_X1 NOT_346( .ZN(g4483), .A(g712) );
  INV_X1 NOT_347( .ZN(g4486), .A(g714) );
  INV_X1 NOT_348( .ZN(g4489), .A(g730) );
  INV_X1 NOT_349( .ZN(g4492), .A(g732) );
  INV_X1 NOT_350( .ZN(g4495), .A(g869) );
  INV_X1 NOT_351( .ZN(g4498), .A(g817) );
  INV_X1 NOT_352( .ZN(g4501), .A(g822) );
  INV_X1 NOT_353( .ZN(g4504), .A(g850) );
  INV_X1 NOT_354( .ZN(II13501), .A(g789) );
  INV_X1 NOT_355( .ZN(g4507), .A(II13501) );
  INV_X1 NOT_356( .ZN(II13504), .A(g793) );
  INV_X1 NOT_357( .ZN(g4508), .A(II13504) );
  INV_X1 NOT_358( .ZN(g4509), .A(g1030) );
  INV_X1 NOT_359( .ZN(g4512), .A(g1056) );
  INV_X1 NOT_360( .ZN(g4515), .A(g1119) );
  INV_X1 NOT_361( .ZN(g4516), .A(g1125) );
  INV_X1 NOT_362( .ZN(g4517), .A(g1390) );
  INV_X1 NOT_363( .ZN(g4520), .A(g1395) );
  INV_X1 NOT_364( .ZN(g4523), .A(g1397) );
  INV_X1 NOT_365( .ZN(g4526), .A(g1415) );
  INV_X8 NOT_366( .ZN(g4529), .A(g1513) );
  INV_X1 NOT_367( .ZN(g4532), .A(g1515) );
  INV_X1 NOT_368( .ZN(g4535), .A(g1541) );
  INV_X1 NOT_369( .ZN(g4538), .A(g1546) );
  INV_X1 NOT_370( .ZN(g4541), .A(g1735) );
  INV_X1 NOT_371( .ZN(g4544), .A(g1804) );
  INV_X1 NOT_372( .ZN(g4545), .A(g1807) );
  INV_X1 NOT_373( .ZN(g4548), .A(g1810) );
  INV_X1 NOT_374( .ZN(g4549), .A(g2081) );
  INV_X1 NOT_375( .ZN(g4552), .A(g2086) );
  INV_X1 NOT_376( .ZN(g4555), .A(g2088) );
  INV_X1 NOT_377( .ZN(g4558), .A(g2206) );
  INV_X1 NOT_378( .ZN(g4561), .A(g2232) );
  INV_X1 NOT_379( .ZN(g4564), .A(g2237) );
  INV_X1 NOT_380( .ZN(g4567), .A(g2239) );
  INV_X1 NOT_381( .ZN(g4570), .A(g2253) );
  INV_X1 NOT_382( .ZN(g4573), .A(g2489) );
  INV_X1 NOT_383( .ZN(g4574), .A(g2495) );
  INV_X1 NOT_384( .ZN(g4575), .A(g2503) );
  INV_X1 NOT_385( .ZN(g4578), .A(g2772) );
  INV_X1 NOT_386( .ZN(g4581), .A(g2777) );
  INV_X1 NOT_387( .ZN(g4584), .A(g2779) );
  INV_X1 NOT_388( .ZN(g4587), .A(g2799) );
  INV_X1 NOT_389( .ZN(II13538), .A(g2870) );
  INV_X1 NOT_390( .ZN(g4590), .A(II13538) );
  INV_X1 NOT_391( .ZN(g4591), .A(g2870) );
  INV_X1 NOT_392( .ZN(g4592), .A(g361) );
  INV_X1 NOT_393( .ZN(g4595), .A(g373) );
  INV_X1 NOT_394( .ZN(g4598), .A(g398) );
  INV_X1 NOT_395( .ZN(g4601), .A(g444) );
  INV_X1 NOT_396( .ZN(g4602), .A(g525) );
  INV_X1 NOT_397( .ZN(g4603), .A(g577) );
  INV_X1 NOT_398( .ZN(g4606), .A(g579) );
  INV_X1 NOT_399( .ZN(g4609), .A(g590) );
  INV_X1 NOT_400( .ZN(g4610), .A(g596) );
  INV_X1 NOT_401( .ZN(g4611), .A(g710) );
  INV_X1 NOT_402( .ZN(g4614), .A(g715) );
  INV_X1 NOT_403( .ZN(g4617), .A(g717) );
  INV_X1 NOT_404( .ZN(g4620), .A(g728) );
  INV_X1 NOT_405( .ZN(g4623), .A(g733) );
  INV_X1 NOT_406( .ZN(g4626), .A(g735) );
  INV_X1 NOT_407( .ZN(g4629), .A(g820) );
  INV_X1 NOT_408( .ZN(g4632), .A(g996) );
  INV_X1 NOT_409( .ZN(g4641), .A(g1033) );
  INV_X1 NOT_410( .ZN(g4644), .A(g1045) );
  INV_X1 NOT_411( .ZN(g4647), .A(g1071) );
  INV_X1 NOT_412( .ZN(g4650), .A(g1122) );
  INV_X1 NOT_413( .ZN(g4651), .A(g1128) );
  INV_X1 NOT_414( .ZN(g4652), .A(g1262) );
  INV_X1 NOT_415( .ZN(g4655), .A(g1273) );
  INV_X1 NOT_416( .ZN(g4656), .A(g1393) );
  INV_X1 NOT_417( .ZN(g4659), .A(g1398) );
  INV_X1 NOT_418( .ZN(g4662), .A(g1400) );
  INV_X1 NOT_419( .ZN(g4665), .A(g1416) );
  INV_X1 NOT_420( .ZN(g4668), .A(g1418) );
  INV_X1 NOT_421( .ZN(g4671), .A(g1563) );
  INV_X8 NOT_422( .ZN(g4674), .A(g1511) );
  INV_X8 NOT_423( .ZN(g4677), .A(g1516) );
  INV_X1 NOT_424( .ZN(g4680), .A(g1544) );
  INV_X1 NOT_425( .ZN(II13575), .A(g1476) );
  INV_X1 NOT_426( .ZN(g4683), .A(II13575) );
  INV_X1 NOT_427( .ZN(II13578), .A(g1481) );
  INV_X1 NOT_428( .ZN(g4684), .A(II13578) );
  INV_X1 NOT_429( .ZN(g4685), .A(g1724) );
  INV_X1 NOT_430( .ZN(g4688), .A(g1750) );
  INV_X1 NOT_431( .ZN(g4691), .A(g1813) );
  INV_X1 NOT_432( .ZN(g4692), .A(g1819) );
  INV_X1 NOT_433( .ZN(g4693), .A(g2084) );
  INV_X1 NOT_434( .ZN(g4696), .A(g2089) );
  INV_X1 NOT_435( .ZN(g4699), .A(g2091) );
  INV_X1 NOT_436( .ZN(g4702), .A(g2109) );
  INV_X1 NOT_437( .ZN(g4705), .A(g2207) );
  INV_X1 NOT_438( .ZN(g4708), .A(g2209) );
  INV_X1 NOT_439( .ZN(g4711), .A(g2235) );
  INV_X1 NOT_440( .ZN(g4714), .A(g2240) );
  INV_X1 NOT_441( .ZN(g4717), .A(g2429) );
  INV_X1 NOT_442( .ZN(g4720), .A(g2498) );
  INV_X1 NOT_443( .ZN(g4721), .A(g2501) );
  INV_X1 NOT_444( .ZN(g4724), .A(g2504) );
  INV_X1 NOT_445( .ZN(g4725), .A(g2775) );
  INV_X1 NOT_446( .ZN(g4728), .A(g2780) );
  INV_X1 NOT_447( .ZN(g4731), .A(g2782) );
  INV_X1 NOT_448( .ZN(g4734), .A(g11) );
  INV_X1 NOT_449( .ZN(II13601), .A(g121) );
  INV_X1 NOT_450( .ZN(g4735), .A(II13601) );
  INV_X1 NOT_451( .ZN(II13604), .A(g125) );
  INV_X1 NOT_452( .ZN(g4736), .A(II13604) );
  INV_X1 NOT_453( .ZN(g4737), .A(g376) );
  INV_X1 NOT_454( .ZN(g4740), .A(g388) );
  INV_X1 NOT_455( .ZN(g4743), .A(g575) );
  INV_X1 NOT_456( .ZN(g4746), .A(g580) );
  INV_X1 NOT_457( .ZN(g4749), .A(g582) );
  INV_X1 NOT_458( .ZN(g4752), .A(g593) );
  INV_X1 NOT_459( .ZN(g4753), .A(g599) );
  INV_X1 NOT_460( .ZN(g4754), .A(g713) );
  INV_X1 NOT_461( .ZN(g4757), .A(g718) );
  INV_X1 NOT_462( .ZN(g4760), .A(g720) );
  INV_X1 NOT_463( .ZN(g4763), .A(g731) );
  INV_X1 NOT_464( .ZN(g4766), .A(g736) );
  INV_X1 NOT_465( .ZN(g4769), .A(g1048) );
  INV_X1 NOT_466( .ZN(g4772), .A(g1060) );
  INV_X1 NOT_467( .ZN(g4775), .A(g1085) );
  INV_X1 NOT_468( .ZN(g4778), .A(g1131) );
  INV_X1 NOT_469( .ZN(g4779), .A(g1211) );
  INV_X1 NOT_470( .ZN(g4780), .A(g1263) );
  INV_X1 NOT_471( .ZN(g4783), .A(g1265) );
  INV_X1 NOT_472( .ZN(g4786), .A(g1276) );
  INV_X1 NOT_473( .ZN(g4787), .A(g1282) );
  INV_X1 NOT_474( .ZN(g4788), .A(g1396) );
  INV_X1 NOT_475( .ZN(g4791), .A(g1401) );
  INV_X1 NOT_476( .ZN(g4794), .A(g1403) );
  INV_X1 NOT_477( .ZN(g4797), .A(g1414) );
  INV_X1 NOT_478( .ZN(g4800), .A(g1419) );
  INV_X1 NOT_479( .ZN(g4803), .A(g1421) );
  INV_X1 NOT_480( .ZN(g4806), .A(g1514) );
  INV_X1 NOT_481( .ZN(g4809), .A(g1690) );
  INV_X1 NOT_482( .ZN(g4818), .A(g1727) );
  INV_X1 NOT_483( .ZN(g4821), .A(g1739) );
  INV_X1 NOT_484( .ZN(g4824), .A(g1765) );
  INV_X1 NOT_485( .ZN(g4827), .A(g1816) );
  INV_X1 NOT_486( .ZN(g4828), .A(g1822) );
  INV_X1 NOT_487( .ZN(g4829), .A(g1956) );
  INV_X1 NOT_488( .ZN(g4832), .A(g1967) );
  INV_X1 NOT_489( .ZN(g4833), .A(g2087) );
  INV_X1 NOT_490( .ZN(g4836), .A(g2092) );
  INV_X1 NOT_491( .ZN(g4839), .A(g2094) );
  INV_X1 NOT_492( .ZN(g4842), .A(g2110) );
  INV_X1 NOT_493( .ZN(g4845), .A(g2112) );
  INV_X1 NOT_494( .ZN(g4848), .A(g2257) );
  INV_X1 NOT_495( .ZN(g4851), .A(g2205) );
  INV_X1 NOT_496( .ZN(g4854), .A(g2210) );
  INV_X1 NOT_497( .ZN(g4857), .A(g2238) );
  INV_X1 NOT_498( .ZN(II13652), .A(g2170) );
  INV_X1 NOT_499( .ZN(g4860), .A(II13652) );
  INV_X1 NOT_500( .ZN(II13655), .A(g2175) );
  INV_X1 NOT_501( .ZN(g4861), .A(II13655) );
  INV_X1 NOT_502( .ZN(g4862), .A(g2418) );
  INV_X1 NOT_503( .ZN(g4865), .A(g2444) );
  INV_X1 NOT_504( .ZN(g4868), .A(g2507) );
  INV_X1 NOT_505( .ZN(g4869), .A(g2513) );
  INV_X1 NOT_506( .ZN(g4870), .A(g2778) );
  INV_X1 NOT_507( .ZN(g4873), .A(g2783) );
  INV_X1 NOT_508( .ZN(g4876), .A(g2785) );
  INV_X1 NOT_509( .ZN(g4879), .A(g2803) );
  INV_X1 NOT_510( .ZN(g4882), .A(g391) );
  INV_X1 NOT_511( .ZN(g4885), .A(g448) );
  INV_X1 NOT_512( .ZN(g4888), .A(g578) );
  INV_X1 NOT_513( .ZN(g4891), .A(g583) );
  INV_X1 NOT_514( .ZN(g4894), .A(g585) );
  INV_X1 NOT_515( .ZN(g4897), .A(g602) );
  INV_X1 NOT_516( .ZN(g4898), .A(g605) );
  INV_X1 NOT_517( .ZN(g4899), .A(g716) );
  INV_X1 NOT_518( .ZN(g4902), .A(g721) );
  INV_X1 NOT_519( .ZN(g4905), .A(g723) );
  INV_X1 NOT_520( .ZN(g4908), .A(g734) );
  INV_X1 NOT_521( .ZN(II13677), .A(g809) );
  INV_X1 NOT_522( .ZN(g4911), .A(II13677) );
  INV_X1 NOT_523( .ZN(II13680), .A(g813) );
  INV_X1 NOT_524( .ZN(g4912), .A(II13680) );
  INV_X1 NOT_525( .ZN(g4913), .A(g1063) );
  INV_X1 NOT_526( .ZN(g4916), .A(g1075) );
  INV_X1 NOT_527( .ZN(g4919), .A(g1261) );
  INV_X1 NOT_528( .ZN(g4922), .A(g1266) );
  INV_X1 NOT_529( .ZN(g4925), .A(g1268) );
  INV_X1 NOT_530( .ZN(g4928), .A(g1279) );
  INV_X1 NOT_531( .ZN(g4929), .A(g1285) );
  INV_X1 NOT_532( .ZN(g4930), .A(g1399) );
  INV_X1 NOT_533( .ZN(g4933), .A(g1404) );
  INV_X1 NOT_534( .ZN(g4936), .A(g1406) );
  INV_X8 NOT_535( .ZN(g4939), .A(g1417) );
  INV_X8 NOT_536( .ZN(g4942), .A(g1422) );
  INV_X8 NOT_537( .ZN(g4945), .A(g1742) );
  INV_X8 NOT_538( .ZN(g4948), .A(g1754) );
  INV_X1 NOT_539( .ZN(g4951), .A(g1779) );
  INV_X1 NOT_540( .ZN(g4954), .A(g1825) );
  INV_X1 NOT_541( .ZN(g4955), .A(g1905) );
  INV_X1 NOT_542( .ZN(g4956), .A(g1957) );
  INV_X1 NOT_543( .ZN(g4959), .A(g1959) );
  INV_X1 NOT_544( .ZN(g4962), .A(g1970) );
  INV_X1 NOT_545( .ZN(g4963), .A(g1976) );
  INV_X1 NOT_546( .ZN(g4964), .A(g2090) );
  INV_X1 NOT_547( .ZN(g4967), .A(g2095) );
  INV_X1 NOT_548( .ZN(g4970), .A(g2097) );
  INV_X1 NOT_549( .ZN(g4973), .A(g2108) );
  INV_X1 NOT_550( .ZN(g4976), .A(g2113) );
  INV_X1 NOT_551( .ZN(g4979), .A(g2115) );
  INV_X1 NOT_552( .ZN(g4982), .A(g2208) );
  INV_X1 NOT_553( .ZN(g4985), .A(g2384) );
  INV_X1 NOT_554( .ZN(g4994), .A(g2421) );
  INV_X1 NOT_555( .ZN(g4997), .A(g2433) );
  INV_X1 NOT_556( .ZN(g5000), .A(g2459) );
  INV_X1 NOT_557( .ZN(g5003), .A(g2510) );
  INV_X1 NOT_558( .ZN(g5004), .A(g2516) );
  INV_X1 NOT_559( .ZN(g5005), .A(g2650) );
  INV_X1 NOT_560( .ZN(g5008), .A(g2661) );
  INV_X1 NOT_561( .ZN(g5009), .A(g2781) );
  INV_X1 NOT_562( .ZN(g5012), .A(g2786) );
  INV_X1 NOT_563( .ZN(g5015), .A(g2788) );
  INV_X1 NOT_564( .ZN(g5018), .A(g2804) );
  INV_X1 NOT_565( .ZN(g5021), .A(g2806) );
  INV_X1 NOT_566( .ZN(g5024), .A(g449) );
  INV_X1 NOT_567( .ZN(g5027), .A(g581) );
  INV_X1 NOT_568( .ZN(g5030), .A(g586) );
  INV_X1 NOT_569( .ZN(g5033), .A(g608) );
  INV_X1 NOT_570( .ZN(g5034), .A(g614) );
  INV_X1 NOT_571( .ZN(g5035), .A(g719) );
  INV_X1 NOT_572( .ZN(g5038), .A(g724) );
  INV_X1 NOT_573( .ZN(g5041), .A(g1078) );
  INV_X1 NOT_574( .ZN(g5044), .A(g1135) );
  INV_X1 NOT_575( .ZN(g5047), .A(g1264) );
  INV_X1 NOT_576( .ZN(g5050), .A(g1269) );
  INV_X1 NOT_577( .ZN(g5053), .A(g1271) );
  INV_X1 NOT_578( .ZN(g5056), .A(g1288) );
  INV_X1 NOT_579( .ZN(g5057), .A(g1291) );
  INV_X1 NOT_580( .ZN(g5058), .A(g1402) );
  INV_X1 NOT_581( .ZN(g5061), .A(g1407) );
  INV_X1 NOT_582( .ZN(g5064), .A(g1409) );
  INV_X1 NOT_583( .ZN(g5067), .A(g1420) );
  INV_X1 NOT_584( .ZN(II13742), .A(g1501) );
  INV_X1 NOT_585( .ZN(g5070), .A(II13742) );
  INV_X1 NOT_586( .ZN(II13745), .A(g1506) );
  INV_X1 NOT_587( .ZN(g5071), .A(II13745) );
  INV_X1 NOT_588( .ZN(g5072), .A(g1757) );
  INV_X1 NOT_589( .ZN(g5075), .A(g1769) );
  INV_X1 NOT_590( .ZN(g5078), .A(g1955) );
  INV_X1 NOT_591( .ZN(g5081), .A(g1960) );
  INV_X1 NOT_592( .ZN(g5084), .A(g1962) );
  INV_X1 NOT_593( .ZN(g5087), .A(g1973) );
  INV_X1 NOT_594( .ZN(g5088), .A(g1979) );
  INV_X1 NOT_595( .ZN(g5089), .A(g2093) );
  INV_X1 NOT_596( .ZN(g5092), .A(g2098) );
  INV_X1 NOT_597( .ZN(g5095), .A(g2100) );
  INV_X1 NOT_598( .ZN(g5098), .A(g2111) );
  INV_X1 NOT_599( .ZN(g5101), .A(g2116) );
  INV_X1 NOT_600( .ZN(g5104), .A(g2436) );
  INV_X1 NOT_601( .ZN(g5107), .A(g2448) );
  INV_X1 NOT_602( .ZN(g5110), .A(g2473) );
  INV_X1 NOT_603( .ZN(g5113), .A(g2519) );
  INV_X16 NOT_604( .ZN(g5114), .A(g2599) );
  INV_X1 NOT_605( .ZN(g5115), .A(g2651) );
  INV_X1 NOT_606( .ZN(g5118), .A(g2653) );
  INV_X1 NOT_607( .ZN(g5121), .A(g2664) );
  INV_X1 NOT_608( .ZN(g5122), .A(g2670) );
  INV_X1 NOT_609( .ZN(g5123), .A(g2784) );
  INV_X1 NOT_610( .ZN(g5126), .A(g2789) );
  INV_X1 NOT_611( .ZN(g5129), .A(g2791) );
  INV_X1 NOT_612( .ZN(g5132), .A(g2802) );
  INV_X1 NOT_613( .ZN(g5135), .A(g2807) );
  INV_X1 NOT_614( .ZN(g5138), .A(g2809) );
  INV_X1 NOT_615( .ZN(II13775), .A(g109) );
  INV_X1 NOT_616( .ZN(g5141), .A(II13775) );
  INV_X1 NOT_617( .ZN(g5142), .A(g447) );
  INV_X1 NOT_618( .ZN(g5145), .A(g584) );
  INV_X1 NOT_619( .ZN(g5148), .A(g611) );
  INV_X1 NOT_620( .ZN(g5149), .A(g617) );
  INV_X1 NOT_621( .ZN(g5150), .A(g722) );
  INV_X1 NOT_622( .ZN(g5153), .A(g1136) );
  INV_X1 NOT_623( .ZN(g5156), .A(g1267) );
  INV_X1 NOT_624( .ZN(g5159), .A(g1272) );
  INV_X1 NOT_625( .ZN(g5162), .A(g1294) );
  INV_X1 NOT_626( .ZN(g5163), .A(g1300) );
  INV_X1 NOT_627( .ZN(g5164), .A(g1405) );
  INV_X1 NOT_628( .ZN(g5167), .A(g1410) );
  INV_X1 NOT_629( .ZN(g5170), .A(g1772) );
  INV_X1 NOT_630( .ZN(g5173), .A(g1829) );
  INV_X1 NOT_631( .ZN(g5176), .A(g1958) );
  INV_X1 NOT_632( .ZN(g5179), .A(g1963) );
  INV_X1 NOT_633( .ZN(g5182), .A(g1965) );
  INV_X1 NOT_634( .ZN(g5185), .A(g1982) );
  INV_X1 NOT_635( .ZN(g5186), .A(g1985) );
  INV_X1 NOT_636( .ZN(g5187), .A(g2096) );
  INV_X1 NOT_637( .ZN(g5190), .A(g2101) );
  INV_X1 NOT_638( .ZN(g5193), .A(g2103) );
  INV_X1 NOT_639( .ZN(g5196), .A(g2114) );
  INV_X1 NOT_640( .ZN(II13801), .A(g2195) );
  INV_X1 NOT_641( .ZN(g5199), .A(II13801) );
  INV_X1 NOT_642( .ZN(II13804), .A(g2200) );
  INV_X1 NOT_643( .ZN(g5200), .A(II13804) );
  INV_X1 NOT_644( .ZN(g5201), .A(g2451) );
  INV_X1 NOT_645( .ZN(g5204), .A(g2463) );
  INV_X1 NOT_646( .ZN(g5207), .A(g2649) );
  INV_X1 NOT_647( .ZN(g5210), .A(g2654) );
  INV_X1 NOT_648( .ZN(g5213), .A(g2656) );
  INV_X1 NOT_649( .ZN(g5216), .A(g2667) );
  INV_X1 NOT_650( .ZN(g5217), .A(g2673) );
  INV_X1 NOT_651( .ZN(g5218), .A(g2787) );
  INV_X1 NOT_652( .ZN(g5221), .A(g2792) );
  INV_X1 NOT_653( .ZN(g5224), .A(g2794) );
  INV_X1 NOT_654( .ZN(g5227), .A(g2805) );
  INV_X1 NOT_655( .ZN(g5230), .A(g2810) );
  INV_X1 NOT_656( .ZN(g5233), .A(g620) );
  INV_X1 NOT_657( .ZN(II13820), .A(g797) );
  INV_X1 NOT_658( .ZN(g5234), .A(II13820) );
  INV_X1 NOT_659( .ZN(g5235), .A(g1134) );
  INV_X1 NOT_660( .ZN(g5238), .A(g1270) );
  INV_X1 NOT_661( .ZN(g5241), .A(g1297) );
  INV_X1 NOT_662( .ZN(g5242), .A(g1303) );
  INV_X1 NOT_663( .ZN(g5243), .A(g1408) );
  INV_X1 NOT_664( .ZN(g5246), .A(g1830) );
  INV_X1 NOT_665( .ZN(g5249), .A(g1961) );
  INV_X1 NOT_666( .ZN(g5252), .A(g1966) );
  INV_X16 NOT_667( .ZN(g5255), .A(g1988) );
  INV_X1 NOT_668( .ZN(g5256), .A(g1994) );
  INV_X1 NOT_669( .ZN(g5257), .A(g2099) );
  INV_X1 NOT_670( .ZN(g5260), .A(g2104) );
  INV_X1 NOT_671( .ZN(g5263), .A(g2466) );
  INV_X1 NOT_672( .ZN(g5266), .A(g2523) );
  INV_X1 NOT_673( .ZN(g5269), .A(g2652) );
  INV_X1 NOT_674( .ZN(g5272), .A(g2657) );
  INV_X1 NOT_675( .ZN(g5275), .A(g2659) );
  INV_X1 NOT_676( .ZN(g5278), .A(g2676) );
  INV_X1 NOT_677( .ZN(g5279), .A(g2679) );
  INV_X1 NOT_678( .ZN(g5280), .A(g2790) );
  INV_X1 NOT_679( .ZN(g5283), .A(g2795) );
  INV_X1 NOT_680( .ZN(g5286), .A(g2797) );
  INV_X1 NOT_681( .ZN(g5289), .A(g2808) );
  INV_X1 NOT_682( .ZN(g5292), .A(g2857) );
  INV_X1 NOT_683( .ZN(g5293), .A(g738) );
  INV_X1 NOT_684( .ZN(g5296), .A(g1306) );
  INV_X1 NOT_685( .ZN(II13849), .A(g1486) );
  INV_X1 NOT_686( .ZN(g5297), .A(II13849) );
  INV_X1 NOT_687( .ZN(g5298), .A(g1828) );
  INV_X1 NOT_688( .ZN(g5301), .A(g1964) );
  INV_X1 NOT_689( .ZN(g5304), .A(g1991) );
  INV_X1 NOT_690( .ZN(g5305), .A(g1997) );
  INV_X1 NOT_691( .ZN(g5306), .A(g2102) );
  INV_X1 NOT_692( .ZN(g5309), .A(g2524) );
  INV_X1 NOT_693( .ZN(g5312), .A(g2655) );
  INV_X1 NOT_694( .ZN(g5315), .A(g2660) );
  INV_X1 NOT_695( .ZN(g5318), .A(g2682) );
  INV_X1 NOT_696( .ZN(g5319), .A(g2688) );
  INV_X1 NOT_697( .ZN(g5320), .A(g2793) );
  INV_X1 NOT_698( .ZN(g5323), .A(g2798) );
  INV_X1 NOT_699( .ZN(g5326), .A(g2873) );
  INV_X1 NOT_700( .ZN(g5327), .A(g739) );
  INV_X1 NOT_701( .ZN(g5330), .A(g1424) );
  INV_X1 NOT_702( .ZN(g5333), .A(g2000) );
  INV_X1 NOT_703( .ZN(II13868), .A(g2180) );
  INV_X1 NOT_704( .ZN(g5334), .A(II13868) );
  INV_X1 NOT_705( .ZN(g5335), .A(g2522) );
  INV_X1 NOT_706( .ZN(g5338), .A(g2658) );
  INV_X1 NOT_707( .ZN(g5341), .A(g2685) );
  INV_X1 NOT_708( .ZN(g5342), .A(g2691) );
  INV_X16 NOT_709( .ZN(g5343), .A(g2796) );
  INV_X1 NOT_710( .ZN(g5346), .A(g3106) );
  INV_X1 NOT_711( .ZN(g5349), .A(g2877) );
  INV_X1 NOT_712( .ZN(g5352), .A(g737) );
  INV_X1 NOT_713( .ZN(g5355), .A(g1425) );
  INV_X1 NOT_714( .ZN(g5358), .A(g2118) );
  INV_X1 NOT_715( .ZN(g5361), .A(g2694) );
  INV_X1 NOT_716( .ZN(g5362), .A(g2817) );
  INV_X1 NOT_717( .ZN(g5363), .A(g3107) );
  INV_X1 NOT_718( .ZN(g5366), .A(g2878) );
  INV_X1 NOT_719( .ZN(g5369), .A(g1423) );
  INV_X1 NOT_720( .ZN(g5372), .A(g2119) );
  INV_X1 NOT_721( .ZN(g5375), .A(g2812) );
  INV_X1 NOT_722( .ZN(g5378), .A(g2933) );
  INV_X1 NOT_723( .ZN(g5379), .A(g3108) );
  INV_X1 NOT_724( .ZN(g5382), .A(g2117) );
  INV_X1 NOT_725( .ZN(g5385), .A(g2813) );
  INV_X1 NOT_726( .ZN(II13892), .A(g3040) );
  INV_X1 NOT_727( .ZN(g5388), .A(II13892) );
  INV_X1 NOT_728( .ZN(g5389), .A(g3040) );
  INV_X1 NOT_729( .ZN(II13896), .A(g343) );
  INV_X1 NOT_730( .ZN(g5390), .A(II13896) );
  INV_X1 NOT_731( .ZN(g5391), .A(g2811) );
  INV_X1 NOT_732( .ZN(g5394), .A(g3054) );
  INV_X1 NOT_733( .ZN(II13901), .A(g346) );
  INV_X1 NOT_734( .ZN(g5395), .A(II13901) );
  INV_X1 NOT_735( .ZN(II13904), .A(g358) );
  INV_X1 NOT_736( .ZN(g5396), .A(II13904) );
  INV_X1 NOT_737( .ZN(II13907), .A(g1030) );
  INV_X1 NOT_738( .ZN(g5397), .A(II13907) );
  INV_X1 NOT_739( .ZN(II13910), .A(g361) );
  INV_X1 NOT_740( .ZN(g5398), .A(II13910) );
  INV_X1 NOT_741( .ZN(II13913), .A(g373) );
  INV_X1 NOT_742( .ZN(g5399), .A(II13913) );
  INV_X1 NOT_743( .ZN(II13916), .A(g1033) );
  INV_X1 NOT_744( .ZN(g5400), .A(II13916) );
  INV_X1 NOT_745( .ZN(II13919), .A(g1045) );
  INV_X1 NOT_746( .ZN(g5401), .A(II13919) );
  INV_X1 NOT_747( .ZN(II13922), .A(g1724) );
  INV_X1 NOT_748( .ZN(g5402), .A(II13922) );
  INV_X1 NOT_749( .ZN(II13925), .A(g376) );
  INV_X1 NOT_750( .ZN(g5403), .A(II13925) );
  INV_X1 NOT_751( .ZN(II13928), .A(g388) );
  INV_X1 NOT_752( .ZN(g5404), .A(II13928) );
  INV_X1 NOT_753( .ZN(II13931), .A(g1048) );
  INV_X1 NOT_754( .ZN(g5405), .A(II13931) );
  INV_X1 NOT_755( .ZN(II13934), .A(g1060) );
  INV_X1 NOT_756( .ZN(g5406), .A(II13934) );
  INV_X1 NOT_757( .ZN(II13937), .A(g1727) );
  INV_X1 NOT_758( .ZN(g5407), .A(II13937) );
  INV_X1 NOT_759( .ZN(II13940), .A(g1739) );
  INV_X1 NOT_760( .ZN(g5408), .A(II13940) );
  INV_X1 NOT_761( .ZN(II13943), .A(g2418) );
  INV_X1 NOT_762( .ZN(g5409), .A(II13943) );
  INV_X1 NOT_763( .ZN(g5410), .A(g3079) );
  INV_X1 NOT_764( .ZN(II13947), .A(g391) );
  INV_X1 NOT_765( .ZN(g5411), .A(II13947) );
  INV_X1 NOT_766( .ZN(II13950), .A(g1063) );
  INV_X1 NOT_767( .ZN(g5412), .A(II13950) );
  INV_X1 NOT_768( .ZN(II13953), .A(g1075) );
  INV_X1 NOT_769( .ZN(g5413), .A(II13953) );
  INV_X1 NOT_770( .ZN(II13956), .A(g1742) );
  INV_X1 NOT_771( .ZN(g5414), .A(II13956) );
  INV_X1 NOT_772( .ZN(II13959), .A(g1754) );
  INV_X1 NOT_773( .ZN(g5415), .A(II13959) );
  INV_X1 NOT_774( .ZN(II13962), .A(g2421) );
  INV_X1 NOT_775( .ZN(g5416), .A(II13962) );
  INV_X1 NOT_776( .ZN(II13965), .A(g2433) );
  INV_X1 NOT_777( .ZN(g5417), .A(II13965) );
  INV_X1 NOT_778( .ZN(II13968), .A(g1078) );
  INV_X1 NOT_779( .ZN(g5418), .A(II13968) );
  INV_X1 NOT_780( .ZN(II13971), .A(g1757) );
  INV_X1 NOT_781( .ZN(g5419), .A(II13971) );
  INV_X1 NOT_782( .ZN(II13974), .A(g1769) );
  INV_X1 NOT_783( .ZN(g5420), .A(II13974) );
  INV_X1 NOT_784( .ZN(II13977), .A(g2436) );
  INV_X1 NOT_785( .ZN(g5421), .A(II13977) );
  INV_X1 NOT_786( .ZN(II13980), .A(g2448) );
  INV_X1 NOT_787( .ZN(g5422), .A(II13980) );
  INV_X1 NOT_788( .ZN(g5423), .A(g2879) );
  INV_X1 NOT_789( .ZN(II13984), .A(g1772) );
  INV_X1 NOT_790( .ZN(g5424), .A(II13984) );
  INV_X1 NOT_791( .ZN(II13987), .A(g2451) );
  INV_X1 NOT_792( .ZN(g5425), .A(II13987) );
  INV_X1 NOT_793( .ZN(II13990), .A(g2463) );
  INV_X1 NOT_794( .ZN(g5426), .A(II13990) );
  INV_X1 NOT_795( .ZN(II13993), .A(g2466) );
  INV_X1 NOT_796( .ZN(g5427), .A(II13993) );
  INV_X1 NOT_797( .ZN(g5428), .A(g3210) );
  INV_X1 NOT_798( .ZN(g5431), .A(g3211) );
  INV_X1 NOT_799( .ZN(g5434), .A(g3084) );
  INV_X1 NOT_800( .ZN(II13999), .A(g276) );
  INV_X1 NOT_801( .ZN(g5437), .A(II13999) );
  INV_X1 NOT_802( .ZN(II14002), .A(g276) );
  INV_X1 NOT_803( .ZN(g5438), .A(II14002) );
  INV_X1 NOT_804( .ZN(g5469), .A(g3085) );
  INV_X1 NOT_805( .ZN(II14006), .A(g963) );
  INV_X1 NOT_806( .ZN(g5472), .A(II14006) );
  INV_X1 NOT_807( .ZN(II14009), .A(g963) );
  INV_X1 NOT_808( .ZN(g5473), .A(II14009) );
  INV_X1 NOT_809( .ZN(g5504), .A(g3086) );
  INV_X1 NOT_810( .ZN(g5507), .A(g3155) );
  INV_X1 NOT_811( .ZN(II14014), .A(g499) );
  INV_X1 NOT_812( .ZN(g5508), .A(II14014) );
  INV_X1 NOT_813( .ZN(II14017), .A(g1657) );
  INV_X1 NOT_814( .ZN(g5511), .A(II14017) );
  INV_X1 NOT_815( .ZN(II14020), .A(g1657) );
  INV_X1 NOT_816( .ZN(g5512), .A(II14020) );
  INV_X1 NOT_817( .ZN(g5543), .A(g3087) );
  INV_X1 NOT_818( .ZN(g5546), .A(g3164) );
  INV_X1 NOT_819( .ZN(g5547), .A(g101) );
  INV_X1 NOT_820( .ZN(g5548), .A(g105) );
  INV_X1 NOT_821( .ZN(II14027), .A(g182) );
  INV_X1 NOT_822( .ZN(g5549), .A(II14027) );
  INV_X1 NOT_823( .ZN(II14030), .A(g182) );
  INV_X1 NOT_824( .ZN(g5550), .A(II14030) );
  INV_X1 NOT_825( .ZN(g5551), .A(g514) );
  INV_X1 NOT_826( .ZN(II14034), .A(g1186) );
  INV_X1 NOT_827( .ZN(g5552), .A(II14034) );
  INV_X1 NOT_828( .ZN(II14037), .A(g2351) );
  INV_X1 NOT_829( .ZN(g5555), .A(II14037) );
  INV_X1 NOT_830( .ZN(II14040), .A(g2351) );
  INV_X1 NOT_831( .ZN(g5556), .A(II14040) );
  INV_X1 NOT_832( .ZN(g5587), .A(g3091) );
  INV_X1 NOT_833( .ZN(g5590), .A(g3158) );
  INV_X1 NOT_834( .ZN(g5591), .A(g3173) );
  INV_X1 NOT_835( .ZN(g5592), .A(g515) );
  INV_X1 NOT_836( .ZN(g5593), .A(g789) );
  INV_X1 NOT_837( .ZN(g5594), .A(g793) );
  INV_X1 NOT_838( .ZN(II14049), .A(g870) );
  INV_X1 NOT_839( .ZN(g5595), .A(II14049) );
  INV_X1 NOT_840( .ZN(II14052), .A(g870) );
  INV_X1 NOT_841( .ZN(g5596), .A(II14052) );
  INV_X1 NOT_842( .ZN(g5597), .A(g1200) );
  INV_X16 NOT_843( .ZN(II14056), .A(g1880) );
  INV_X1 NOT_844( .ZN(g5598), .A(II14056) );
  INV_X1 NOT_845( .ZN(g5601), .A(g3092) );
  INV_X1 NOT_846( .ZN(g5604), .A(g3167) );
  INV_X1 NOT_847( .ZN(g5605), .A(g3182) );
  INV_X1 NOT_848( .ZN(g5606), .A(g79) );
  INV_X1 NOT_849( .ZN(g5609), .A(g1201) );
  INV_X1 NOT_850( .ZN(g5610), .A(g1476) );
  INV_X1 NOT_851( .ZN(g5611), .A(g1481) );
  INV_X1 NOT_852( .ZN(II14066), .A(g1564) );
  INV_X1 NOT_853( .ZN(g5612), .A(II14066) );
  INV_X1 NOT_854( .ZN(II14069), .A(g1564) );
  INV_X1 NOT_855( .ZN(g5613), .A(II14069) );
  INV_X1 NOT_856( .ZN(g5614), .A(g1894) );
  INV_X1 NOT_857( .ZN(II14073), .A(g2574) );
  INV_X1 NOT_858( .ZN(g5615), .A(II14073) );
  INV_X1 NOT_859( .ZN(g5618), .A(g3093) );
  INV_X1 NOT_860( .ZN(g5621), .A(g3161) );
  INV_X1 NOT_861( .ZN(g5622), .A(g3176) );
  INV_X1 NOT_862( .ZN(g5623), .A(g70) );
  INV_X1 NOT_863( .ZN(g5626), .A(g121) );
  INV_X1 NOT_864( .ZN(g5627), .A(g125) );
  INV_X1 NOT_865( .ZN(g5628), .A(g300) );
  INV_X1 NOT_866( .ZN(II14083), .A(g325) );
  INV_X1 NOT_867( .ZN(g5629), .A(II14083) );
  INV_X1 NOT_868( .ZN(g5631), .A(g767) );
  INV_X1 NOT_869( .ZN(g5634), .A(g1895) );
  INV_X1 NOT_870( .ZN(g5635), .A(g2170) );
  INV_X1 NOT_871( .ZN(g5636), .A(g2175) );
  INV_X1 NOT_872( .ZN(II14091), .A(g2258) );
  INV_X1 NOT_873( .ZN(g5637), .A(II14091) );
  INV_X1 NOT_874( .ZN(II14094), .A(g2258) );
  INV_X1 NOT_875( .ZN(g5638), .A(II14094) );
  INV_X1 NOT_876( .ZN(g5639), .A(g2588) );
  INV_X1 NOT_877( .ZN(g5640), .A(g3170) );
  INV_X1 NOT_878( .ZN(g5641), .A(g3185) );
  INV_X1 NOT_879( .ZN(g5642), .A(g61) );
  INV_X1 NOT_880( .ZN(g5645), .A(g101) );
  INV_X1 NOT_881( .ZN(g5646), .A(g213) );
  INV_X1 NOT_882( .ZN(g5647), .A(g301) );
  INV_X1 NOT_883( .ZN(II14104), .A(g331) );
  INV_X1 NOT_884( .ZN(g5648), .A(II14104) );
  INV_X1 NOT_885( .ZN(g5651), .A(g758) );
  INV_X1 NOT_886( .ZN(g5654), .A(g809) );
  INV_X1 NOT_887( .ZN(g5655), .A(g813) );
  INV_X1 NOT_888( .ZN(g5656), .A(g987) );
  INV_X1 NOT_889( .ZN(II14113), .A(g1012) );
  INV_X1 NOT_890( .ZN(g5657), .A(II14113) );
  INV_X1 NOT_891( .ZN(g5659), .A(g1453) );
  INV_X1 NOT_892( .ZN(g5662), .A(g2589) );
  INV_X1 NOT_893( .ZN(g5663), .A(g3179) );
  INV_X1 NOT_894( .ZN(g5664), .A(g65) );
  INV_X1 NOT_895( .ZN(g5665), .A(g105) );
  INV_X1 NOT_896( .ZN(g5666), .A(g216) );
  INV_X1 NOT_897( .ZN(g5667), .A(g222) );
  INV_X1 NOT_898( .ZN(g5668), .A(g299) );
  INV_X1 NOT_899( .ZN(g5675), .A(g302) );
  INV_X1 NOT_900( .ZN(g5679), .A(g506) );
  INV_X1 NOT_901( .ZN(g5680), .A(g749) );
  INV_X1 NOT_902( .ZN(g5683), .A(g789) );
  INV_X1 NOT_903( .ZN(g5684), .A(g900) );
  INV_X1 NOT_904( .ZN(g5685), .A(g988) );
  INV_X1 NOT_905( .ZN(II14134), .A(g1018) );
  INV_X1 NOT_906( .ZN(g5686), .A(II14134) );
  INV_X1 NOT_907( .ZN(g5689), .A(g1444) );
  INV_X1 NOT_908( .ZN(g5692), .A(g1501) );
  INV_X1 NOT_909( .ZN(g5693), .A(g1506) );
  INV_X1 NOT_910( .ZN(g5694), .A(g1681) );
  INV_X1 NOT_911( .ZN(II14143), .A(g1706) );
  INV_X1 NOT_912( .ZN(g5695), .A(II14143) );
  INV_X1 NOT_913( .ZN(g5697), .A(g2147) );
  INV_X1 NOT_914( .ZN(g5700), .A(g3088) );
  INV_X1 NOT_915( .ZN(II14149), .A(g3231) );
  INV_X1 NOT_916( .ZN(g5701), .A(II14149) );
  INV_X1 NOT_917( .ZN(g5702), .A(g56) );
  INV_X1 NOT_918( .ZN(g5703), .A(g109) );
  INV_X1 NOT_919( .ZN(g5704), .A(g219) );
  INV_X1 NOT_920( .ZN(g5705), .A(g225) );
  INV_X1 NOT_921( .ZN(g5706), .A(g231) );
  INV_X1 NOT_922( .ZN(g5707), .A(g109) );
  INV_X1 NOT_923( .ZN(g5708), .A(g303) );
  INV_X1 NOT_924( .ZN(g5712), .A(g305) );
  INV_X1 NOT_925( .ZN(II14163), .A(g113) );
  INV_X1 NOT_926( .ZN(g5713), .A(II14163) );
  INV_X1 NOT_927( .ZN(g5714), .A(g507) );
  INV_X1 NOT_928( .ZN(g5715), .A(g541) );
  INV_X1 NOT_929( .ZN(g5716), .A(g753) );
  INV_X1 NOT_930( .ZN(g5717), .A(g793) );
  INV_X1 NOT_931( .ZN(g5718), .A(g903) );
  INV_X1 NOT_932( .ZN(g5719), .A(g909) );
  INV_X1 NOT_933( .ZN(g5720), .A(g986) );
  INV_X1 NOT_934( .ZN(g5727), .A(g989) );
  INV_X1 NOT_935( .ZN(g5731), .A(g1192) );
  INV_X8 NOT_936( .ZN(g5732), .A(g1435) );
  INV_X8 NOT_937( .ZN(g5735), .A(g1476) );
  INV_X1 NOT_938( .ZN(g5736), .A(g1594) );
  INV_X1 NOT_939( .ZN(g5737), .A(g1682) );
  INV_X1 NOT_940( .ZN(II14182), .A(g1712) );
  INV_X1 NOT_941( .ZN(g5738), .A(II14182) );
  INV_X1 NOT_942( .ZN(g5741), .A(g2138) );
  INV_X1 NOT_943( .ZN(g5744), .A(g2195) );
  INV_X1 NOT_944( .ZN(g5745), .A(g2200) );
  INV_X1 NOT_945( .ZN(g5746), .A(g2375) );
  INV_X1 NOT_946( .ZN(II14191), .A(g2400) );
  INV_X1 NOT_947( .ZN(g5747), .A(II14191) );
  INV_X1 NOT_948( .ZN(II14195), .A(g3212) );
  INV_X1 NOT_949( .ZN(g5749), .A(II14195) );
  INV_X1 NOT_950( .ZN(g5750), .A(g92) );
  INV_X1 NOT_951( .ZN(g5751), .A(g52) );
  INV_X1 NOT_952( .ZN(g5752), .A(g113) );
  INV_X1 NOT_953( .ZN(g5753), .A(g228) );
  INV_X1 NOT_954( .ZN(g5754), .A(g234) );
  INV_X1 NOT_955( .ZN(g5755), .A(g240) );
  INV_X1 NOT_956( .ZN(g5756), .A(g304) );
  INV_X1 NOT_957( .ZN(g5759), .A(g508) );
  INV_X1 NOT_958( .ZN(g5760), .A(g744) );
  INV_X1 NOT_959( .ZN(g5761), .A(g797) );
  INV_X1 NOT_960( .ZN(g5762), .A(g906) );
  INV_X1 NOT_961( .ZN(g5763), .A(g912) );
  INV_X1 NOT_962( .ZN(g5764), .A(g918) );
  INV_X1 NOT_963( .ZN(g5765), .A(g797) );
  INV_X1 NOT_964( .ZN(g5766), .A(g990) );
  INV_X1 NOT_965( .ZN(g5770), .A(g992) );
  INV_X1 NOT_966( .ZN(II14219), .A(g801) );
  INV_X1 NOT_967( .ZN(g5771), .A(II14219) );
  INV_X1 NOT_968( .ZN(g5772), .A(g1193) );
  INV_X1 NOT_969( .ZN(g5773), .A(g1227) );
  INV_X1 NOT_970( .ZN(g5774), .A(g1439) );
  INV_X1 NOT_971( .ZN(g5775), .A(g1481) );
  INV_X1 NOT_972( .ZN(g5776), .A(g1597) );
  INV_X1 NOT_973( .ZN(g5777), .A(g1603) );
  INV_X1 NOT_974( .ZN(g5778), .A(g1680) );
  INV_X1 NOT_975( .ZN(g5785), .A(g1683) );
  INV_X1 NOT_976( .ZN(g5789), .A(g1886) );
  INV_X1 NOT_977( .ZN(g5790), .A(g2129) );
  INV_X1 NOT_978( .ZN(g5793), .A(g2170) );
  INV_X1 NOT_979( .ZN(g5794), .A(g2288) );
  INV_X1 NOT_980( .ZN(g5795), .A(g2376) );
  INV_X1 NOT_981( .ZN(II14238), .A(g2406) );
  INV_X1 NOT_982( .ZN(g5796), .A(II14238) );
  INV_X1 NOT_983( .ZN(II14243), .A(g3221) );
  INV_X1 NOT_984( .ZN(g5799), .A(II14243) );
  INV_X1 NOT_985( .ZN(II14246), .A(g3227) );
  INV_X1 NOT_986( .ZN(g5800), .A(II14246) );
  INV_X1 NOT_987( .ZN(II14249), .A(g3216) );
  INV_X1 NOT_988( .ZN(g5801), .A(II14249) );
  INV_X1 NOT_989( .ZN(g5802), .A(g83) );
  INV_X1 NOT_990( .ZN(g5803), .A(g117) );
  INV_X1 NOT_991( .ZN(g5804), .A(g237) );
  INV_X1 NOT_992( .ZN(g5805), .A(g243) );
  INV_X1 NOT_993( .ZN(g5806), .A(g249) );
  INV_X1 NOT_994( .ZN(g5808), .A(g509) );
  INV_X1 NOT_995( .ZN(g5809), .A(g780) );
  INV_X1 NOT_996( .ZN(g5810), .A(g740) );
  INV_X1 NOT_997( .ZN(g5811), .A(g801) );
  INV_X1 NOT_998( .ZN(g5812), .A(g915) );
  INV_X1 NOT_999( .ZN(g5813), .A(g921) );
  INV_X1 NOT_1000( .ZN(g5814), .A(g927) );
  INV_X1 NOT_1001( .ZN(g5815), .A(g991) );
  INV_X1 NOT_1002( .ZN(g5818), .A(g1194) );
  INV_X1 NOT_1003( .ZN(g5819), .A(g1430) );
  INV_X1 NOT_1004( .ZN(g5820), .A(g1486) );
  INV_X1 NOT_1005( .ZN(g5821), .A(g1600) );
  INV_X1 NOT_1006( .ZN(g5822), .A(g1606) );
  INV_X1 NOT_1007( .ZN(g5823), .A(g1612) );
  INV_X1 NOT_1008( .ZN(g5824), .A(g1486) );
  INV_X1 NOT_1009( .ZN(g5825), .A(g1684) );
  INV_X1 NOT_1010( .ZN(g5829), .A(g1686) );
  INV_X1 NOT_1011( .ZN(II14280), .A(g1491) );
  INV_X1 NOT_1012( .ZN(g5830), .A(II14280) );
  INV_X1 NOT_1013( .ZN(g5831), .A(g1887) );
  INV_X1 NOT_1014( .ZN(g5832), .A(g1921) );
  INV_X1 NOT_1015( .ZN(g5833), .A(g2133) );
  INV_X1 NOT_1016( .ZN(g5834), .A(g2175) );
  INV_X1 NOT_1017( .ZN(g5835), .A(g2291) );
  INV_X1 NOT_1018( .ZN(g5836), .A(g2297) );
  INV_X1 NOT_1019( .ZN(g5837), .A(g2374) );
  INV_X1 NOT_1020( .ZN(g5844), .A(g2377) );
  INV_X1 NOT_1021( .ZN(g5848), .A(g2580) );
  INV_X1 NOT_1022( .ZN(II14295), .A(g3228) );
  INV_X1 NOT_1023( .ZN(g5849), .A(II14295) );
  INV_X1 NOT_1024( .ZN(II14298), .A(g3217) );
  INV_X1 NOT_1025( .ZN(g5850), .A(II14298) );
  INV_X1 NOT_1026( .ZN(g5851), .A(g74) );
  INV_X1 NOT_1027( .ZN(g5852), .A(g121) );
  INV_X1 NOT_1028( .ZN(g5853), .A(g246) );
  INV_X1 NOT_1029( .ZN(g5854), .A(g252) );
  INV_X1 NOT_1030( .ZN(g5855), .A(g258) );
  INV_X1 NOT_1031( .ZN(II14306), .A(g97) );
  INV_X1 NOT_1032( .ZN(g5856), .A(II14306) );
  INV_X1 NOT_1033( .ZN(g5857), .A(g538) );
  INV_X1 NOT_1034( .ZN(g5858), .A(g771) );
  INV_X1 NOT_1035( .ZN(g5859), .A(g805) );
  INV_X1 NOT_1036( .ZN(g5860), .A(g924) );
  INV_X1 NOT_1037( .ZN(g5861), .A(g930) );
  INV_X1 NOT_1038( .ZN(g5862), .A(g936) );
  INV_X1 NOT_1039( .ZN(g5864), .A(g1195) );
  INV_X1 NOT_1040( .ZN(g5865), .A(g1466) );
  INV_X1 NOT_1041( .ZN(g5866), .A(g1426) );
  INV_X1 NOT_1042( .ZN(g5867), .A(g1491) );
  INV_X1 NOT_1043( .ZN(g5868), .A(g1609) );
  INV_X1 NOT_1044( .ZN(g5869), .A(g1615) );
  INV_X1 NOT_1045( .ZN(g5870), .A(g1621) );
  INV_X1 NOT_1046( .ZN(g5871), .A(g1685) );
  INV_X1 NOT_1047( .ZN(g5874), .A(g1888) );
  INV_X1 NOT_1048( .ZN(g5875), .A(g2124) );
  INV_X1 NOT_1049( .ZN(g5876), .A(g2180) );
  INV_X1 NOT_1050( .ZN(g5877), .A(g2294) );
  INV_X1 NOT_1051( .ZN(g5878), .A(g2300) );
  INV_X1 NOT_1052( .ZN(g5879), .A(g2306) );
  INV_X1 NOT_1053( .ZN(g5880), .A(g2180) );
  INV_X1 NOT_1054( .ZN(g5881), .A(g2378) );
  INV_X1 NOT_1055( .ZN(g5885), .A(g2380) );
  INV_X1 NOT_1056( .ZN(II14338), .A(g2185) );
  INV_X1 NOT_1057( .ZN(g5886), .A(II14338) );
  INV_X1 NOT_1058( .ZN(g5887), .A(g2581) );
  INV_X1 NOT_1059( .ZN(g5888), .A(g2615) );
  INV_X1 NOT_1060( .ZN(II14343), .A(g3219) );
  INV_X1 NOT_1061( .ZN(g5889), .A(II14343) );
  INV_X1 NOT_1062( .ZN(g5890), .A(g88) );
  INV_X1 NOT_1063( .ZN(g5893), .A(g125) );
  INV_X1 NOT_1064( .ZN(g5894), .A(g186) );
  INV_X1 NOT_1065( .ZN(g5895), .A(g255) );
  INV_X1 NOT_1066( .ZN(g5896), .A(g261) );
  INV_X1 NOT_1067( .ZN(g5897), .A(g267) );
  INV_X1 NOT_1068( .ZN(g5898), .A(g762) );
  INV_X1 NOT_1069( .ZN(g5899), .A(g809) );
  INV_X1 NOT_1070( .ZN(g5900), .A(g933) );
  INV_X1 NOT_1071( .ZN(g5901), .A(g939) );
  INV_X8 NOT_1072( .ZN(g5902), .A(g945) );
  INV_X8 NOT_1073( .ZN(II14357), .A(g785) );
  INV_X1 NOT_1074( .ZN(g5903), .A(II14357) );
  INV_X1 NOT_1075( .ZN(g5904), .A(g1224) );
  INV_X1 NOT_1076( .ZN(g5905), .A(g1457) );
  INV_X1 NOT_1077( .ZN(g5906), .A(g1496) );
  INV_X1 NOT_1078( .ZN(g5907), .A(g1618) );
  INV_X1 NOT_1079( .ZN(g5908), .A(g1624) );
  INV_X1 NOT_1080( .ZN(g5909), .A(g1630) );
  INV_X1 NOT_1081( .ZN(g5911), .A(g1889) );
  INV_X1 NOT_1082( .ZN(g5912), .A(g2160) );
  INV_X1 NOT_1083( .ZN(g5913), .A(g2120) );
  INV_X1 NOT_1084( .ZN(g5914), .A(g2185) );
  INV_X1 NOT_1085( .ZN(g5915), .A(g2303) );
  INV_X1 NOT_1086( .ZN(g5916), .A(g2309) );
  INV_X1 NOT_1087( .ZN(g5917), .A(g2315) );
  INV_X1 NOT_1088( .ZN(g5918), .A(g2379) );
  INV_X1 NOT_1089( .ZN(g5921), .A(g2582) );
  INV_X1 NOT_1090( .ZN(II14378), .A(g3234) );
  INV_X1 NOT_1091( .ZN(g5922), .A(II14378) );
  INV_X1 NOT_1092( .ZN(II14381), .A(g3223) );
  INV_X1 NOT_1093( .ZN(g5923), .A(II14381) );
  INV_X1 NOT_1094( .ZN(II14384), .A(g3218) );
  INV_X1 NOT_1095( .ZN(g5924), .A(II14384) );
  INV_X1 NOT_1096( .ZN(g5925), .A(g189) );
  INV_X1 NOT_1097( .ZN(g5926), .A(g195) );
  INV_X1 NOT_1098( .ZN(g5927), .A(g264) );
  INV_X1 NOT_1099( .ZN(g5928), .A(g270) );
  INV_X1 NOT_1100( .ZN(g5929), .A(g776) );
  INV_X1 NOT_1101( .ZN(g5932), .A(g813) );
  INV_X1 NOT_1102( .ZN(g5933), .A(g873) );
  INV_X1 NOT_1103( .ZN(g5934), .A(g942) );
  INV_X1 NOT_1104( .ZN(g5935), .A(g948) );
  INV_X1 NOT_1105( .ZN(g5936), .A(g954) );
  INV_X1 NOT_1106( .ZN(g5937), .A(g1448) );
  INV_X1 NOT_1107( .ZN(g5938), .A(g1501) );
  INV_X1 NOT_1108( .ZN(g5939), .A(g1627) );
  INV_X1 NOT_1109( .ZN(g5940), .A(g1633) );
  INV_X1 NOT_1110( .ZN(g5941), .A(g1639) );
  INV_X1 NOT_1111( .ZN(II14402), .A(g1471) );
  INV_X1 NOT_1112( .ZN(g5942), .A(II14402) );
  INV_X1 NOT_1113( .ZN(g5943), .A(g1918) );
  INV_X1 NOT_1114( .ZN(g5944), .A(g2151) );
  INV_X1 NOT_1115( .ZN(g5945), .A(g2190) );
  INV_X1 NOT_1116( .ZN(g5946), .A(g2312) );
  INV_X1 NOT_1117( .ZN(g5947), .A(g2318) );
  INV_X1 NOT_1118( .ZN(g5948), .A(g2324) );
  INV_X1 NOT_1119( .ZN(g5950), .A(g2583) );
  INV_X1 NOT_1120( .ZN(II14413), .A(g3233) );
  INV_X1 NOT_1121( .ZN(g5951), .A(II14413) );
  INV_X1 NOT_1122( .ZN(II14416), .A(g3222) );
  INV_X1 NOT_1123( .ZN(g5952), .A(II14416) );
  INV_X1 NOT_1124( .ZN(g5953), .A(g97) );
  INV_X1 NOT_1125( .ZN(g5954), .A(g192) );
  INV_X1 NOT_1126( .ZN(g5955), .A(g198) );
  INV_X1 NOT_1127( .ZN(g5956), .A(g204) );
  INV_X1 NOT_1128( .ZN(g5957), .A(g273) );
  INV_X1 NOT_1129( .ZN(II14424), .A(g117) );
  INV_X1 NOT_1130( .ZN(g5958), .A(II14424) );
  INV_X1 NOT_1131( .ZN(g5959), .A(g876) );
  INV_X1 NOT_1132( .ZN(g5960), .A(g882) );
  INV_X1 NOT_1133( .ZN(g5961), .A(g951) );
  INV_X1 NOT_1134( .ZN(g5962), .A(g957) );
  INV_X1 NOT_1135( .ZN(g5963), .A(g1462) );
  INV_X1 NOT_1136( .ZN(g5966), .A(g1506) );
  INV_X1 NOT_1137( .ZN(g5967), .A(g1567) );
  INV_X1 NOT_1138( .ZN(g5968), .A(g1636) );
  INV_X1 NOT_1139( .ZN(g5969), .A(g1642) );
  INV_X1 NOT_1140( .ZN(g5970), .A(g1648) );
  INV_X1 NOT_1141( .ZN(g5971), .A(g2142) );
  INV_X1 NOT_1142( .ZN(g5972), .A(g2195) );
  INV_X1 NOT_1143( .ZN(g5973), .A(g2321) );
  INV_X1 NOT_1144( .ZN(g5974), .A(g2327) );
  INV_X1 NOT_1145( .ZN(g5975), .A(g2333) );
  INV_X1 NOT_1146( .ZN(II14442), .A(g2165) );
  INV_X1 NOT_1147( .ZN(g5976), .A(II14442) );
  INV_X1 NOT_1148( .ZN(g5977), .A(g2612) );
  INV_X1 NOT_1149( .ZN(II14446), .A(g3230) );
  INV_X1 NOT_1150( .ZN(g5978), .A(II14446) );
  INV_X1 NOT_1151( .ZN(II14449), .A(g3224) );
  INV_X1 NOT_1152( .ZN(g5979), .A(II14449) );
  INV_X1 NOT_1153( .ZN(g5980), .A(g201) );
  INV_X1 NOT_1154( .ZN(g5981), .A(g207) );
  INV_X1 NOT_1155( .ZN(g5982), .A(g785) );
  INV_X1 NOT_1156( .ZN(g5983), .A(g879) );
  INV_X1 NOT_1157( .ZN(g5984), .A(g885) );
  INV_X1 NOT_1158( .ZN(g5985), .A(g891) );
  INV_X1 NOT_1159( .ZN(g5986), .A(g960) );
  INV_X1 NOT_1160( .ZN(II14459), .A(g805) );
  INV_X1 NOT_1161( .ZN(g5987), .A(II14459) );
  INV_X1 NOT_1162( .ZN(g5988), .A(g1570) );
  INV_X1 NOT_1163( .ZN(g5989), .A(g1576) );
  INV_X1 NOT_1164( .ZN(g5990), .A(g1645) );
  INV_X1 NOT_1165( .ZN(g5991), .A(g1651) );
  INV_X1 NOT_1166( .ZN(g5992), .A(g2156) );
  INV_X1 NOT_1167( .ZN(g5995), .A(g2200) );
  INV_X1 NOT_1168( .ZN(g5996), .A(g2261) );
  INV_X1 NOT_1169( .ZN(g5997), .A(g2330) );
  INV_X1 NOT_1170( .ZN(g5998), .A(g2336) );
  INV_X1 NOT_1171( .ZN(g5999), .A(g2342) );
  INV_X1 NOT_1172( .ZN(II14472), .A(g3080) );
  INV_X1 NOT_1173( .ZN(g6000), .A(II14472) );
  INV_X1 NOT_1174( .ZN(II14475), .A(g3225) );
  INV_X1 NOT_1175( .ZN(g6014), .A(II14475) );
  INV_X1 NOT_1176( .ZN(II14478), .A(g3213) );
  INV_X1 NOT_1177( .ZN(g6015), .A(II14478) );
  INV_X1 NOT_1178( .ZN(g6016), .A(g210) );
  INV_X1 NOT_1179( .ZN(g6017), .A(g888) );
  INV_X1 NOT_1180( .ZN(g6018), .A(g894) );
  INV_X1 NOT_1181( .ZN(g6019), .A(g1471) );
  INV_X1 NOT_1182( .ZN(g6020), .A(g1573) );
  INV_X8 NOT_1183( .ZN(g6021), .A(g1579) );
  INV_X8 NOT_1184( .ZN(g6022), .A(g1585) );
  INV_X8 NOT_1185( .ZN(g6023), .A(g1654) );
  INV_X1 NOT_1186( .ZN(II14489), .A(g1496) );
  INV_X1 NOT_1187( .ZN(g6024), .A(II14489) );
  INV_X1 NOT_1188( .ZN(g6025), .A(g2264) );
  INV_X1 NOT_1189( .ZN(g6026), .A(g2270) );
  INV_X1 NOT_1190( .ZN(g6027), .A(g2339) );
  INV_X1 NOT_1191( .ZN(g6028), .A(g2345) );
  INV_X1 NOT_1192( .ZN(II14496), .A(g3226) );
  INV_X1 NOT_1193( .ZN(g6029), .A(II14496) );
  INV_X1 NOT_1194( .ZN(II14499), .A(g3214) );
  INV_X1 NOT_1195( .ZN(g6030), .A(II14499) );
  INV_X1 NOT_1196( .ZN(II14502), .A(g471) );
  INV_X1 NOT_1197( .ZN(g6031), .A(II14502) );
  INV_X1 NOT_1198( .ZN(g6032), .A(g897) );
  INV_X1 NOT_1199( .ZN(g6033), .A(g1582) );
  INV_X1 NOT_1200( .ZN(g6034), .A(g1588) );
  INV_X1 NOT_1201( .ZN(g6035), .A(g2165) );
  INV_X1 NOT_1202( .ZN(g6036), .A(g2267) );
  INV_X1 NOT_1203( .ZN(g6037), .A(g2273) );
  INV_X1 NOT_1204( .ZN(g6038), .A(g2279) );
  INV_X1 NOT_1205( .ZN(g6039), .A(g2348) );
  INV_X1 NOT_1206( .ZN(II14513), .A(g2190) );
  INV_X1 NOT_1207( .ZN(g6040), .A(II14513) );
  INV_X1 NOT_1208( .ZN(II14516), .A(g3215) );
  INV_X1 NOT_1209( .ZN(g6041), .A(II14516) );
  INV_X1 NOT_1210( .ZN(II14519), .A(g1158) );
  INV_X1 NOT_1211( .ZN(g6042), .A(II14519) );
  INV_X1 NOT_1212( .ZN(g6043), .A(g1591) );
  INV_X1 NOT_1213( .ZN(g6044), .A(g2276) );
  INV_X1 NOT_1214( .ZN(g6045), .A(g2282) );
  INV_X1 NOT_1215( .ZN(II14525), .A(g1852) );
  INV_X1 NOT_1216( .ZN(g6046), .A(II14525) );
  INV_X1 NOT_1217( .ZN(g6047), .A(g2285) );
  INV_X1 NOT_1218( .ZN(II14529), .A(g3142) );
  INV_X1 NOT_1219( .ZN(g6048), .A(II14529) );
  INV_X1 NOT_1220( .ZN(II14532), .A(g354) );
  INV_X1 NOT_1221( .ZN(g6051), .A(II14532) );
  INV_X1 NOT_1222( .ZN(II14535), .A(g2546) );
  INV_X1 NOT_1223( .ZN(g6052), .A(II14535) );
  INV_X1 NOT_1224( .ZN(II14538), .A(g369) );
  INV_X1 NOT_1225( .ZN(g6053), .A(II14538) );
  INV_X1 NOT_1226( .ZN(II14541), .A(g455) );
  INV_X1 NOT_1227( .ZN(g6054), .A(II14541) );
  INV_X1 NOT_1228( .ZN(II14544), .A(g1041) );
  INV_X1 NOT_1229( .ZN(g6055), .A(II14544) );
  INV_X1 NOT_1230( .ZN(II14547), .A(g384) );
  INV_X1 NOT_1231( .ZN(g6056), .A(II14547) );
  INV_X1 NOT_1232( .ZN(II14550), .A(g458) );
  INV_X1 NOT_1233( .ZN(g6057), .A(II14550) );
  INV_X1 NOT_1234( .ZN(II14553), .A(g1056) );
  INV_X1 NOT_1235( .ZN(g6058), .A(II14553) );
  INV_X1 NOT_1236( .ZN(II14556), .A(g1142) );
  INV_X1 NOT_1237( .ZN(g6059), .A(II14556) );
  INV_X1 NOT_1238( .ZN(II14559), .A(g1735) );
  INV_X1 NOT_1239( .ZN(g6060), .A(II14559) );
  INV_X1 NOT_1240( .ZN(II14562), .A(g398) );
  INV_X1 NOT_1241( .ZN(g6061), .A(II14562) );
  INV_X1 NOT_1242( .ZN(II14565), .A(g461) );
  INV_X1 NOT_1243( .ZN(g6062), .A(II14565) );
  INV_X1 NOT_1244( .ZN(II14568), .A(g1071) );
  INV_X1 NOT_1245( .ZN(g6063), .A(II14568) );
  INV_X1 NOT_1246( .ZN(II14571), .A(g1145) );
  INV_X1 NOT_1247( .ZN(g6064), .A(II14571) );
  INV_X1 NOT_1248( .ZN(II14574), .A(g1750) );
  INV_X1 NOT_1249( .ZN(g6065), .A(II14574) );
  INV_X1 NOT_1250( .ZN(II14577), .A(g1836) );
  INV_X1 NOT_1251( .ZN(g6066), .A(II14577) );
  INV_X1 NOT_1252( .ZN(II14580), .A(g2429) );
  INV_X1 NOT_1253( .ZN(g6067), .A(II14580) );
  INV_X1 NOT_1254( .ZN(g6068), .A(g499) );
  INV_X1 NOT_1255( .ZN(II14584), .A(g465) );
  INV_X1 NOT_1256( .ZN(g6079), .A(II14584) );
  INV_X1 NOT_1257( .ZN(II14587), .A(g1085) );
  INV_X1 NOT_1258( .ZN(g6080), .A(II14587) );
  INV_X1 NOT_1259( .ZN(II14590), .A(g1148) );
  INV_X1 NOT_1260( .ZN(g6081), .A(II14590) );
  INV_X1 NOT_1261( .ZN(II14593), .A(g1765) );
  INV_X1 NOT_1262( .ZN(g6082), .A(II14593) );
  INV_X1 NOT_1263( .ZN(II14596), .A(g1839) );
  INV_X1 NOT_1264( .ZN(g6083), .A(II14596) );
  INV_X1 NOT_1265( .ZN(II14599), .A(g2444) );
  INV_X1 NOT_1266( .ZN(g6084), .A(II14599) );
  INV_X1 NOT_1267( .ZN(II14602), .A(g2530) );
  INV_X1 NOT_1268( .ZN(g6085), .A(II14602) );
  INV_X1 NOT_1269( .ZN(II14605), .A(g468) );
  INV_X1 NOT_1270( .ZN(g6086), .A(II14605) );
  INV_X1 NOT_1271( .ZN(g6087), .A(g1186) );
  INV_X1 NOT_1272( .ZN(II14609), .A(g1152) );
  INV_X1 NOT_1273( .ZN(g6098), .A(II14609) );
  INV_X1 NOT_1274( .ZN(II14612), .A(g1779) );
  INV_X1 NOT_1275( .ZN(g6099), .A(II14612) );
  INV_X1 NOT_1276( .ZN(II14615), .A(g1842) );
  INV_X1 NOT_1277( .ZN(g6100), .A(II14615) );
  INV_X1 NOT_1278( .ZN(II14618), .A(g2459) );
  INV_X1 NOT_1279( .ZN(g6101), .A(II14618) );
  INV_X1 NOT_1280( .ZN(II14621), .A(g2533) );
  INV_X1 NOT_1281( .ZN(g6102), .A(II14621) );
  INV_X1 NOT_1282( .ZN(II14624), .A(g1155) );
  INV_X1 NOT_1283( .ZN(g6103), .A(II14624) );
  INV_X1 NOT_1284( .ZN(g6104), .A(g1880) );
  INV_X8 NOT_1285( .ZN(II14628), .A(g1846) );
  INV_X8 NOT_1286( .ZN(g6115), .A(II14628) );
  INV_X8 NOT_1287( .ZN(II14631), .A(g2473) );
  INV_X8 NOT_1288( .ZN(g6116), .A(II14631) );
  INV_X8 NOT_1289( .ZN(II14634), .A(g2536) );
  INV_X1 NOT_1290( .ZN(g6117), .A(II14634) );
  INV_X1 NOT_1291( .ZN(II14637), .A(g1849) );
  INV_X1 NOT_1292( .ZN(g6118), .A(II14637) );
  INV_X1 NOT_1293( .ZN(g6119), .A(g2574) );
  INV_X1 NOT_1294( .ZN(II14641), .A(g2540) );
  INV_X1 NOT_1295( .ZN(g6130), .A(II14641) );
  INV_X1 NOT_1296( .ZN(II14644), .A(g3142) );
  INV_X1 NOT_1297( .ZN(g6131), .A(II14644) );
  INV_X1 NOT_1298( .ZN(II14647), .A(g2543) );
  INV_X1 NOT_1299( .ZN(g6134), .A(II14647) );
  INV_X1 NOT_1300( .ZN(II14650), .A(g525) );
  INV_X1 NOT_1301( .ZN(g6135), .A(II14650) );
  INV_X1 NOT_1302( .ZN(g6136), .A(g672) );
  INV_X1 NOT_1303( .ZN(II14654), .A(g3220) );
  INV_X1 NOT_1304( .ZN(g6139), .A(II14654) );
  INV_X1 NOT_1305( .ZN(g6140), .A(g524) );
  INV_X1 NOT_1306( .ZN(g6141), .A(g554) );
  INV_X1 NOT_1307( .ZN(g6142), .A(g679) );
  INV_X1 NOT_1308( .ZN(II14660), .A(g1211) );
  INV_X1 NOT_1309( .ZN(g6145), .A(II14660) );
  INV_X1 NOT_1310( .ZN(g6146), .A(g1358) );
  INV_X1 NOT_1311( .ZN(g6149), .A(g3097) );
  INV_X1 NOT_1312( .ZN(II14665), .A(g3147) );
  INV_X1 NOT_1313( .ZN(g6153), .A(II14665) );
  INV_X1 NOT_1314( .ZN(II14668), .A(g3232) );
  INV_X1 NOT_1315( .ZN(g6156), .A(II14668) );
  INV_X1 NOT_1316( .ZN(g6157), .A(g686) );
  INV_X1 NOT_1317( .ZN(g6161), .A(g1210) );
  INV_X1 NOT_1318( .ZN(g6162), .A(g1240) );
  INV_X1 NOT_1319( .ZN(g6163), .A(g1365) );
  INV_X1 NOT_1320( .ZN(II14675), .A(g1905) );
  INV_X1 NOT_1321( .ZN(g6166), .A(II14675) );
  INV_X1 NOT_1322( .ZN(g6167), .A(g2052) );
  INV_X1 NOT_1323( .ZN(g6170), .A(g3098) );
  INV_X1 NOT_1324( .ZN(g6173), .A(g557) );
  INV_X1 NOT_1325( .ZN(g6177), .A(g633) );
  INV_X1 NOT_1326( .ZN(g6180), .A(g692) );
  INV_X1 NOT_1327( .ZN(g6183), .A(g291) );
  INV_X1 NOT_1328( .ZN(g6184), .A(g1372) );
  INV_X1 NOT_1329( .ZN(g6188), .A(g1904) );
  INV_X1 NOT_1330( .ZN(g6189), .A(g1934) );
  INV_X1 NOT_1331( .ZN(g6190), .A(g2059) );
  INV_X1 NOT_1332( .ZN(II14688), .A(g2599) );
  INV_X1 NOT_1333( .ZN(g6193), .A(II14688) );
  INV_X1 NOT_1334( .ZN(g6194), .A(g2746) );
  INV_X1 NOT_1335( .ZN(g6197), .A(g3099) );
  INV_X1 NOT_1336( .ZN(g6200), .A(g542) );
  INV_X1 NOT_1337( .ZN(g6201), .A(g646) );
  INV_X1 NOT_1338( .ZN(g6204), .A(g289) );
  INV_X1 NOT_1339( .ZN(g6205), .A(g1243) );
  INV_X1 NOT_1340( .ZN(g6209), .A(g1319) );
  INV_X1 NOT_1341( .ZN(g6212), .A(g1378) );
  INV_X1 NOT_1342( .ZN(g6215), .A(g978) );
  INV_X1 NOT_1343( .ZN(g6216), .A(g2066) );
  INV_X1 NOT_1344( .ZN(g6220), .A(g2598) );
  INV_X1 NOT_1345( .ZN(g6221), .A(g2628) );
  INV_X1 NOT_1346( .ZN(g6222), .A(g2753) );
  INV_X1 NOT_1347( .ZN(II14704), .A(g2818) );
  INV_X1 NOT_1348( .ZN(g6225), .A(II14704) );
  INV_X1 NOT_1349( .ZN(g6226), .A(g2818) );
  INV_X1 NOT_1350( .ZN(g6227), .A(g3100) );
  INV_X1 NOT_1351( .ZN(II14709), .A(g3229) );
  INV_X1 NOT_1352( .ZN(g6230), .A(II14709) );
  INV_X1 NOT_1353( .ZN(II14712), .A(g138) );
  INV_X1 NOT_1354( .ZN(g6231), .A(II14712) );
  INV_X1 NOT_1355( .ZN(II14715), .A(g138) );
  INV_X1 NOT_1356( .ZN(g6232), .A(II14715) );
  INV_X1 NOT_1357( .ZN(g6281), .A(g510) );
  INV_X1 NOT_1358( .ZN(g6284), .A(g640) );
  INV_X1 NOT_1359( .ZN(g6288), .A(g287) );
  INV_X1 NOT_1360( .ZN(g6289), .A(g1228) );
  INV_X1 NOT_1361( .ZN(g6290), .A(g1332) );
  INV_X1 NOT_1362( .ZN(g6293), .A(g976) );
  INV_X1 NOT_1363( .ZN(g6294), .A(g1937) );
  INV_X1 NOT_1364( .ZN(g6298), .A(g2013) );
  INV_X1 NOT_1365( .ZN(g6301), .A(g2072) );
  INV_X1 NOT_1366( .ZN(g6304), .A(g1672) );
  INV_X1 NOT_1367( .ZN(g6305), .A(g2760) );
  INV_X1 NOT_1368( .ZN(g6309), .A(g14) );
  INV_X1 NOT_1369( .ZN(g6310), .A(g3101) );
  INV_X1 NOT_1370( .ZN(II14731), .A(g135) );
  INV_X1 NOT_1371( .ZN(g6313), .A(II14731) );
  INV_X1 NOT_1372( .ZN(II14734), .A(g135) );
  INV_X1 NOT_1373( .ZN(g6314), .A(II14734) );
  INV_X1 NOT_1374( .ZN(g6363), .A(g653) );
  INV_X1 NOT_1375( .ZN(g6367), .A(g285) );
  INV_X1 NOT_1376( .ZN(II14739), .A(g826) );
  INV_X1 NOT_1377( .ZN(g6368), .A(II14739) );
  INV_X1 NOT_1378( .ZN(II14742), .A(g826) );
  INV_X1 NOT_1379( .ZN(g6369), .A(II14742) );
  INV_X1 NOT_1380( .ZN(g6418), .A(g1196) );
  INV_X1 NOT_1381( .ZN(g6421), .A(g1326) );
  INV_X1 NOT_1382( .ZN(g6425), .A(g974) );
  INV_X1 NOT_1383( .ZN(g6426), .A(g1922) );
  INV_X1 NOT_1384( .ZN(g6427), .A(g2026) );
  INV_X1 NOT_1385( .ZN(g6430), .A(g1670) );
  INV_X1 NOT_1386( .ZN(g6431), .A(g2631) );
  INV_X1 NOT_1387( .ZN(g6435), .A(g2707) );
  INV_X1 NOT_1388( .ZN(g6438), .A(g2766) );
  INV_X1 NOT_1389( .ZN(g6441), .A(g2366) );
  INV_X1 NOT_1390( .ZN(II14755), .A(g2821) );
  INV_X1 NOT_1391( .ZN(g6442), .A(II14755) );
  INV_X1 NOT_1392( .ZN(g6443), .A(g2821) );
  INV_X1 NOT_1393( .ZN(g6444), .A(g3102) );
  INV_X1 NOT_1394( .ZN(II14760), .A(g405) );
  INV_X1 NOT_1395( .ZN(g6447), .A(II14760) );
  INV_X1 NOT_1396( .ZN(II14763), .A(g405) );
  INV_X1 NOT_1397( .ZN(g6448), .A(II14763) );
  INV_X1 NOT_1398( .ZN(II14766), .A(g545) );
  INV_X1 NOT_1399( .ZN(g6485), .A(II14766) );
  INV_X1 NOT_1400( .ZN(II14769), .A(g545) );
  INV_X1 NOT_1401( .ZN(g6486), .A(II14769) );
  INV_X1 NOT_1402( .ZN(g6512), .A(g544) );
  INV_X1 NOT_1403( .ZN(g6513), .A(g660) );
  INV_X1 NOT_1404( .ZN(g6517), .A(g283) );
  INV_X1 NOT_1405( .ZN(II14775), .A(g823) );
  INV_X1 NOT_1406( .ZN(g6518), .A(II14775) );
  INV_X1 NOT_1407( .ZN(II14778), .A(g823) );
  INV_X1 NOT_1408( .ZN(g6519), .A(II14778) );
  INV_X1 NOT_1409( .ZN(g6568), .A(g1339) );
  INV_X8 NOT_1410( .ZN(g6572), .A(g972) );
  INV_X8 NOT_1411( .ZN(II14783), .A(g1520) );
  INV_X8 NOT_1412( .ZN(g6573), .A(II14783) );
  INV_X1 NOT_1413( .ZN(II14786), .A(g1520) );
  INV_X1 NOT_1414( .ZN(g6574), .A(II14786) );
  INV_X1 NOT_1415( .ZN(g6623), .A(g1890) );
  INV_X1 NOT_1416( .ZN(g6626), .A(g2020) );
  INV_X1 NOT_1417( .ZN(g6630), .A(g1668) );
  INV_X1 NOT_1418( .ZN(g6631), .A(g2616) );
  INV_X1 NOT_1419( .ZN(g6632), .A(g2720) );
  INV_X1 NOT_1420( .ZN(g6635), .A(g2364) );
  INV_X1 NOT_1421( .ZN(g6636), .A(g1491) );
  INV_X1 NOT_1422( .ZN(g6637), .A(g5) );
  INV_X1 NOT_1423( .ZN(g6638), .A(g3103) );
  INV_X1 NOT_1424( .ZN(g6641), .A(g113) );
  INV_X1 NOT_1425( .ZN(II14799), .A(g551) );
  INV_X1 NOT_1426( .ZN(g6642), .A(II14799) );
  INV_X1 NOT_1427( .ZN(II14802), .A(g551) );
  INV_X1 NOT_1428( .ZN(g6643), .A(II14802) );
  INV_X1 NOT_1429( .ZN(g6672), .A(g464) );
  INV_X1 NOT_1430( .ZN(g6675), .A(g458) );
  INV_X1 NOT_1431( .ZN(g6676), .A(g559) );
  INV_X1 NOT_1432( .ZN(II14808), .A(g623) );
  INV_X1 NOT_1433( .ZN(g6677), .A(II14808) );
  INV_X1 NOT_1434( .ZN(II14811), .A(g623) );
  INV_X1 NOT_1435( .ZN(g6678), .A(II14811) );
  INV_X1 NOT_1436( .ZN(g6707), .A(g666) );
  INV_X1 NOT_1437( .ZN(g6711), .A(g281) );
  INV_X1 NOT_1438( .ZN(II14816), .A(g1092) );
  INV_X1 NOT_1439( .ZN(g6712), .A(II14816) );
  INV_X1 NOT_1440( .ZN(II14819), .A(g1092) );
  INV_X1 NOT_1441( .ZN(g6713), .A(II14819) );
  INV_X1 NOT_1442( .ZN(II14822), .A(g1231) );
  INV_X1 NOT_1443( .ZN(g6750), .A(II14822) );
  INV_X1 NOT_1444( .ZN(II14825), .A(g1231) );
  INV_X1 NOT_1445( .ZN(g6751), .A(II14825) );
  INV_X1 NOT_1446( .ZN(g6776), .A(g1230) );
  INV_X1 NOT_1447( .ZN(g6777), .A(g1346) );
  INV_X1 NOT_1448( .ZN(g6781), .A(g970) );
  INV_X1 NOT_1449( .ZN(II14831), .A(g1517) );
  INV_X1 NOT_1450( .ZN(g6782), .A(II14831) );
  INV_X1 NOT_1451( .ZN(II14834), .A(g1517) );
  INV_X1 NOT_1452( .ZN(g6783), .A(II14834) );
  INV_X1 NOT_1453( .ZN(g6832), .A(g2033) );
  INV_X1 NOT_1454( .ZN(g6836), .A(g1666) );
  INV_X1 NOT_1455( .ZN(II14839), .A(g2214) );
  INV_X1 NOT_1456( .ZN(g6837), .A(II14839) );
  INV_X1 NOT_1457( .ZN(II14842), .A(g2214) );
  INV_X1 NOT_1458( .ZN(g6838), .A(II14842) );
  INV_X1 NOT_1459( .ZN(g6887), .A(g2584) );
  INV_X1 NOT_1460( .ZN(g6890), .A(g2714) );
  INV_X1 NOT_1461( .ZN(g6894), .A(g2362) );
  INV_X1 NOT_1462( .ZN(II14848), .A(g2824) );
  INV_X1 NOT_1463( .ZN(g6895), .A(II14848) );
  INV_X1 NOT_1464( .ZN(g6896), .A(g2824) );
  INV_X1 NOT_1465( .ZN(g6897), .A(g1486) );
  INV_X1 NOT_1466( .ZN(g6898), .A(g2993) );
  INV_X1 NOT_1467( .ZN(g6901), .A(g3006) );
  INV_X1 NOT_1468( .ZN(g6905), .A(g3104) );
  INV_X1 NOT_1469( .ZN(g6908), .A(g484) );
  INV_X1 NOT_1470( .ZN(II14857), .A(g626) );
  INV_X1 NOT_1471( .ZN(g6911), .A(II14857) );
  INV_X1 NOT_1472( .ZN(II14860), .A(g626) );
  INV_X1 NOT_1473( .ZN(g6912), .A(II14860) );
  INV_X1 NOT_1474( .ZN(g6942), .A(g279) );
  INV_X1 NOT_1475( .ZN(g6943), .A(g801) );
  INV_X1 NOT_1476( .ZN(II14865), .A(g1237) );
  INV_X1 NOT_1477( .ZN(g6944), .A(II14865) );
  INV_X1 NOT_1478( .ZN(II14868), .A(g1237) );
  INV_X1 NOT_1479( .ZN(g6945), .A(II14868) );
  INV_X1 NOT_1480( .ZN(g6974), .A(g1151) );
  INV_X1 NOT_1481( .ZN(g6977), .A(g1145) );
  INV_X1 NOT_1482( .ZN(g6978), .A(g1245) );
  INV_X1 NOT_1483( .ZN(II14874), .A(g1309) );
  INV_X1 NOT_1484( .ZN(g6979), .A(II14874) );
  INV_X1 NOT_1485( .ZN(II14877), .A(g1309) );
  INV_X1 NOT_1486( .ZN(g6980), .A(II14877) );
  INV_X1 NOT_1487( .ZN(g7009), .A(g1352) );
  INV_X1 NOT_1488( .ZN(g7013), .A(g968) );
  INV_X1 NOT_1489( .ZN(II14882), .A(g1786) );
  INV_X1 NOT_1490( .ZN(g7014), .A(II14882) );
  INV_X1 NOT_1491( .ZN(II14885), .A(g1786) );
  INV_X1 NOT_1492( .ZN(g7015), .A(II14885) );
  INV_X1 NOT_1493( .ZN(II14888), .A(g1925) );
  INV_X1 NOT_1494( .ZN(g7052), .A(II14888) );
  INV_X1 NOT_1495( .ZN(II14891), .A(g1925) );
  INV_X1 NOT_1496( .ZN(g7053), .A(II14891) );
  INV_X1 NOT_1497( .ZN(g7078), .A(g1924) );
  INV_X1 NOT_1498( .ZN(g7079), .A(g2040) );
  INV_X1 NOT_1499( .ZN(g7083), .A(g1664) );
  INV_X1 NOT_1500( .ZN(II14897), .A(g2211) );
  INV_X1 NOT_1501( .ZN(g7084), .A(II14897) );
  INV_X1 NOT_1502( .ZN(II14900), .A(g2211) );
  INV_X1 NOT_1503( .ZN(g7085), .A(II14900) );
  INV_X1 NOT_1504( .ZN(g7134), .A(g2727) );
  INV_X1 NOT_1505( .ZN(g7138), .A(g2360) );
  INV_X1 NOT_1506( .ZN(g7139), .A(g1481) );
  INV_X1 NOT_1507( .ZN(g7140), .A(g2170) );
  INV_X1 NOT_1508( .ZN(g7141), .A(g2195) );
  INV_X1 NOT_1509( .ZN(g7142), .A(g8) );
  INV_X1 NOT_1510( .ZN(g7143), .A(g2998) );
  INV_X1 NOT_1511( .ZN(g7146), .A(g3013) );
  INV_X1 NOT_1512( .ZN(g7149), .A(g3105) );
  INV_X1 NOT_1513( .ZN(g7152), .A(g3136) );
  INV_X1 NOT_1514( .ZN(g7153), .A(g480) );
  INV_X1 NOT_1515( .ZN(g7156), .A(g461) );
  INV_X1 NOT_1516( .ZN(g7157), .A(g453) );
  INV_X1 NOT_1517( .ZN(g7158), .A(g1171) );
  INV_X1 NOT_1518( .ZN(II14917), .A(g1312) );
  INV_X1 NOT_1519( .ZN(g7161), .A(II14917) );
  INV_X1 NOT_1520( .ZN(II14920), .A(g1312) );
  INV_X1 NOT_1521( .ZN(g7162), .A(II14920) );
  INV_X4 NOT_1522( .ZN(g7192), .A(g966) );
  INV_X4 NOT_1523( .ZN(g7193), .A(g1491) );
  INV_X1 NOT_1524( .ZN(II14925), .A(g1931) );
  INV_X1 NOT_1525( .ZN(g7194), .A(II14925) );
  INV_X1 NOT_1526( .ZN(II14928), .A(g1931) );
  INV_X1 NOT_1527( .ZN(g7195), .A(II14928) );
  INV_X1 NOT_1528( .ZN(g7224), .A(g1845) );
  INV_X1 NOT_1529( .ZN(g7227), .A(g1839) );
  INV_X1 NOT_1530( .ZN(g7228), .A(g1939) );
  INV_X1 NOT_1531( .ZN(II14934), .A(g2003) );
  INV_X1 NOT_1532( .ZN(g7229), .A(II14934) );
  INV_X1 NOT_1533( .ZN(II14937), .A(g2003) );
  INV_X1 NOT_1534( .ZN(g7230), .A(II14937) );
  INV_X1 NOT_1535( .ZN(g7259), .A(g2046) );
  INV_X1 NOT_1536( .ZN(g7263), .A(g1662) );
  INV_X1 NOT_1537( .ZN(II14942), .A(g2480) );
  INV_X1 NOT_1538( .ZN(g7264), .A(II14942) );
  INV_X1 NOT_1539( .ZN(II14945), .A(g2480) );
  INV_X1 NOT_1540( .ZN(g7265), .A(II14945) );
  INV_X1 NOT_1541( .ZN(II14948), .A(g2619) );
  INV_X1 NOT_1542( .ZN(g7302), .A(II14948) );
  INV_X1 NOT_1543( .ZN(II14951), .A(g2619) );
  INV_X1 NOT_1544( .ZN(g7303), .A(II14951) );
  INV_X1 NOT_1545( .ZN(g7328), .A(g2618) );
  INV_X1 NOT_1546( .ZN(g7329), .A(g2734) );
  INV_X1 NOT_1547( .ZN(g7333), .A(g2358) );
  INV_X1 NOT_1548( .ZN(II14957), .A(g2827) );
  INV_X1 NOT_1549( .ZN(g7334), .A(II14957) );
  INV_X1 NOT_1550( .ZN(g7335), .A(g2827) );
  INV_X1 NOT_1551( .ZN(g7336), .A(g1476) );
  INV_X1 NOT_1552( .ZN(g7337), .A(g2190) );
  INV_X1 NOT_1553( .ZN(g7338), .A(g3002) );
  INV_X1 NOT_1554( .ZN(g7342), .A(g3024) );
  INV_X1 NOT_1555( .ZN(g7345), .A(g3139) );
  INV_X1 NOT_1556( .ZN(g7346), .A(g97) );
  INV_X1 NOT_1557( .ZN(g7347), .A(g490) );
  INV_X1 NOT_1558( .ZN(g7348), .A(g451) );
  INV_X1 NOT_1559( .ZN(g7349), .A(g1167) );
  INV_X1 NOT_1560( .ZN(g7352), .A(g1148) );
  INV_X1 NOT_1561( .ZN(g7353), .A(g1140) );
  INV_X1 NOT_1562( .ZN(g7354), .A(g1865) );
  INV_X1 NOT_1563( .ZN(II14973), .A(g2006) );
  INV_X1 NOT_1564( .ZN(g7357), .A(II14973) );
  INV_X1 NOT_1565( .ZN(II14976), .A(g2006) );
  INV_X1 NOT_1566( .ZN(g7358), .A(II14976) );
  INV_X1 NOT_1567( .ZN(g7388), .A(g1660) );
  INV_X1 NOT_1568( .ZN(g7389), .A(g2185) );
  INV_X1 NOT_1569( .ZN(II14981), .A(g2625) );
  INV_X1 NOT_1570( .ZN(g7390), .A(II14981) );
  INV_X1 NOT_1571( .ZN(II14984), .A(g2625) );
  INV_X1 NOT_1572( .ZN(g7391), .A(II14984) );
  INV_X1 NOT_1573( .ZN(g7420), .A(g2539) );
  INV_X1 NOT_1574( .ZN(g7423), .A(g2533) );
  INV_X1 NOT_1575( .ZN(g7424), .A(g2633) );
  INV_X1 NOT_1576( .ZN(II14990), .A(g2697) );
  INV_X1 NOT_1577( .ZN(g7425), .A(II14990) );
  INV_X1 NOT_1578( .ZN(II14993), .A(g2697) );
  INV_X1 NOT_1579( .ZN(g7426), .A(II14993) );
  INV_X1 NOT_1580( .ZN(g7455), .A(g2740) );
  INV_X1 NOT_1581( .ZN(g7459), .A(g2356) );
  INV_X1 NOT_1582( .ZN(g7460), .A(g1471) );
  INV_X1 NOT_1583( .ZN(g7461), .A(g2175) );
  INV_X1 NOT_1584( .ZN(g7462), .A(g2912) );
  INV_X1 NOT_1585( .ZN(g7465), .A(g2) );
  INV_X1 NOT_1586( .ZN(g7466), .A(g3010) );
  INV_X1 NOT_1587( .ZN(g7471), .A(g3036) );
  INV_X1 NOT_1588( .ZN(g7475), .A(g493) );
  INV_X1 NOT_1589( .ZN(g7476), .A(g785) );
  INV_X4 NOT_1590( .ZN(g7477), .A(g1177) );
  INV_X4 NOT_1591( .ZN(g7478), .A(g1138) );
  INV_X1 NOT_1592( .ZN(g7479), .A(g1861) );
  INV_X1 NOT_1593( .ZN(g7482), .A(g1842) );
  INV_X1 NOT_1594( .ZN(g7483), .A(g1834) );
  INV_X1 NOT_1595( .ZN(g7484), .A(g2559) );
  INV_X1 NOT_1596( .ZN(II15012), .A(g2700) );
  INV_X1 NOT_1597( .ZN(g7487), .A(II15012) );
  INV_X1 NOT_1598( .ZN(II15015), .A(g2700) );
  INV_X1 NOT_1599( .ZN(g7488), .A(II15015) );
  INV_X1 NOT_1600( .ZN(g7518), .A(g2354) );
  INV_X1 NOT_1601( .ZN(II15019), .A(g2830) );
  INV_X1 NOT_1602( .ZN(g7519), .A(II15019) );
  INV_X1 NOT_1603( .ZN(g7520), .A(g2830) );
  INV_X1 NOT_1604( .ZN(g7521), .A(g2200) );
  INV_X1 NOT_1605( .ZN(g7522), .A(g2917) );
  INV_X1 NOT_1606( .ZN(g7527), .A(g3018) );
  INV_X1 NOT_1607( .ZN(g7529), .A(g465) );
  INV_X1 NOT_1608( .ZN(g7530), .A(g496) );
  INV_X1 NOT_1609( .ZN(g7531), .A(g1180) );
  INV_X1 NOT_1610( .ZN(g7532), .A(g1471) );
  INV_X1 NOT_1611( .ZN(g7533), .A(g1871) );
  INV_X1 NOT_1612( .ZN(g7534), .A(g1832) );
  INV_X1 NOT_1613( .ZN(g7535), .A(g2555) );
  INV_X1 NOT_1614( .ZN(g7538), .A(g2536) );
  INV_X1 NOT_1615( .ZN(g7539), .A(g2528) );
  INV_X1 NOT_1616( .ZN(g7540), .A(g1506) );
  INV_X1 NOT_1617( .ZN(g7541), .A(g2180) );
  INV_X1 NOT_1618( .ZN(g7542), .A(g2883) );
  INV_X1 NOT_1619( .ZN(g7545), .A(g2920) );
  INV_X1 NOT_1620( .ZN(g7548), .A(g2990) );
  INV_X1 NOT_1621( .ZN(g7549), .A(g3028) );
  INV_X1 NOT_1622( .ZN(g7553), .A(g3114) );
  INV_X1 NOT_1623( .ZN(g7554), .A(g117) );
  INV_X1 NOT_1624( .ZN(g7555), .A(g1152) );
  INV_X1 NOT_1625( .ZN(g7556), .A(g1183) );
  INV_X1 NOT_1626( .ZN(g7557), .A(g1874) );
  INV_X1 NOT_1627( .ZN(g7558), .A(g2165) );
  INV_X1 NOT_1628( .ZN(g7559), .A(g2565) );
  INV_X1 NOT_1629( .ZN(g7560), .A(g2526) );
  INV_X1 NOT_1630( .ZN(g7561), .A(g1501) );
  INV_X1 NOT_1631( .ZN(g7562), .A(g2888) );
  INV_X1 NOT_1632( .ZN(g7566), .A(g2896) );
  INV_X1 NOT_1633( .ZN(g7570), .A(g3032) );
  INV_X1 NOT_1634( .ZN(g7573), .A(g3120) );
  INV_X1 NOT_1635( .ZN(g7574), .A(g3128) );
  INV_X1 NOT_1636( .ZN(g7576), .A(g468) );
  INV_X1 NOT_1637( .ZN(g7577), .A(g805) );
  INV_X1 NOT_1638( .ZN(g7578), .A(g1846) );
  INV_X1 NOT_1639( .ZN(g7579), .A(g1877) );
  INV_X1 NOT_1640( .ZN(g7580), .A(g2568) );
  INV_X1 NOT_1641( .ZN(g7581), .A(g1496) );
  INV_X1 NOT_1642( .ZN(g7582), .A(g2185) );
  INV_X1 NOT_1643( .ZN(g7583), .A(g2892) );
  INV_X1 NOT_1644( .ZN(g7587), .A(g2903) );
  INV_X1 NOT_1645( .ZN(g7590), .A(g1155) );
  INV_X1 NOT_1646( .ZN(g7591), .A(g1496) );
  INV_X1 NOT_1647( .ZN(g7592), .A(g2540) );
  INV_X1 NOT_1648( .ZN(g7593), .A(g2571) );
  INV_X1 NOT_1649( .ZN(g7594), .A(g2165) );
  INV_X1 NOT_1650( .ZN(g7595), .A(g2900) );
  INV_X1 NOT_1651( .ZN(g7600), .A(g2908) );
  INV_X1 NOT_1652( .ZN(g7603), .A(g3133) );
  INV_X1 NOT_1653( .ZN(g7604), .A(g471) );
  INV_X1 NOT_1654( .ZN(g7605), .A(g1849) );
  INV_X1 NOT_1655( .ZN(g7606), .A(g2190) );
  INV_X1 NOT_1656( .ZN(g7607), .A(g2924) );
  INV_X1 NOT_1657( .ZN(g7610), .A(g312) );
  INV_X1 NOT_1658( .ZN(g7613), .A(g1158) );
  INV_X1 NOT_1659( .ZN(g7614), .A(g2543) );
  INV_X1 NOT_1660( .ZN(g7615), .A(g3123) );
  INV_X1 NOT_1661( .ZN(g7616), .A(g313) );
  INV_X1 NOT_1662( .ZN(g7619), .A(g999) );
  INV_X1 NOT_1663( .ZN(g7622), .A(g1852) );
  INV_X1 NOT_1664( .ZN(g7623), .A(g314) );
  INV_X1 NOT_1665( .ZN(g7626), .A(g315) );
  INV_X1 NOT_1666( .ZN(g7629), .A(g403) );
  INV_X1 NOT_1667( .ZN(g7632), .A(g1000) );
  INV_X1 NOT_1668( .ZN(g7635), .A(g1693) );
  INV_X1 NOT_1669( .ZN(g7638), .A(g2546) );
  INV_X1 NOT_1670( .ZN(g7639), .A(g3094) );
  INV_X1 NOT_1671( .ZN(g7642), .A(g3125) );
  INV_X1 NOT_1672( .ZN(g7643), .A(g316) );
  INV_X1 NOT_1673( .ZN(g7646), .A(g318) );
  INV_X1 NOT_1674( .ZN(g7649), .A(g404) );
  INV_X1 NOT_1675( .ZN(g7652), .A(g1001) );
  INV_X1 NOT_1676( .ZN(g7655), .A(g1002) );
  INV_X1 NOT_1677( .ZN(g7658), .A(g1090) );
  INV_X1 NOT_1678( .ZN(g7661), .A(g1694) );
  INV_X1 NOT_1679( .ZN(g7664), .A(g2387) );
  INV_X1 NOT_1680( .ZN(g7667), .A(g3095) );
  INV_X1 NOT_1681( .ZN(g7670), .A(g317) );
  INV_X1 NOT_1682( .ZN(g7673), .A(g319) );
  INV_X1 NOT_1683( .ZN(g7676), .A(g402) );
  INV_X1 NOT_1684( .ZN(g7679), .A(g1003) );
  INV_X1 NOT_1685( .ZN(g7682), .A(g1005) );
  INV_X1 NOT_1686( .ZN(g7685), .A(g1091) );
  INV_X1 NOT_1687( .ZN(g7688), .A(g1695) );
  INV_X1 NOT_1688( .ZN(g7691), .A(g1696) );
  INV_X1 NOT_1689( .ZN(g7694), .A(g1784) );
  INV_X1 NOT_1690( .ZN(g7697), .A(g2388) );
  INV_X1 NOT_1691( .ZN(g7700), .A(g3096) );
  INV_X1 NOT_1692( .ZN(g7703), .A(g320) );
  INV_X1 NOT_1693( .ZN(g7706), .A(g1004) );
  INV_X1 NOT_1694( .ZN(g7709), .A(g1006) );
  INV_X1 NOT_1695( .ZN(g7712), .A(g1089) );
  INV_X1 NOT_1696( .ZN(g7715), .A(g1697) );
  INV_X1 NOT_1697( .ZN(g7718), .A(g1699) );
  INV_X1 NOT_1698( .ZN(g7721), .A(g1785) );
  INV_X1 NOT_1699( .ZN(g7724), .A(g2389) );
  INV_X1 NOT_1700( .ZN(g7727), .A(g2390) );
  INV_X1 NOT_1701( .ZN(g7730), .A(g2478) );
  INV_X1 NOT_1702( .ZN(g7733), .A(g1007) );
  INV_X1 NOT_1703( .ZN(g7736), .A(g1698) );
  INV_X1 NOT_1704( .ZN(g7739), .A(g1700) );
  INV_X1 NOT_1705( .ZN(g7742), .A(g1783) );
  INV_X1 NOT_1706( .ZN(g7745), .A(g2391) );
  INV_X1 NOT_1707( .ZN(g7748), .A(g2393) );
  INV_X4 NOT_1708( .ZN(g7751), .A(g2479) );
  INV_X4 NOT_1709( .ZN(g7754), .A(g322) );
  INV_X4 NOT_1710( .ZN(g7757), .A(g1701) );
  INV_X4 NOT_1711( .ZN(g7760), .A(g2392) );
  INV_X1 NOT_1712( .ZN(g7763), .A(g2394) );
  INV_X1 NOT_1713( .ZN(g7766), .A(g2477) );
  INV_X1 NOT_1714( .ZN(g7769), .A(g323) );
  INV_X1 NOT_1715( .ZN(g7772), .A(g659) );
  INV_X1 NOT_1716( .ZN(g7776), .A(g1009) );
  INV_X1 NOT_1717( .ZN(g7779), .A(g2395) );
  INV_X1 NOT_1718( .ZN(g7782), .A(g321) );
  INV_X1 NOT_1719( .ZN(g7785), .A(g1010) );
  INV_X1 NOT_1720( .ZN(g7788), .A(g1345) );
  INV_X1 NOT_1721( .ZN(g7792), .A(g1703) );
  INV_X1 NOT_1722( .ZN(g7796), .A(g1008) );
  INV_X1 NOT_1723( .ZN(g7799), .A(g1704) );
  INV_X1 NOT_1724( .ZN(g7802), .A(g2039) );
  INV_X1 NOT_1725( .ZN(g7806), .A(g2397) );
  INV_X1 NOT_1726( .ZN(g7809), .A(g1702) );
  INV_X1 NOT_1727( .ZN(g7812), .A(g2398) );
  INV_X1 NOT_1728( .ZN(g7815), .A(g2733) );
  INV_X1 NOT_1729( .ZN(g7819), .A(g479) );
  INV_X1 NOT_1730( .ZN(g7822), .A(g510) );
  INV_X1 NOT_1731( .ZN(g7823), .A(g2396) );
  INV_X1 NOT_1732( .ZN(g7826), .A(g2987) );
  INV_X1 NOT_1733( .ZN(g7827), .A(g478) );
  INV_X1 NOT_1734( .ZN(g7830), .A(g1166) );
  INV_X1 NOT_1735( .ZN(g7833), .A(g1196) );
  INV_X1 NOT_1736( .ZN(g7834), .A(g2953) );
  INV_X1 NOT_1737( .ZN(g7837), .A(g3044) );
  INV_X1 NOT_1738( .ZN(g7838), .A(g477) );
  INV_X1 NOT_1739( .ZN(g7841), .A(g630) );
  INV_X1 NOT_1740( .ZN(g7842), .A(g1165) );
  INV_X1 NOT_1741( .ZN(g7845), .A(g1860) );
  INV_X1 NOT_1742( .ZN(g7848), .A(g1890) );
  INV_X1 NOT_1743( .ZN(g7849), .A(g2956) );
  INV_X1 NOT_1744( .ZN(g7852), .A(g2981) );
  INV_X1 NOT_1745( .ZN(g7856), .A(g3045) );
  INV_X1 NOT_1746( .ZN(g7857), .A(g3055) );
  INV_X1 NOT_1747( .ZN(g7858), .A(g1164) );
  INV_X1 NOT_1748( .ZN(g7861), .A(g1316) );
  INV_X1 NOT_1749( .ZN(g7862), .A(g1859) );
  INV_X1 NOT_1750( .ZN(g7865), .A(g2554) );
  INV_X1 NOT_1751( .ZN(g7868), .A(g2584) );
  INV_X1 NOT_1752( .ZN(g7869), .A(g2959) );
  INV_X1 NOT_1753( .ZN(g7872), .A(g2874) );
  INV_X1 NOT_1754( .ZN(g7877), .A(g3046) );
  INV_X1 NOT_1755( .ZN(g7878), .A(g3056) );
  INV_X1 NOT_1756( .ZN(g7879), .A(g3065) );
  INV_X1 NOT_1757( .ZN(g7880), .A(g3201) );
  INV_X1 NOT_1758( .ZN(g7888), .A(g1858) );
  INV_X1 NOT_1759( .ZN(g7891), .A(g2010) );
  INV_X1 NOT_1760( .ZN(g7892), .A(g2553) );
  INV_X1 NOT_1761( .ZN(g7897), .A(g3047) );
  INV_X1 NOT_1762( .ZN(g7898), .A(g3057) );
  INV_X1 NOT_1763( .ZN(g7899), .A(g3066) );
  INV_X1 NOT_1764( .ZN(g7900), .A(g3075) );
  INV_X1 NOT_1765( .ZN(II15222), .A(g3151) );
  INV_X1 NOT_1766( .ZN(g7901), .A(II15222) );
  INV_X1 NOT_1767( .ZN(g7906), .A(g488) );
  INV_X1 NOT_1768( .ZN(II15226), .A(g474) );
  INV_X1 NOT_1769( .ZN(g7909), .A(II15226) );
  INV_X1 NOT_1770( .ZN(g7910), .A(g474) );
  INV_X1 NOT_1771( .ZN(II15230), .A(g499) );
  INV_X1 NOT_1772( .ZN(g7911), .A(II15230) );
  INV_X1 NOT_1773( .ZN(g7912), .A(g2552) );
  INV_X1 NOT_1774( .ZN(g7915), .A(g2704) );
  INV_X1 NOT_1775( .ZN(g7916), .A(g2935) );
  INV_X1 NOT_1776( .ZN(g7919), .A(g2963) );
  INV_X1 NOT_1777( .ZN(g7924), .A(g3048) );
  INV_X1 NOT_1778( .ZN(g7925), .A(g3058) );
  INV_X1 NOT_1779( .ZN(g7926), .A(g3067) );
  INV_X1 NOT_1780( .ZN(g7927), .A(g3076) );
  INV_X1 NOT_1781( .ZN(g7928), .A(g3204) );
  INV_X1 NOT_1782( .ZN(II15256), .A(g2950) );
  INV_X1 NOT_1783( .ZN(g7936), .A(II15256) );
  INV_X1 NOT_1784( .ZN(g7949), .A(g165) );
  INV_X1 NOT_1785( .ZN(g7950), .A(g142) );
  INV_X1 NOT_1786( .ZN(g7953), .A(g487) );
  INV_X1 NOT_1787( .ZN(II15262), .A(g481) );
  INV_X1 NOT_1788( .ZN(g7956), .A(II15262) );
  INV_X1 NOT_1789( .ZN(g7957), .A(g481) );
  INV_X1 NOT_1790( .ZN(g7958), .A(g1175) );
  INV_X1 NOT_1791( .ZN(II15267), .A(g1161) );
  INV_X1 NOT_1792( .ZN(g7961), .A(II15267) );
  INV_X1 NOT_1793( .ZN(g7962), .A(g1161) );
  INV_X1 NOT_1794( .ZN(II15271), .A(g1186) );
  INV_X1 NOT_1795( .ZN(g7963), .A(II15271) );
  INV_X1 NOT_1796( .ZN(g7964), .A(g2938) );
  INV_X1 NOT_1797( .ZN(g7967), .A(g2966) );
  INV_X1 NOT_1798( .ZN(g7971), .A(g3049) );
  INV_X1 NOT_1799( .ZN(g7972), .A(g3059) );
  INV_X1 NOT_1800( .ZN(g7973), .A(g3068) );
  INV_X1 NOT_1801( .ZN(g7974), .A(g3077) );
  INV_X1 NOT_1802( .ZN(g7975), .A(g39) );
  INV_X1 NOT_1803( .ZN(II15288), .A(g3109) );
  INV_X1 NOT_1804( .ZN(g7976), .A(II15288) );
  INV_X1 NOT_1805( .ZN(g7989), .A(g3191) );
  INV_X1 NOT_1806( .ZN(g7990), .A(g143) );
  INV_X1 NOT_1807( .ZN(g7993), .A(g145) );
  INV_X1 NOT_1808( .ZN(g7996), .A(g486) );
  INV_X1 NOT_1809( .ZN(g7999), .A(g485) );
  INV_X1 NOT_1810( .ZN(g8000), .A(g853) );
  INV_X1 NOT_1811( .ZN(g8001), .A(g830) );
  INV_X1 NOT_1812( .ZN(g8004), .A(g1174) );
  INV_X1 NOT_1813( .ZN(II15299), .A(g1168) );
  INV_X1 NOT_1814( .ZN(g8007), .A(II15299) );
  INV_X1 NOT_1815( .ZN(g8008), .A(g1168) );
  INV_X1 NOT_1816( .ZN(g8009), .A(g1869) );
  INV_X1 NOT_1817( .ZN(II15304), .A(g1855) );
  INV_X1 NOT_1818( .ZN(g8012), .A(II15304) );
  INV_X1 NOT_1819( .ZN(g8013), .A(g1855) );
  INV_X1 NOT_1820( .ZN(II15308), .A(g1880) );
  INV_X1 NOT_1821( .ZN(g8014), .A(II15308) );
  INV_X1 NOT_1822( .ZN(g8015), .A(g2941) );
  INV_X1 NOT_1823( .ZN(g8018), .A(g2969) );
  INV_X1 NOT_1824( .ZN(II15313), .A(g2930) );
  INV_X4 NOT_1825( .ZN(g8021), .A(II15313) );
  INV_X4 NOT_1826( .ZN(g8022), .A(g2930) );
  INV_X4 NOT_1827( .ZN(II15317), .A(g2842) );
  INV_X4 NOT_1828( .ZN(g8023), .A(II15317) );
  INV_X1 NOT_1829( .ZN(g8024), .A(g2842) );
  INV_X1 NOT_1830( .ZN(g8025), .A(g3050) );
  INV_X1 NOT_1831( .ZN(g8026), .A(g3060) );
  INV_X1 NOT_1832( .ZN(g8027), .A(g3069) );
  INV_X1 NOT_1833( .ZN(g8028), .A(g3078) );
  INV_X1 NOT_1834( .ZN(g8029), .A(g3083) );
  INV_X1 NOT_1835( .ZN(II15326), .A(g3117) );
  INV_X1 NOT_1836( .ZN(g8030), .A(II15326) );
  INV_X1 NOT_1837( .ZN(II15329), .A(g3117) );
  INV_X1 NOT_1838( .ZN(g8031), .A(II15329) );
  INV_X1 NOT_1839( .ZN(g8044), .A(g3194) );
  INV_X1 NOT_1840( .ZN(g8045), .A(g3207) );
  INV_X1 NOT_1841( .ZN(g8053), .A(g141) );
  INV_X1 NOT_1842( .ZN(g8056), .A(g146) );
  INV_X1 NOT_1843( .ZN(g8059), .A(g148) );
  INV_X1 NOT_1844( .ZN(g8062), .A(g169) );
  INV_X1 NOT_1845( .ZN(g8065), .A(g831) );
  INV_X1 NOT_1846( .ZN(g8068), .A(g833) );
  INV_X1 NOT_1847( .ZN(g8071), .A(g1173) );
  INV_X1 NOT_1848( .ZN(g8074), .A(g1172) );
  INV_X1 NOT_1849( .ZN(g8075), .A(g1547) );
  INV_X1 NOT_1850( .ZN(g8076), .A(g1524) );
  INV_X1 NOT_1851( .ZN(g8079), .A(g1868) );
  INV_X1 NOT_1852( .ZN(II15345), .A(g1862) );
  INV_X1 NOT_1853( .ZN(g8082), .A(II15345) );
  INV_X1 NOT_1854( .ZN(g8083), .A(g1862) );
  INV_X1 NOT_1855( .ZN(g8084), .A(g2563) );
  INV_X1 NOT_1856( .ZN(II15350), .A(g2549) );
  INV_X1 NOT_1857( .ZN(g8087), .A(II15350) );
  INV_X1 NOT_1858( .ZN(g8088), .A(g2549) );
  INV_X1 NOT_1859( .ZN(II15354), .A(g2574) );
  INV_X1 NOT_1860( .ZN(g8089), .A(II15354) );
  INV_X1 NOT_1861( .ZN(g8090), .A(g2944) );
  INV_X1 NOT_1862( .ZN(g8093), .A(g2972) );
  INV_X1 NOT_1863( .ZN(II15359), .A(g2858) );
  INV_X1 NOT_1864( .ZN(g8096), .A(II15359) );
  INV_X1 NOT_1865( .ZN(g8097), .A(g2858) );
  INV_X1 NOT_1866( .ZN(g8098), .A(g3051) );
  INV_X1 NOT_1867( .ZN(g8099), .A(g3061) );
  INV_X1 NOT_1868( .ZN(g8100), .A(g3070) );
  INV_X1 NOT_1869( .ZN(g8101), .A(g2997) );
  INV_X1 NOT_1870( .ZN(g8102), .A(g27) );
  INV_X1 NOT_1871( .ZN(g8103), .A(g185) );
  INV_X1 NOT_1872( .ZN(II15369), .A(g3129) );
  INV_X1 NOT_1873( .ZN(g8106), .A(II15369) );
  INV_X1 NOT_1874( .ZN(II15372), .A(g3129) );
  INV_X1 NOT_1875( .ZN(g8107), .A(II15372) );
  INV_X1 NOT_1876( .ZN(g8120), .A(g3197) );
  INV_X1 NOT_1877( .ZN(g8123), .A(g144) );
  INV_X1 NOT_1878( .ZN(g8126), .A(g149) );
  INV_X1 NOT_1879( .ZN(g8129), .A(g151) );
  INV_X1 NOT_1880( .ZN(g8132), .A(g170) );
  INV_X1 NOT_1881( .ZN(g8135), .A(g172) );
  INV_X1 NOT_1882( .ZN(g8138), .A(g829) );
  INV_X1 NOT_1883( .ZN(g8141), .A(g834) );
  INV_X1 NOT_1884( .ZN(g8144), .A(g836) );
  INV_X1 NOT_1885( .ZN(g8147), .A(g857) );
  INV_X1 NOT_1886( .ZN(g8150), .A(g1525) );
  INV_X1 NOT_1887( .ZN(g8153), .A(g1527) );
  INV_X1 NOT_1888( .ZN(g8156), .A(g1867) );
  INV_X4 NOT_1889( .ZN(g8159), .A(g1866) );
  INV_X1 NOT_1890( .ZN(g8160), .A(g2241) );
  INV_X1 NOT_1891( .ZN(g8161), .A(g2218) );
  INV_X1 NOT_1892( .ZN(g8164), .A(g2562) );
  INV_X1 NOT_1893( .ZN(II15392), .A(g2556) );
  INV_X1 NOT_1894( .ZN(g8167), .A(II15392) );
  INV_X1 NOT_1895( .ZN(g8168), .A(g2556) );
  INV_X1 NOT_1896( .ZN(g8169), .A(g2947) );
  INV_X1 NOT_1897( .ZN(g8172), .A(g2975) );
  INV_X1 NOT_1898( .ZN(II15398), .A(g2845) );
  INV_X1 NOT_1899( .ZN(g8175), .A(II15398) );
  INV_X1 NOT_1900( .ZN(g8176), .A(g2845) );
  INV_X1 NOT_1901( .ZN(g8177), .A(g3043) );
  INV_X1 NOT_1902( .ZN(g8178), .A(g3052) );
  INV_X1 NOT_1903( .ZN(g8179), .A(g3062) );
  INV_X1 NOT_1904( .ZN(g8180), .A(g3071) );
  INV_X1 NOT_1905( .ZN(g8181), .A(g48) );
  INV_X1 NOT_1906( .ZN(g8182), .A(g3198) );
  INV_X1 NOT_1907( .ZN(g8183), .A(g3188) );
  INV_X1 NOT_1908( .ZN(g8191), .A(g147) );
  INV_X1 NOT_1909( .ZN(g8194), .A(g152) );
  INV_X1 NOT_1910( .ZN(g8197), .A(g154) );
  INV_X1 NOT_1911( .ZN(g8200), .A(g168) );
  INV_X1 NOT_1912( .ZN(g8203), .A(g173) );
  INV_X1 NOT_1913( .ZN(g8206), .A(g175) );
  INV_X1 NOT_1914( .ZN(g8209), .A(g832) );
  INV_X1 NOT_1915( .ZN(g8212), .A(g837) );
  INV_X1 NOT_1916( .ZN(g8215), .A(g839) );
  INV_X1 NOT_1917( .ZN(g8218), .A(g858) );
  INV_X1 NOT_1918( .ZN(g8221), .A(g860) );
  INV_X1 NOT_1919( .ZN(g8224), .A(g1523) );
  INV_X1 NOT_1920( .ZN(g8227), .A(g1528) );
  INV_X1 NOT_1921( .ZN(g8230), .A(g1530) );
  INV_X1 NOT_1922( .ZN(g8233), .A(g1551) );
  INV_X1 NOT_1923( .ZN(g8236), .A(g2219) );
  INV_X1 NOT_1924( .ZN(g8239), .A(g2221) );
  INV_X1 NOT_1925( .ZN(g8242), .A(g2561) );
  INV_X1 NOT_1926( .ZN(g8245), .A(g2560) );
  INV_X1 NOT_1927( .ZN(g8246), .A(g2978) );
  INV_X1 NOT_1928( .ZN(II15429), .A(g2833) );
  INV_X1 NOT_1929( .ZN(g8249), .A(II15429) );
  INV_X1 NOT_1930( .ZN(g8250), .A(g2833) );
  INV_X1 NOT_1931( .ZN(II15433), .A(g2861) );
  INV_X1 NOT_1932( .ZN(g8251), .A(II15433) );
  INV_X1 NOT_1933( .ZN(g8252), .A(g2861) );
  INV_X1 NOT_1934( .ZN(g8253), .A(g3053) );
  INV_X1 NOT_1935( .ZN(g8254), .A(g3063) );
  INV_X1 NOT_1936( .ZN(g8255), .A(g3072) );
  INV_X1 NOT_1937( .ZN(g8256), .A(g30) );
  INV_X1 NOT_1938( .ZN(g8257), .A(g3201) );
  INV_X1 NOT_1939( .ZN(II15442), .A(g3235) );
  INV_X1 NOT_1940( .ZN(g8258), .A(II15442) );
  INV_X1 NOT_1941( .ZN(II15445), .A(g3236) );
  INV_X1 NOT_1942( .ZN(g8259), .A(II15445) );
  INV_X1 NOT_1943( .ZN(II15448), .A(g3237) );
  INV_X1 NOT_1944( .ZN(g8260), .A(II15448) );
  INV_X1 NOT_1945( .ZN(II15451), .A(g3238) );
  INV_X1 NOT_1946( .ZN(g8261), .A(II15451) );
  INV_X1 NOT_1947( .ZN(II15454), .A(g3239) );
  INV_X1 NOT_1948( .ZN(g8262), .A(II15454) );
  INV_X1 NOT_1949( .ZN(II15457), .A(g3240) );
  INV_X1 NOT_1950( .ZN(g8263), .A(II15457) );
  INV_X1 NOT_1951( .ZN(II15460), .A(g3241) );
  INV_X1 NOT_1952( .ZN(g8264), .A(II15460) );
  INV_X1 NOT_1953( .ZN(II15463), .A(g3242) );
  INV_X1 NOT_1954( .ZN(g8265), .A(II15463) );
  INV_X1 NOT_1955( .ZN(II15466), .A(g3243) );
  INV_X1 NOT_1956( .ZN(g8266), .A(II15466) );
  INV_X1 NOT_1957( .ZN(II15469), .A(g3244) );
  INV_X1 NOT_1958( .ZN(g8267), .A(II15469) );
  INV_X1 NOT_1959( .ZN(II15472), .A(g3245) );
  INV_X1 NOT_1960( .ZN(g8268), .A(II15472) );
  INV_X1 NOT_1961( .ZN(II15475), .A(g3246) );
  INV_X1 NOT_1962( .ZN(g8269), .A(II15475) );
  INV_X1 NOT_1963( .ZN(II15478), .A(g3247) );
  INV_X1 NOT_1964( .ZN(g8270), .A(II15478) );
  INV_X1 NOT_1965( .ZN(II15481), .A(g3248) );
  INV_X1 NOT_1966( .ZN(g8271), .A(II15481) );
  INV_X1 NOT_1967( .ZN(II15484), .A(g3249) );
  INV_X1 NOT_1968( .ZN(g8272), .A(II15484) );
  INV_X1 NOT_1969( .ZN(II15487), .A(g3250) );
  INV_X1 NOT_1970( .ZN(g8273), .A(II15487) );
  INV_X1 NOT_1971( .ZN(II15490), .A(g3251) );
  INV_X1 NOT_1972( .ZN(g8274), .A(II15490) );
  INV_X1 NOT_1973( .ZN(II15493), .A(g3252) );
  INV_X1 NOT_1974( .ZN(g8275), .A(II15493) );
  INV_X1 NOT_1975( .ZN(g8276), .A(g3253) );
  INV_X1 NOT_1976( .ZN(g8277), .A(g3305) );
  INV_X1 NOT_1977( .ZN(g8278), .A(g3337) );
  INV_X1 NOT_1978( .ZN(II15499), .A(g7911) );
  INV_X1 NOT_1979( .ZN(g8284), .A(II15499) );
  INV_X1 NOT_1980( .ZN(g8285), .A(g3365) );
  INV_X1 NOT_1981( .ZN(g8286), .A(g3461) );
  INV_X1 NOT_1982( .ZN(g8287), .A(g3493) );
  INV_X1 NOT_1983( .ZN(II15505), .A(g7963) );
  INV_X1 NOT_1984( .ZN(g8293), .A(II15505) );
  INV_X1 NOT_1985( .ZN(g8294), .A(g3521) );
  INV_X1 NOT_1986( .ZN(g8295), .A(g3617) );
  INV_X1 NOT_1987( .ZN(g8296), .A(g3649) );
  INV_X1 NOT_1988( .ZN(II15511), .A(g8014) );
  INV_X1 NOT_1989( .ZN(g8302), .A(II15511) );
  INV_X4 NOT_1990( .ZN(g8303), .A(g3677) );
  INV_X4 NOT_1991( .ZN(g8304), .A(g3773) );
  INV_X1 NOT_1992( .ZN(g8305), .A(g3805) );
  INV_X1 NOT_1993( .ZN(II15517), .A(g8089) );
  INV_X1 NOT_1994( .ZN(g8311), .A(II15517) );
  INV_X1 NOT_1995( .ZN(g8312), .A(g3833) );
  INV_X1 NOT_1996( .ZN(g8313), .A(g3897) );
  INV_X1 NOT_1997( .ZN(g8317), .A(g3919) );
  INV_X1 NOT_1998( .ZN(II15523), .A(g3254) );
  INV_X1 NOT_1999( .ZN(g8321), .A(II15523) );
  INV_X1 NOT_2000( .ZN(II15526), .A(g6314) );
  INV_X1 NOT_2001( .ZN(g8324), .A(II15526) );
  INV_X1 NOT_2002( .ZN(II15532), .A(g3410) );
  INV_X1 NOT_2003( .ZN(g8330), .A(II15532) );
  INV_X1 NOT_2004( .ZN(II15535), .A(g6519) );
  INV_X1 NOT_2005( .ZN(g8333), .A(II15535) );
  INV_X1 NOT_2006( .ZN(II15538), .A(g6369) );
  INV_X1 NOT_2007( .ZN(g8336), .A(II15538) );
  INV_X1 NOT_2008( .ZN(II15543), .A(g3410) );
  INV_X1 NOT_2009( .ZN(g8341), .A(II15543) );
  INV_X1 NOT_2010( .ZN(II15546), .A(g6783) );
  INV_X1 NOT_2011( .ZN(g8344), .A(II15546) );
  INV_X1 NOT_2012( .ZN(II15549), .A(g6574) );
  INV_X1 NOT_2013( .ZN(g8347), .A(II15549) );
  INV_X1 NOT_2014( .ZN(II15553), .A(g3566) );
  INV_X1 NOT_2015( .ZN(g8351), .A(II15553) );
  INV_X1 NOT_2016( .ZN(II15556), .A(g6783) );
  INV_X1 NOT_2017( .ZN(g8354), .A(II15556) );
  INV_X1 NOT_2018( .ZN(II15559), .A(g7015) );
  INV_X1 NOT_2019( .ZN(g8357), .A(II15559) );
  INV_X1 NOT_2020( .ZN(II15562), .A(g5778) );
  INV_X1 NOT_2021( .ZN(g8360), .A(II15562) );
  INV_X1 NOT_2022( .ZN(II15565), .A(g6838) );
  INV_X1 NOT_2023( .ZN(g8363), .A(II15565) );
  INV_X1 NOT_2024( .ZN(II15568), .A(g3722) );
  INV_X1 NOT_2025( .ZN(g8366), .A(II15568) );
  INV_X1 NOT_2026( .ZN(II15571), .A(g7085) );
  INV_X1 NOT_2027( .ZN(g8369), .A(II15571) );
  INV_X1 NOT_2028( .ZN(II15574), .A(g6838) );
  INV_X1 NOT_2029( .ZN(g8372), .A(II15574) );
  INV_X1 NOT_2030( .ZN(II15577), .A(g7265) );
  INV_X1 NOT_2031( .ZN(g8375), .A(II15577) );
  INV_X1 NOT_2032( .ZN(II15580), .A(g5837) );
  INV_X1 NOT_2033( .ZN(g8378), .A(II15580) );
  INV_X1 NOT_2034( .ZN(II15584), .A(g3254) );
  INV_X1 NOT_2035( .ZN(g8382), .A(II15584) );
  INV_X1 NOT_2036( .ZN(II15590), .A(g3410) );
  INV_X1 NOT_2037( .ZN(g8388), .A(II15590) );
  INV_X1 NOT_2038( .ZN(II15593), .A(g6519) );
  INV_X1 NOT_2039( .ZN(g8391), .A(II15593) );
  INV_X1 NOT_2040( .ZN(II15599), .A(g3566) );
  INV_X1 NOT_2041( .ZN(g8397), .A(II15599) );
  INV_X1 NOT_2042( .ZN(II15602), .A(g6783) );
  INV_X1 NOT_2043( .ZN(g8400), .A(II15602) );
  INV_X1 NOT_2044( .ZN(II15605), .A(g6574) );
  INV_X1 NOT_2045( .ZN(g8403), .A(II15605) );
  INV_X1 NOT_2046( .ZN(II15610), .A(g3566) );
  INV_X1 NOT_2047( .ZN(g8408), .A(II15610) );
  INV_X1 NOT_2048( .ZN(II15613), .A(g7085) );
  INV_X1 NOT_2049( .ZN(g8411), .A(II15613) );
  INV_X1 NOT_2050( .ZN(II15616), .A(g6838) );
  INV_X1 NOT_2051( .ZN(g8414), .A(II15616) );
  INV_X16 NOT_2052( .ZN(II15620), .A(g3722) );
  INV_X16 NOT_2053( .ZN(g8418), .A(II15620) );
  INV_X1 NOT_2054( .ZN(II15623), .A(g7085) );
  INV_X1 NOT_2055( .ZN(g8421), .A(II15623) );
  INV_X1 NOT_2056( .ZN(II15626), .A(g7265) );
  INV_X1 NOT_2057( .ZN(g8424), .A(II15626) );
  INV_X1 NOT_2058( .ZN(II15629), .A(g5837) );
  INV_X1 NOT_2059( .ZN(g8427), .A(II15629) );
  INV_X1 NOT_2060( .ZN(II15636), .A(g3410) );
  INV_X1 NOT_2061( .ZN(g8434), .A(II15636) );
  INV_X1 NOT_2062( .ZN(II15642), .A(g3566) );
  INV_X1 NOT_2063( .ZN(g8440), .A(II15642) );
  INV_X1 NOT_2064( .ZN(II15645), .A(g6783) );
  INV_X1 NOT_2065( .ZN(g8443), .A(II15645) );
  INV_X1 NOT_2066( .ZN(II15651), .A(g3722) );
  INV_X1 NOT_2067( .ZN(g8449), .A(II15651) );
  INV_X1 NOT_2068( .ZN(II15654), .A(g7085) );
  INV_X1 NOT_2069( .ZN(g8452), .A(II15654) );
  INV_X1 NOT_2070( .ZN(II15657), .A(g6838) );
  INV_X1 NOT_2071( .ZN(g8455), .A(II15657) );
  INV_X1 NOT_2072( .ZN(II15662), .A(g3722) );
  INV_X1 NOT_2073( .ZN(g8460), .A(II15662) );
  INV_X1 NOT_2074( .ZN(II15671), .A(g3566) );
  INV_X1 NOT_2075( .ZN(g8469), .A(II15671) );
  INV_X1 NOT_2076( .ZN(II15677), .A(g3722) );
  INV_X1 NOT_2077( .ZN(g8475), .A(II15677) );
  INV_X1 NOT_2078( .ZN(II15680), .A(g7085) );
  INV_X1 NOT_2079( .ZN(g8478), .A(II15680) );
  INV_X1 NOT_2080( .ZN(II15696), .A(g3722) );
  INV_X1 NOT_2081( .ZN(g8494), .A(II15696) );
  INV_X1 NOT_2082( .ZN(g8514), .A(g6139) );
  INV_X1 NOT_2083( .ZN(g8530), .A(g6156) );
  INV_X1 NOT_2084( .ZN(g8568), .A(g6230) );
  INV_X1 NOT_2085( .ZN(II15771), .A(g6000) );
  INV_X1 NOT_2086( .ZN(g8569), .A(II15771) );
  INV_X1 NOT_2087( .ZN(II15779), .A(g6000) );
  INV_X1 NOT_2088( .ZN(g8575), .A(II15779) );
  INV_X1 NOT_2089( .ZN(II15784), .A(g6000) );
  INV_X1 NOT_2090( .ZN(g8578), .A(II15784) );
  INV_X1 NOT_2091( .ZN(II15787), .A(g6000) );
  INV_X1 NOT_2092( .ZN(g8579), .A(II15787) );
  INV_X1 NOT_2093( .ZN(g8580), .A(g6281) );
  INV_X1 NOT_2094( .ZN(g8587), .A(g6418) );
  INV_X1 NOT_2095( .ZN(g8594), .A(g6623) );
  INV_X1 NOT_2096( .ZN(II15794), .A(g3338) );
  INV_X1 NOT_2097( .ZN(g8602), .A(II15794) );
  INV_X1 NOT_2098( .ZN(g8605), .A(g6887) );
  INV_X1 NOT_2099( .ZN(II15800), .A(g3494) );
  INV_X1 NOT_2100( .ZN(g8614), .A(II15800) );
  INV_X1 NOT_2101( .ZN(II15803), .A(g8107) );
  INV_X1 NOT_2102( .ZN(g8617), .A(II15803) );
  INV_X1 NOT_2103( .ZN(II15806), .A(g5550) );
  INV_X1 NOT_2104( .ZN(g8620), .A(II15806) );
  INV_X1 NOT_2105( .ZN(II15810), .A(g3338) );
  INV_X1 NOT_2106( .ZN(g8622), .A(II15810) );
  INV_X1 NOT_2107( .ZN(II15815), .A(g3650) );
  INV_X1 NOT_2108( .ZN(g8627), .A(II15815) );
  INV_X1 NOT_2109( .ZN(II15818), .A(g5596) );
  INV_X1 NOT_2110( .ZN(g8630), .A(II15818) );
  INV_X1 NOT_2111( .ZN(II15822), .A(g3494) );
  INV_X16 NOT_2112( .ZN(g8632), .A(II15822) );
  INV_X1 NOT_2113( .ZN(II15827), .A(g3806) );
  INV_X1 NOT_2114( .ZN(g8637), .A(II15827) );
  INV_X1 NOT_2115( .ZN(II15830), .A(g8031) );
  INV_X1 NOT_2116( .ZN(g8640), .A(II15830) );
  INV_X1 NOT_2117( .ZN(II15833), .A(g3338) );
  INV_X1 NOT_2118( .ZN(g8643), .A(II15833) );
  INV_X1 NOT_2119( .ZN(II15836), .A(g3366) );
  INV_X1 NOT_2120( .ZN(g8646), .A(II15836) );
  INV_X1 NOT_2121( .ZN(II15839), .A(g5613) );
  INV_X1 NOT_2122( .ZN(g8649), .A(II15839) );
  INV_X1 NOT_2123( .ZN(II15843), .A(g3650) );
  INV_X1 NOT_2124( .ZN(g8651), .A(II15843) );
  INV_X1 NOT_2125( .ZN(II15847), .A(g3878) );
  INV_X1 NOT_2126( .ZN(g8655), .A(II15847) );
  INV_X1 NOT_2127( .ZN(II15850), .A(g5627) );
  INV_X1 NOT_2128( .ZN(g8658), .A(II15850) );
  INV_X1 NOT_2129( .ZN(II15853), .A(g3494) );
  INV_X1 NOT_2130( .ZN(g8659), .A(II15853) );
  INV_X1 NOT_2131( .ZN(II15856), .A(g3522) );
  INV_X1 NOT_2132( .ZN(g8662), .A(II15856) );
  INV_X1 NOT_2133( .ZN(II15859), .A(g5638) );
  INV_X1 NOT_2134( .ZN(g8665), .A(II15859) );
  INV_X1 NOT_2135( .ZN(II15863), .A(g3806) );
  INV_X1 NOT_2136( .ZN(g8667), .A(II15863) );
  INV_X1 NOT_2137( .ZN(II15866), .A(g3878) );
  INV_X1 NOT_2138( .ZN(g8670), .A(II15866) );
  INV_X1 NOT_2139( .ZN(II15869), .A(g7976) );
  INV_X1 NOT_2140( .ZN(g8673), .A(II15869) );
  INV_X1 NOT_2141( .ZN(II15873), .A(g5655) );
  INV_X1 NOT_2142( .ZN(g8677), .A(II15873) );
  INV_X1 NOT_2143( .ZN(II15876), .A(g3650) );
  INV_X1 NOT_2144( .ZN(g8678), .A(II15876) );
  INV_X1 NOT_2145( .ZN(II15879), .A(g3678) );
  INV_X1 NOT_2146( .ZN(g8681), .A(II15879) );
  INV_X1 NOT_2147( .ZN(II15882), .A(g3878) );
  INV_X1 NOT_2148( .ZN(g8684), .A(II15882) );
  INV_X1 NOT_2149( .ZN(II15887), .A(g5693) );
  INV_X1 NOT_2150( .ZN(g8689), .A(II15887) );
  INV_X1 NOT_2151( .ZN(II15890), .A(g3806) );
  INV_X1 NOT_2152( .ZN(g8690), .A(II15890) );
  INV_X1 NOT_2153( .ZN(II15893), .A(g3834) );
  INV_X32 NOT_2154( .ZN(g8693), .A(II15893) );
  INV_X32 NOT_2155( .ZN(II15896), .A(g3878) );
  INV_X32 NOT_2156( .ZN(g8696), .A(II15896) );
  INV_X32 NOT_2157( .ZN(II15899), .A(g5626) );
  INV_X1 NOT_2158( .ZN(g8699), .A(II15899) );
  INV_X1 NOT_2159( .ZN(II15902), .A(g6486) );
  INV_X1 NOT_2160( .ZN(g8700), .A(II15902) );
  INV_X1 NOT_2161( .ZN(II15909), .A(g5745) );
  INV_X1 NOT_2162( .ZN(g8707), .A(II15909) );
  INV_X1 NOT_2163( .ZN(II15912), .A(g3878) );
  INV_X1 NOT_2164( .ZN(g8708), .A(II15912) );
  INV_X1 NOT_2165( .ZN(II15915), .A(g3878) );
  INV_X1 NOT_2166( .ZN(g8711), .A(II15915) );
  INV_X1 NOT_2167( .ZN(II15918), .A(g6643) );
  INV_X1 NOT_2168( .ZN(g8714), .A(II15918) );
  INV_X1 NOT_2169( .ZN(II15922), .A(g5654) );
  INV_X1 NOT_2170( .ZN(g8718), .A(II15922) );
  INV_X1 NOT_2171( .ZN(II15925), .A(g6751) );
  INV_X1 NOT_2172( .ZN(g8719), .A(II15925) );
  INV_X1 NOT_2173( .ZN(II15932), .A(g5423) );
  INV_X1 NOT_2174( .ZN(g8726), .A(II15932) );
  INV_X1 NOT_2175( .ZN(II15935), .A(g3878) );
  INV_X1 NOT_2176( .ZN(g8745), .A(II15935) );
  INV_X1 NOT_2177( .ZN(II15938), .A(g3338) );
  INV_X1 NOT_2178( .ZN(g8748), .A(II15938) );
  INV_X1 NOT_2179( .ZN(II15942), .A(g6945) );
  INV_X1 NOT_2180( .ZN(g8752), .A(II15942) );
  INV_X1 NOT_2181( .ZN(II15946), .A(g5692) );
  INV_X1 NOT_2182( .ZN(g8756), .A(II15946) );
  INV_X1 NOT_2183( .ZN(II15949), .A(g7053) );
  INV_X1 NOT_2184( .ZN(g8757), .A(II15949) );
  INV_X1 NOT_2185( .ZN(II15955), .A(g3878) );
  INV_X1 NOT_2186( .ZN(g8763), .A(II15955) );
  INV_X1 NOT_2187( .ZN(II15958), .A(g3878) );
  INV_X1 NOT_2188( .ZN(g8766), .A(II15958) );
  INV_X1 NOT_2189( .ZN(II15961), .A(g6051) );
  INV_X1 NOT_2190( .ZN(g8769), .A(II15961) );
  INV_X1 NOT_2191( .ZN(II15964), .A(g7554) );
  INV_X1 NOT_2192( .ZN(g8770), .A(II15964) );
  INV_X1 NOT_2193( .ZN(II15967), .A(g3494) );
  INV_X1 NOT_2194( .ZN(g8771), .A(II15967) );
  INV_X1 NOT_2195( .ZN(II15971), .A(g7195) );
  INV_X1 NOT_2196( .ZN(g8775), .A(II15971) );
  INV_X1 NOT_2197( .ZN(II15975), .A(g5744) );
  INV_X1 NOT_2198( .ZN(g8779), .A(II15975) );
  INV_X1 NOT_2199( .ZN(II15978), .A(g7303) );
  INV_X1 NOT_2200( .ZN(g8780), .A(II15978) );
  INV_X1 NOT_2201( .ZN(II15983), .A(g3878) );
  INV_X1 NOT_2202( .ZN(g8785), .A(II15983) );
  INV_X1 NOT_2203( .ZN(II15986), .A(g3878) );
  INV_X1 NOT_2204( .ZN(g8788), .A(II15986) );
  INV_X1 NOT_2205( .ZN(II15989), .A(g6053) );
  INV_X1 NOT_2206( .ZN(g8791), .A(II15989) );
  INV_X1 NOT_2207( .ZN(II15992), .A(g6055) );
  INV_X1 NOT_2208( .ZN(g8792), .A(II15992) );
  INV_X1 NOT_2209( .ZN(II15995), .A(g7577) );
  INV_X1 NOT_2210( .ZN(g8793), .A(II15995) );
  INV_X1 NOT_2211( .ZN(II15998), .A(g3650) );
  INV_X1 NOT_2212( .ZN(g8794), .A(II15998) );
  INV_X1 NOT_2213( .ZN(II16002), .A(g7391) );
  INV_X1 NOT_2214( .ZN(g8798), .A(II16002) );
  INV_X1 NOT_2215( .ZN(II16006), .A(g3878) );
  INV_X1 NOT_2216( .ZN(g8802), .A(II16006) );
  INV_X1 NOT_2217( .ZN(II16009), .A(g3878) );
  INV_X1 NOT_2218( .ZN(g8805), .A(II16009) );
  INV_X1 NOT_2219( .ZN(II16012), .A(g5390) );
  INV_X1 NOT_2220( .ZN(g8808), .A(II16012) );
  INV_X1 NOT_2221( .ZN(II16015), .A(g6056) );
  INV_X1 NOT_2222( .ZN(g8809), .A(II16015) );
  INV_X1 NOT_2223( .ZN(II16018), .A(g6058) );
  INV_X1 NOT_2224( .ZN(g8810), .A(II16018) );
  INV_X1 NOT_2225( .ZN(II16021), .A(g6060) );
  INV_X1 NOT_2226( .ZN(g8811), .A(II16021) );
  INV_X1 NOT_2227( .ZN(II16024), .A(g7591) );
  INV_X1 NOT_2228( .ZN(g8812), .A(II16024) );
  INV_X1 NOT_2229( .ZN(II16027), .A(g3806) );
  INV_X1 NOT_2230( .ZN(g8813), .A(II16027) );
  INV_X1 NOT_2231( .ZN(II16031), .A(g3878) );
  INV_X1 NOT_2232( .ZN(g8817), .A(II16031) );
  INV_X1 NOT_2233( .ZN(II16034), .A(g5396) );
  INV_X1 NOT_2234( .ZN(g8820), .A(II16034) );
  INV_X1 NOT_2235( .ZN(II16037), .A(g6061) );
  INV_X1 NOT_2236( .ZN(g8821), .A(II16037) );
  INV_X1 NOT_2237( .ZN(g8822), .A(g4602) );
  INV_X1 NOT_2238( .ZN(II16041), .A(g6486) );
  INV_X1 NOT_2239( .ZN(g8823), .A(II16041) );
  INV_X1 NOT_2240( .ZN(II16044), .A(g5397) );
  INV_X1 NOT_2241( .ZN(g8824), .A(II16044) );
  INV_X1 NOT_2242( .ZN(II16047), .A(g6063) );
  INV_X1 NOT_2243( .ZN(g8825), .A(II16047) );
  INV_X1 NOT_2244( .ZN(II16050), .A(g6065) );
  INV_X1 NOT_2245( .ZN(g8826), .A(II16050) );
  INV_X1 NOT_2246( .ZN(II16053), .A(g6067) );
  INV_X1 NOT_2247( .ZN(g8827), .A(II16053) );
  INV_X1 NOT_2248( .ZN(II16056), .A(g7606) );
  INV_X1 NOT_2249( .ZN(g8828), .A(II16056) );
  INV_X1 NOT_2250( .ZN(II16059), .A(g3878) );
  INV_X1 NOT_2251( .ZN(g8829), .A(II16059) );
  INV_X1 NOT_2252( .ZN(II16062), .A(g3900) );
  INV_X1 NOT_2253( .ZN(g8832), .A(II16062) );
  INV_X1 NOT_2254( .ZN(II16065), .A(g7936) );
  INV_X1 NOT_2255( .ZN(g8835), .A(II16065) );
  INV_X1 NOT_2256( .ZN(II16068), .A(g5438) );
  INV_X1 NOT_2257( .ZN(g8836), .A(II16068) );
  INV_X1 NOT_2258( .ZN(II16071), .A(g5395) );
  INV_X1 NOT_2259( .ZN(g8839), .A(II16071) );
  INV_X1 NOT_2260( .ZN(II16074), .A(g5399) );
  INV_X1 NOT_2261( .ZN(g8840), .A(II16074) );
  INV_X1 NOT_2262( .ZN(II16079), .A(g6086) );
  INV_X1 NOT_2263( .ZN(g8843), .A(II16079) );
  INV_X1 NOT_2264( .ZN(II16082), .A(g5401) );
  INV_X1 NOT_2265( .ZN(g8844), .A(II16082) );
  INV_X1 NOT_2266( .ZN(II16085), .A(g6080) );
  INV_X1 NOT_2267( .ZN(g8845), .A(II16085) );
  INV_X1 NOT_2268( .ZN(g8846), .A(g4779) );
  INV_X1 NOT_2269( .ZN(II16089), .A(g6751) );
  INV_X1 NOT_2270( .ZN(g8847), .A(II16089) );
  INV_X1 NOT_2271( .ZN(II16092), .A(g5402) );
  INV_X1 NOT_2272( .ZN(g8850), .A(II16092) );
  INV_X1 NOT_2273( .ZN(II16095), .A(g6082) );
  INV_X1 NOT_2274( .ZN(g8851), .A(II16095) );
  INV_X1 NOT_2275( .ZN(II16098), .A(g6084) );
  INV_X1 NOT_2276( .ZN(g8852), .A(II16098) );
  INV_X1 NOT_2277( .ZN(II16101), .A(g3878) );
  INV_X1 NOT_2278( .ZN(g8853), .A(II16101) );
  INV_X1 NOT_2279( .ZN(II16104), .A(g6448) );
  INV_X1 NOT_2280( .ZN(g8856), .A(II16104) );
  INV_X1 NOT_2281( .ZN(II16107), .A(g5398) );
  INV_X1 NOT_2282( .ZN(g8859), .A(II16107) );
  INV_X1 NOT_2283( .ZN(II16110), .A(g5404) );
  INV_X1 NOT_2284( .ZN(g8860), .A(II16110) );
  INV_X1 NOT_2285( .ZN(II16114), .A(g7936) );
  INV_X1 NOT_2286( .ZN(g8862), .A(II16114) );
  INV_X1 NOT_2287( .ZN(II16117), .A(g5473) );
  INV_X1 NOT_2288( .ZN(g8863), .A(II16117) );
  INV_X1 NOT_2289( .ZN(II16120), .A(g5400) );
  INV_X1 NOT_2290( .ZN(g8866), .A(II16120) );
  INV_X1 NOT_2291( .ZN(II16123), .A(g5406) );
  INV_X1 NOT_2292( .ZN(g8867), .A(II16123) );
  INV_X1 NOT_2293( .ZN(II16128), .A(g6103) );
  INV_X1 NOT_2294( .ZN(g8870), .A(II16128) );
  INV_X1 NOT_2295( .ZN(II16131), .A(g5408) );
  INV_X1 NOT_2296( .ZN(g8871), .A(II16131) );
  INV_X1 NOT_2297( .ZN(II16134), .A(g6099) );
  INV_X1 NOT_2298( .ZN(g8872), .A(II16134) );
  INV_X1 NOT_2299( .ZN(g8873), .A(g4955) );
  INV_X1 NOT_2300( .ZN(II16138), .A(g7053) );
  INV_X1 NOT_2301( .ZN(g8874), .A(II16138) );
  INV_X1 NOT_2302( .ZN(II16141), .A(g5409) );
  INV_X1 NOT_2303( .ZN(g8877), .A(II16141) );
  INV_X1 NOT_2304( .ZN(II16144), .A(g6101) );
  INV_X1 NOT_2305( .ZN(g8878), .A(II16144) );
  INV_X1 NOT_2306( .ZN(II16147), .A(g3878) );
  INV_X1 NOT_2307( .ZN(g8879), .A(II16147) );
  INV_X1 NOT_2308( .ZN(II16150), .A(g3900) );
  INV_X1 NOT_2309( .ZN(g8882), .A(II16150) );
  INV_X1 NOT_2310( .ZN(II16153), .A(g3306) );
  INV_X1 NOT_2311( .ZN(g8885), .A(II16153) );
  INV_X1 NOT_2312( .ZN(II16156), .A(g5438) );
  INV_X1 NOT_2313( .ZN(g8888), .A(II16156) );
  INV_X1 NOT_2314( .ZN(II16159), .A(g5403) );
  INV_X1 NOT_2315( .ZN(g8891), .A(II16159) );
  INV_X1 NOT_2316( .ZN(II16163), .A(g6031) );
  INV_X1 NOT_2317( .ZN(g8893), .A(II16163) );
  INV_X1 NOT_2318( .ZN(II16166), .A(g6713) );
  INV_X1 NOT_2319( .ZN(g8894), .A(II16166) );
  INV_X1 NOT_2320( .ZN(II16169), .A(g5405) );
  INV_X1 NOT_2321( .ZN(g8897), .A(II16169) );
  INV_X1 NOT_2322( .ZN(II16172), .A(g5413) );
  INV_X1 NOT_2323( .ZN(g8898), .A(II16172) );
  INV_X1 NOT_2324( .ZN(II16176), .A(g7936) );
  INV_X1 NOT_2325( .ZN(g8900), .A(II16176) );
  INV_X1 NOT_2326( .ZN(II16179), .A(g5512) );
  INV_X1 NOT_2327( .ZN(g8901), .A(II16179) );
  INV_X1 NOT_2328( .ZN(II16182), .A(g5407) );
  INV_X1 NOT_2329( .ZN(g8904), .A(II16182) );
  INV_X1 NOT_2330( .ZN(II16185), .A(g5415) );
  INV_X1 NOT_2331( .ZN(g8905), .A(II16185) );
  INV_X1 NOT_2332( .ZN(II16190), .A(g6118) );
  INV_X1 NOT_2333( .ZN(g8908), .A(II16190) );
  INV_X1 NOT_2334( .ZN(II16193), .A(g5417) );
  INV_X1 NOT_2335( .ZN(g8909), .A(II16193) );
  INV_X1 NOT_2336( .ZN(II16196), .A(g6116) );
  INV_X1 NOT_2337( .ZN(g8910), .A(II16196) );
  INV_X1 NOT_2338( .ZN(g8911), .A(g5114) );
  INV_X1 NOT_2339( .ZN(II16200), .A(g7303) );
  INV_X1 NOT_2340( .ZN(g8912), .A(II16200) );
  INV_X1 NOT_2341( .ZN(II16203), .A(g3878) );
  INV_X1 NOT_2342( .ZN(g8915), .A(II16203) );
  INV_X1 NOT_2343( .ZN(II16206), .A(g6448) );
  INV_X1 NOT_2344( .ZN(g8918), .A(II16206) );
  INV_X1 NOT_2345( .ZN(II16209), .A(g5438) );
  INV_X1 NOT_2346( .ZN(g8921), .A(II16209) );
  INV_X1 NOT_2347( .ZN(II16212), .A(g5411) );
  INV_X1 NOT_2348( .ZN(g8924), .A(II16212) );
  INV_X1 NOT_2349( .ZN(II16215), .A(g3462) );
  INV_X1 NOT_2350( .ZN(g8925), .A(II16215) );
  INV_X1 NOT_2351( .ZN(II16218), .A(g5473) );
  INV_X1 NOT_2352( .ZN(g8928), .A(II16218) );
  INV_X1 NOT_2353( .ZN(II16221), .A(g5412) );
  INV_X1 NOT_2354( .ZN(g8931), .A(II16221) );
  INV_X1 NOT_2355( .ZN(II16225), .A(g6042) );
  INV_X1 NOT_2356( .ZN(g8933), .A(II16225) );
  INV_X1 NOT_2357( .ZN(II16228), .A(g7015) );
  INV_X1 NOT_2358( .ZN(g8934), .A(II16228) );
  INV_X1 NOT_2359( .ZN(II16231), .A(g5414) );
  INV_X1 NOT_2360( .ZN(g8937), .A(II16231) );
  INV_X1 NOT_2361( .ZN(II16234), .A(g5420) );
  INV_X1 NOT_2362( .ZN(g8938), .A(II16234) );
  INV_X1 NOT_2363( .ZN(II16238), .A(g7936) );
  INV_X1 NOT_2364( .ZN(g8940), .A(II16238) );
  INV_X1 NOT_2365( .ZN(II16241), .A(g5556) );
  INV_X1 NOT_2366( .ZN(g8941), .A(II16241) );
  INV_X1 NOT_2367( .ZN(II16244), .A(g5416) );
  INV_X1 NOT_2368( .ZN(g8944), .A(II16244) );
  INV_X1 NOT_2369( .ZN(II16247), .A(g5422) );
  INV_X1 NOT_2370( .ZN(g8945), .A(II16247) );
  INV_X1 NOT_2371( .ZN(II16252), .A(g6134) );
  INV_X1 NOT_2372( .ZN(g8948), .A(II16252) );
  INV_X1 NOT_2373( .ZN(II16255), .A(g3900) );
  INV_X1 NOT_2374( .ZN(g8949), .A(II16255) );
  INV_X1 NOT_2375( .ZN(II16258), .A(g3306) );
  INV_X1 NOT_2376( .ZN(g8952), .A(II16258) );
  INV_X1 NOT_2377( .ZN(II16261), .A(g6448) );
  INV_X1 NOT_2378( .ZN(g8955), .A(II16261) );
  INV_X1 NOT_2379( .ZN(II16264), .A(g6713) );
  INV_X1 NOT_2380( .ZN(g8958), .A(II16264) );
  INV_X1 NOT_2381( .ZN(II16267), .A(g5473) );
  INV_X1 NOT_2382( .ZN(g8961), .A(II16267) );
  INV_X1 NOT_2383( .ZN(II16270), .A(g5418) );
  INV_X1 NOT_2384( .ZN(g8964), .A(II16270) );
  INV_X1 NOT_2385( .ZN(II16273), .A(g3618) );
  INV_X1 NOT_2386( .ZN(g8965), .A(II16273) );
  INV_X1 NOT_2387( .ZN(II16276), .A(g5512) );
  INV_X1 NOT_2388( .ZN(g8968), .A(II16276) );
  INV_X1 NOT_2389( .ZN(II16279), .A(g5419) );
  INV_X1 NOT_2390( .ZN(g8971), .A(II16279) );
  INV_X1 NOT_2391( .ZN(II16283), .A(g6046) );
  INV_X1 NOT_2392( .ZN(g8973), .A(II16283) );
  INV_X1 NOT_2393( .ZN(II16286), .A(g7265) );
  INV_X1 NOT_2394( .ZN(g8974), .A(II16286) );
  INV_X1 NOT_2395( .ZN(II16289), .A(g5421) );
  INV_X1 NOT_2396( .ZN(g8977), .A(II16289) );
  INV_X1 NOT_2397( .ZN(II16292), .A(g5426) );
  INV_X32 NOT_2398( .ZN(g8978), .A(II16292) );
  INV_X32 NOT_2399( .ZN(II16296), .A(g3306) );
  INV_X1 NOT_2400( .ZN(g8980), .A(II16296) );
  INV_X1 NOT_2401( .ZN(g8983), .A(g6486) );
  INV_X1 NOT_2402( .ZN(II16300), .A(g3462) );
  INV_X1 NOT_2403( .ZN(g8984), .A(II16300) );
  INV_X1 NOT_2404( .ZN(II16303), .A(g6713) );
  INV_X1 NOT_2405( .ZN(g8987), .A(II16303) );
  INV_X1 NOT_2406( .ZN(II16306), .A(g7015) );
  INV_X1 NOT_2407( .ZN(g8990), .A(II16306) );
  INV_X1 NOT_2408( .ZN(II16309), .A(g5512) );
  INV_X1 NOT_2409( .ZN(g8993), .A(II16309) );
  INV_X1 NOT_2410( .ZN(II16312), .A(g5424) );
  INV_X1 NOT_2411( .ZN(g8996), .A(II16312) );
  INV_X1 NOT_2412( .ZN(II16315), .A(g3774) );
  INV_X1 NOT_2413( .ZN(g8997), .A(II16315) );
  INV_X1 NOT_2414( .ZN(II16318), .A(g5556) );
  INV_X1 NOT_2415( .ZN(g9000), .A(II16318) );
  INV_X1 NOT_2416( .ZN(II16321), .A(g5425) );
  INV_X1 NOT_2417( .ZN(g9003), .A(II16321) );
  INV_X1 NOT_2418( .ZN(II16325), .A(g6052) );
  INV_X1 NOT_2419( .ZN(g9005), .A(II16325) );
  INV_X1 NOT_2420( .ZN(II16328), .A(g3900) );
  INV_X1 NOT_2421( .ZN(g9006), .A(II16328) );
  INV_X1 NOT_2422( .ZN(II16332), .A(g3462) );
  INV_X1 NOT_2423( .ZN(g9010), .A(II16332) );
  INV_X1 NOT_2424( .ZN(II16335), .A(g3618) );
  INV_X1 NOT_2425( .ZN(g9013), .A(II16335) );
  INV_X1 NOT_2426( .ZN(II16338), .A(g7015) );
  INV_X1 NOT_2427( .ZN(g9016), .A(II16338) );
  INV_X1 NOT_2428( .ZN(II16341), .A(g7265) );
  INV_X1 NOT_2429( .ZN(g9019), .A(II16341) );
  INV_X1 NOT_2430( .ZN(II16344), .A(g5556) );
  INV_X1 NOT_2431( .ZN(g9022), .A(II16344) );
  INV_X1 NOT_2432( .ZN(II16347), .A(g5427) );
  INV_X1 NOT_2433( .ZN(g9025), .A(II16347) );
  INV_X1 NOT_2434( .ZN(g9027), .A(g5679) );
  INV_X1 NOT_2435( .ZN(II16354), .A(g3618) );
  INV_X1 NOT_2436( .ZN(g9035), .A(II16354) );
  INV_X1 NOT_2437( .ZN(II16357), .A(g3774) );
  INV_X1 NOT_2438( .ZN(g9038), .A(II16357) );
  INV_X1 NOT_2439( .ZN(II16360), .A(g7265) );
  INV_X1 NOT_2440( .ZN(g9041), .A(II16360) );
  INV_X1 NOT_2441( .ZN(II16363), .A(g3900) );
  INV_X1 NOT_2442( .ZN(g9044), .A(II16363) );
  INV_X1 NOT_2443( .ZN(g9050), .A(g5731) );
  INV_X1 NOT_2444( .ZN(II16372), .A(g3774) );
  INV_X1 NOT_2445( .ZN(g9058), .A(II16372) );
  INV_X1 NOT_2446( .ZN(g9067), .A(g5789) );
  INV_X1 NOT_2447( .ZN(g9084), .A(g5848) );
  INV_X1 NOT_2448( .ZN(II16432), .A(g3366) );
  INV_X1 NOT_2449( .ZN(g9128), .A(II16432) );
  INV_X1 NOT_2450( .ZN(II16438), .A(g3522) );
  INV_X1 NOT_2451( .ZN(g9134), .A(II16438) );
  INV_X1 NOT_2452( .ZN(II16444), .A(g3678) );
  INV_X1 NOT_2453( .ZN(g9140), .A(II16444) );
  INV_X1 NOT_2454( .ZN(II16450), .A(g3834) );
  INV_X1 NOT_2455( .ZN(g9146), .A(II16450) );
  INV_X1 NOT_2456( .ZN(II16453), .A(g7936) );
  INV_X1 NOT_2457( .ZN(g9149), .A(II16453) );
  INV_X1 NOT_2458( .ZN(g9150), .A(g5893) );
  INV_X1 NOT_2459( .ZN(II16457), .A(g7936) );
  INV_X1 NOT_2460( .ZN(g9159), .A(II16457) );
  INV_X1 NOT_2461( .ZN(g9160), .A(g6170) );
  INV_X1 NOT_2462( .ZN(g9161), .A(g5852) );
  INV_X1 NOT_2463( .ZN(II16462), .A(g5438) );
  INV_X1 NOT_2464( .ZN(g9170), .A(II16462) );
  INV_X1 NOT_2465( .ZN(II16465), .A(g6000) );
  INV_X1 NOT_2466( .ZN(g9173), .A(II16465) );
  INV_X1 NOT_2467( .ZN(g9174), .A(g5932) );
  INV_X1 NOT_2468( .ZN(II16469), .A(g7936) );
  INV_X1 NOT_2469( .ZN(g9183), .A(II16469) );
  INV_X1 NOT_2470( .ZN(II16472), .A(g7901) );
  INV_X1 NOT_2471( .ZN(g9184), .A(II16472) );
  INV_X1 NOT_2472( .ZN(g9187), .A(g5803) );
  INV_X1 NOT_2473( .ZN(II16476), .A(g6448) );
  INV_X1 NOT_2474( .ZN(g9196), .A(II16476) );
  INV_X1 NOT_2475( .ZN(II16479), .A(g5438) );
  INV_X1 NOT_2476( .ZN(g9199), .A(II16479) );
  INV_X1 NOT_2477( .ZN(II16482), .A(g6000) );
  INV_X1 NOT_2478( .ZN(g9202), .A(II16482) );
  INV_X1 NOT_2479( .ZN(g9203), .A(g5899) );
  INV_X1 NOT_2480( .ZN(II16486), .A(g5473) );
  INV_X1 NOT_2481( .ZN(g9212), .A(II16486) );
  INV_X1 NOT_2482( .ZN(II16489), .A(g6000) );
  INV_X1 NOT_2483( .ZN(g9215), .A(II16489) );
  INV_X1 NOT_2484( .ZN(g9216), .A(g5966) );
  INV_X1 NOT_2485( .ZN(II16493), .A(g7936) );
  INV_X1 NOT_2486( .ZN(g9225), .A(II16493) );
  INV_X1 NOT_2487( .ZN(g9226), .A(g5434) );
  INV_X1 NOT_2488( .ZN(g9227), .A(g5587) );
  INV_X1 NOT_2489( .ZN(g9228), .A(g7667) );
  INV_X1 NOT_2490( .ZN(II16499), .A(g7901) );
  INV_X1 NOT_2491( .ZN(g9229), .A(II16499) );
  INV_X1 NOT_2492( .ZN(g9232), .A(g5752) );
  INV_X1 NOT_2493( .ZN(II16504), .A(g3306) );
  INV_X1 NOT_2494( .ZN(g9242), .A(II16504) );
  INV_X1 NOT_2495( .ZN(II16507), .A(g6448) );
  INV_X1 NOT_2496( .ZN(g9245), .A(II16507) );
  INV_X1 NOT_2497( .ZN(g9248), .A(g5859) );
  INV_X1 NOT_2498( .ZN(II16511), .A(g6713) );
  INV_X1 NOT_2499( .ZN(g9257), .A(II16511) );
  INV_X1 NOT_2500( .ZN(II16514), .A(g5473) );
  INV_X1 NOT_2501( .ZN(g9260), .A(II16514) );
  INV_X1 NOT_2502( .ZN(II16517), .A(g6000) );
  INV_X1 NOT_2503( .ZN(g9263), .A(II16517) );
  INV_X1 NOT_2504( .ZN(g9264), .A(g5938) );
  INV_X1 NOT_2505( .ZN(II16521), .A(g5512) );
  INV_X1 NOT_2506( .ZN(g9273), .A(II16521) );
  INV_X1 NOT_2507( .ZN(II16524), .A(g6000) );
  INV_X1 NOT_2508( .ZN(g9276), .A(II16524) );
  INV_X1 NOT_2509( .ZN(g9277), .A(g5995) );
  INV_X1 NOT_2510( .ZN(g9286), .A(g6197) );
  INV_X1 NOT_2511( .ZN(g9287), .A(g6638) );
  INV_X1 NOT_2512( .ZN(g9288), .A(g5363) );
  INV_X1 NOT_2513( .ZN(g9289), .A(g5379) );
  INV_X1 NOT_2514( .ZN(II16532), .A(g7901) );
  INV_X1 NOT_2515( .ZN(g9290), .A(II16532) );
  INV_X1 NOT_2516( .ZN(g9293), .A(g5703) );
  INV_X1 NOT_2517( .ZN(II16538), .A(g3306) );
  INV_X1 NOT_2518( .ZN(g9303), .A(II16538) );
  INV_X1 NOT_2519( .ZN(II16541), .A(g5438) );
  INV_X1 NOT_2520( .ZN(g9306), .A(II16541) );
  INV_X1 NOT_2521( .ZN(II16544), .A(g6054) );
  INV_X1 NOT_2522( .ZN(g9309), .A(II16544) );
  INV_X1 NOT_2523( .ZN(g9310), .A(g5811) );
  INV_X1 NOT_2524( .ZN(II16549), .A(g3462) );
  INV_X1 NOT_2525( .ZN(g9320), .A(II16549) );
  INV_X1 NOT_2526( .ZN(II16552), .A(g6713) );
  INV_X32 NOT_2527( .ZN(g9323), .A(II16552) );
  INV_X32 NOT_2528( .ZN(g9326), .A(g5906) );
  INV_X1 NOT_2529( .ZN(II16556), .A(g7015) );
  INV_X1 NOT_2530( .ZN(g9335), .A(II16556) );
  INV_X1 NOT_2531( .ZN(II16559), .A(g5512) );
  INV_X1 NOT_2532( .ZN(g9338), .A(II16559) );
  INV_X1 NOT_2533( .ZN(II16562), .A(g6000) );
  INV_X1 NOT_2534( .ZN(g9341), .A(II16562) );
  INV_X1 NOT_2535( .ZN(g9342), .A(g5972) );
  INV_X1 NOT_2536( .ZN(II16566), .A(g5556) );
  INV_X1 NOT_2537( .ZN(g9351), .A(II16566) );
  INV_X1 NOT_2538( .ZN(II16569), .A(g6000) );
  INV_X1 NOT_2539( .ZN(g9354), .A(II16569) );
  INV_X1 NOT_2540( .ZN(g9355), .A(g7639) );
  INV_X1 NOT_2541( .ZN(g9356), .A(g5665) );
  INV_X1 NOT_2542( .ZN(II16578), .A(g6448) );
  INV_X1 NOT_2543( .ZN(g9368), .A(II16578) );
  INV_X1 NOT_2544( .ZN(II16581), .A(g5438) );
  INV_X1 NOT_2545( .ZN(g9371), .A(II16581) );
  INV_X1 NOT_2546( .ZN(g9374), .A(g5761) );
  INV_X1 NOT_2547( .ZN(II16587), .A(g3462) );
  INV_X1 NOT_2548( .ZN(g9384), .A(II16587) );
  INV_X1 NOT_2549( .ZN(II16590), .A(g5473) );
  INV_X1 NOT_2550( .ZN(g9387), .A(II16590) );
  INV_X1 NOT_2551( .ZN(II16593), .A(g6059) );
  INV_X1 NOT_2552( .ZN(g9390), .A(II16593) );
  INV_X1 NOT_2553( .ZN(g9391), .A(g5867) );
  INV_X1 NOT_2554( .ZN(II16598), .A(g3618) );
  INV_X1 NOT_2555( .ZN(g9401), .A(II16598) );
  INV_X1 NOT_2556( .ZN(II16601), .A(g7015) );
  INV_X1 NOT_2557( .ZN(g9404), .A(II16601) );
  INV_X1 NOT_2558( .ZN(g9407), .A(g5945) );
  INV_X1 NOT_2559( .ZN(II16605), .A(g7265) );
  INV_X1 NOT_2560( .ZN(g9416), .A(II16605) );
  INV_X1 NOT_2561( .ZN(II16608), .A(g5556) );
  INV_X1 NOT_2562( .ZN(g9419), .A(II16608) );
  INV_X1 NOT_2563( .ZN(II16611), .A(g6000) );
  INV_X1 NOT_2564( .ZN(g9422), .A(II16611) );
  INV_X1 NOT_2565( .ZN(g9423), .A(g5428) );
  INV_X1 NOT_2566( .ZN(g9424), .A(g5469) );
  INV_X1 NOT_2567( .ZN(g9425), .A(g5346) );
  INV_X1 NOT_2568( .ZN(g9426), .A(g5543) );
  INV_X1 NOT_2569( .ZN(g9427), .A(g5645) );
  INV_X1 NOT_2570( .ZN(II16624), .A(g3306) );
  INV_X1 NOT_2571( .ZN(g9443), .A(II16624) );
  INV_X1 NOT_2572( .ZN(II16627), .A(g6448) );
  INV_X1 NOT_2573( .ZN(g9446), .A(II16627) );
  INV_X1 NOT_2574( .ZN(II16630), .A(g6057) );
  INV_X1 NOT_2575( .ZN(g9449), .A(II16630) );
  INV_X1 NOT_2576( .ZN(II16633), .A(g6486) );
  INV_X1 NOT_2577( .ZN(g9450), .A(II16633) );
  INV_X1 NOT_2578( .ZN(g9453), .A(g5717) );
  INV_X1 NOT_2579( .ZN(II16641), .A(g6713) );
  INV_X1 NOT_2580( .ZN(g9465), .A(II16641) );
  INV_X1 NOT_2581( .ZN(II16644), .A(g5473) );
  INV_X1 NOT_2582( .ZN(g9468), .A(II16644) );
  INV_X1 NOT_2583( .ZN(g9471), .A(g5820) );
  INV_X1 NOT_2584( .ZN(II16650), .A(g3618) );
  INV_X1 NOT_2585( .ZN(g9481), .A(II16650) );
  INV_X1 NOT_2586( .ZN(II16653), .A(g5512) );
  INV_X1 NOT_2587( .ZN(g9484), .A(II16653) );
  INV_X1 NOT_2588( .ZN(II16656), .A(g6066) );
  INV_X1 NOT_2589( .ZN(g9487), .A(II16656) );
  INV_X1 NOT_2590( .ZN(g9488), .A(g5914) );
  INV_X1 NOT_2591( .ZN(II16661), .A(g3774) );
  INV_X1 NOT_2592( .ZN(g9498), .A(II16661) );
  INV_X1 NOT_2593( .ZN(II16664), .A(g7265) );
  INV_X1 NOT_2594( .ZN(g9501), .A(II16664) );
  INV_X1 NOT_2595( .ZN(g9504), .A(g6149) );
  INV_X1 NOT_2596( .ZN(g9505), .A(g6227) );
  INV_X1 NOT_2597( .ZN(g9506), .A(g6444) );
  INV_X1 NOT_2598( .ZN(g9507), .A(g5953) );
  INV_X1 NOT_2599( .ZN(II16677), .A(g3306) );
  INV_X1 NOT_2600( .ZN(g9524), .A(II16677) );
  INV_X1 NOT_2601( .ZN(g9527), .A(g5508) );
  INV_X1 NOT_2602( .ZN(II16681), .A(g6643) );
  INV_X1 NOT_2603( .ZN(g9528), .A(II16681) );
  INV_X1 NOT_2604( .ZN(II16684), .A(g6486) );
  INV_X1 NOT_2605( .ZN(g9531), .A(II16684) );
  INV_X1 NOT_2606( .ZN(g9569), .A(g5683) );
  INV_X1 NOT_2607( .ZN(II16694), .A(g3462) );
  INV_X1 NOT_2608( .ZN(g9585), .A(II16694) );
  INV_X1 NOT_2609( .ZN(II16697), .A(g6713) );
  INV_X1 NOT_2610( .ZN(g9588), .A(II16697) );
  INV_X1 NOT_2611( .ZN(II16700), .A(g6064) );
  INV_X1 NOT_2612( .ZN(g9591), .A(II16700) );
  INV_X1 NOT_2613( .ZN(II16703), .A(g6751) );
  INV_X1 NOT_2614( .ZN(g9592), .A(II16703) );
  INV_X1 NOT_2615( .ZN(g9595), .A(g5775) );
  INV_X1 NOT_2616( .ZN(II16711), .A(g7015) );
  INV_X1 NOT_2617( .ZN(g9607), .A(II16711) );
  INV_X1 NOT_2618( .ZN(II16714), .A(g5512) );
  INV_X1 NOT_2619( .ZN(g9610), .A(II16714) );
  INV_X1 NOT_2620( .ZN(g9613), .A(g5876) );
  INV_X1 NOT_2621( .ZN(II16720), .A(g3774) );
  INV_X1 NOT_2622( .ZN(g9623), .A(II16720) );
  INV_X1 NOT_2623( .ZN(II16723), .A(g5556) );
  INV_X1 NOT_2624( .ZN(g9626), .A(II16723) );
  INV_X1 NOT_2625( .ZN(II16726), .A(g6085) );
  INV_X1 NOT_2626( .ZN(g9629), .A(II16726) );
  INV_X1 NOT_2627( .ZN(II16741), .A(g6062) );
  INV_X1 NOT_2628( .ZN(g9640), .A(II16741) );
  INV_X1 NOT_2629( .ZN(II16744), .A(g3338) );
  INV_X1 NOT_2630( .ZN(g9641), .A(II16744) );
  INV_X1 NOT_2631( .ZN(II16747), .A(g6643) );
  INV_X1 NOT_2632( .ZN(g9644), .A(II16747) );
  INV_X1 NOT_2633( .ZN(g9649), .A(g5982) );
  INV_X1 NOT_2634( .ZN(II16759), .A(g3462) );
  INV_X1 NOT_2635( .ZN(g9666), .A(II16759) );
  INV_X1 NOT_2636( .ZN(g9669), .A(g5552) );
  INV_X1 NOT_2637( .ZN(II16763), .A(g6945) );
  INV_X1 NOT_2638( .ZN(g9670), .A(II16763) );
  INV_X1 NOT_2639( .ZN(II16766), .A(g6751) );
  INV_X1 NOT_2640( .ZN(g9673), .A(II16766) );
  INV_X1 NOT_2641( .ZN(g9711), .A(g5735) );
  INV_X1 NOT_2642( .ZN(II16776), .A(g3618) );
  INV_X1 NOT_2643( .ZN(g9727), .A(II16776) );
  INV_X1 NOT_2644( .ZN(II16779), .A(g7015) );
  INV_X1 NOT_2645( .ZN(g9730), .A(II16779) );
  INV_X1 NOT_2646( .ZN(II16782), .A(g6083) );
  INV_X1 NOT_2647( .ZN(g9733), .A(II16782) );
  INV_X1 NOT_2648( .ZN(II16785), .A(g7053) );
  INV_X1 NOT_2649( .ZN(g9734), .A(II16785) );
  INV_X1 NOT_2650( .ZN(g9737), .A(g5834) );
  INV_X1 NOT_2651( .ZN(II16793), .A(g7265) );
  INV_X1 NOT_2652( .ZN(g9749), .A(II16793) );
  INV_X1 NOT_2653( .ZN(II16796), .A(g5556) );
  INV_X1 NOT_2654( .ZN(g9752), .A(II16796) );
  INV_X1 NOT_2655( .ZN(g9755), .A(g5431) );
  INV_X1 NOT_2656( .ZN(g9756), .A(g5504) );
  INV_X1 NOT_2657( .ZN(g9757), .A(g5601) );
  INV_X1 NOT_2658( .ZN(g9758), .A(g5618) );
  INV_X1 NOT_2659( .ZN(II16811), .A(g3338) );
  INV_X1 NOT_2660( .ZN(g9767), .A(II16811) );
  INV_X1 NOT_2661( .ZN(II16814), .A(g6486) );
  INV_X1 NOT_2662( .ZN(g9770), .A(II16814) );
  INV_X1 NOT_2663( .ZN(II16832), .A(g6081) );
  INV_X1 NOT_2664( .ZN(g9786), .A(II16832) );
  INV_X1 NOT_2665( .ZN(II16835), .A(g3494) );
  INV_X1 NOT_2666( .ZN(g9787), .A(II16835) );
  INV_X1 NOT_2667( .ZN(II16838), .A(g6945) );
  INV_X1 NOT_2668( .ZN(g9790), .A(II16838) );
  INV_X1 NOT_2669( .ZN(g9795), .A(g6019) );
  INV_X1 NOT_2670( .ZN(II16850), .A(g3618) );
  INV_X1 NOT_2671( .ZN(g9812), .A(II16850) );
  INV_X1 NOT_2672( .ZN(g9815), .A(g5598) );
  INV_X1 NOT_2673( .ZN(II16854), .A(g7195) );
  INV_X1 NOT_2674( .ZN(g9816), .A(II16854) );
  INV_X1 NOT_2675( .ZN(II16857), .A(g7053) );
  INV_X1 NOT_2676( .ZN(g9819), .A(II16857) );
  INV_X1 NOT_2677( .ZN(g9857), .A(g5793) );
  INV_X1 NOT_2678( .ZN(II16867), .A(g3774) );
  INV_X1 NOT_2679( .ZN(g9873), .A(II16867) );
  INV_X1 NOT_2680( .ZN(II16870), .A(g7265) );
  INV_X1 NOT_2681( .ZN(g9876), .A(II16870) );
  INV_X1 NOT_2682( .ZN(II16873), .A(g6102) );
  INV_X1 NOT_2683( .ZN(g9879), .A(II16873) );
  INV_X1 NOT_2684( .ZN(II16876), .A(g7303) );
  INV_X1 NOT_2685( .ZN(g9880), .A(II16876) );
  INV_X1 NOT_2686( .ZN(g9884), .A(g6310) );
  INV_X1 NOT_2687( .ZN(g9885), .A(g6905) );
  INV_X1 NOT_2688( .ZN(g9886), .A(g7149) );
  INV_X1 NOT_2689( .ZN(II16897), .A(g6643) );
  INV_X1 NOT_2690( .ZN(g9895), .A(II16897) );
  INV_X1 NOT_2691( .ZN(II16900), .A(g6486) );
  INV_X1 NOT_2692( .ZN(g9898), .A(II16900) );
  INV_X1 NOT_2693( .ZN(II16915), .A(g3494) );
  INV_X32 NOT_2694( .ZN(g9913), .A(II16915) );
  INV_X32 NOT_2695( .ZN(II16918), .A(g6751) );
  INV_X1 NOT_2696( .ZN(g9916), .A(II16918) );
  INV_X1 NOT_2697( .ZN(II16936), .A(g6100) );
  INV_X1 NOT_2698( .ZN(g9932), .A(II16936) );
  INV_X1 NOT_2699( .ZN(II16939), .A(g3650) );
  INV_X1 NOT_2700( .ZN(g9933), .A(II16939) );
  INV_X1 NOT_2701( .ZN(II16942), .A(g7195) );
  INV_X1 NOT_2702( .ZN(g9936), .A(II16942) );
  INV_X1 NOT_2703( .ZN(g9941), .A(g6035) );
  INV_X1 NOT_2704( .ZN(II16954), .A(g3774) );
  INV_X1 NOT_2705( .ZN(g9958), .A(II16954) );
  INV_X1 NOT_2706( .ZN(g9961), .A(g5615) );
  INV_X1 NOT_2707( .ZN(II16958), .A(g7391) );
  INV_X1 NOT_2708( .ZN(g9962), .A(II16958) );
  INV_X1 NOT_2709( .ZN(II16961), .A(g7303) );
  INV_X1 NOT_2710( .ZN(g9965), .A(II16961) );
  INV_X1 NOT_2711( .ZN(II16972), .A(g3900) );
  INV_X1 NOT_2712( .ZN(g10004), .A(II16972) );
  INV_X1 NOT_2713( .ZN(g10015), .A(g5292) );
  INV_X1 NOT_2714( .ZN(II16984), .A(g7936) );
  INV_X1 NOT_2715( .ZN(g10016), .A(II16984) );
  INV_X1 NOT_2716( .ZN(II16987), .A(g6079) );
  INV_X1 NOT_2717( .ZN(g10017), .A(II16987) );
  INV_X1 NOT_2718( .ZN(II16990), .A(g3338) );
  INV_X1 NOT_2719( .ZN(g10018), .A(II16990) );
  INV_X1 NOT_2720( .ZN(II16993), .A(g6643) );
  INV_X1 NOT_2721( .ZN(g10021), .A(II16993) );
  INV_X1 NOT_2722( .ZN(II17009), .A(g6945) );
  INV_X1 NOT_2723( .ZN(g10049), .A(II17009) );
  INV_X1 NOT_2724( .ZN(II17012), .A(g6751) );
  INV_X1 NOT_2725( .ZN(g10052), .A(II17012) );
  INV_X1 NOT_2726( .ZN(II17027), .A(g3650) );
  INV_X1 NOT_2727( .ZN(g10067), .A(II17027) );
  INV_X1 NOT_2728( .ZN(II17030), .A(g7053) );
  INV_X1 NOT_2729( .ZN(g10070), .A(II17030) );
  INV_X1 NOT_2730( .ZN(II17048), .A(g6117) );
  INV_X1 NOT_2731( .ZN(g10086), .A(II17048) );
  INV_X1 NOT_2732( .ZN(II17051), .A(g3806) );
  INV_X1 NOT_2733( .ZN(g10087), .A(II17051) );
  INV_X1 NOT_2734( .ZN(II17054), .A(g7391) );
  INV_X1 NOT_2735( .ZN(g10090), .A(II17054) );
  INV_X1 NOT_2736( .ZN(II17066), .A(g3900) );
  INV_X1 NOT_2737( .ZN(g10096), .A(II17066) );
  INV_X1 NOT_2738( .ZN(g10099), .A(g7700) );
  INV_X1 NOT_2739( .ZN(II17070), .A(g7528) );
  INV_X1 NOT_2740( .ZN(g10100), .A(II17070) );
  INV_X1 NOT_2741( .ZN(II17081), .A(g3338) );
  INV_X1 NOT_2742( .ZN(g10109), .A(II17081) );
  INV_X1 NOT_2743( .ZN(g10124), .A(g5326) );
  INV_X1 NOT_2744( .ZN(II17097), .A(g7936) );
  INV_X1 NOT_2745( .ZN(g10125), .A(II17097) );
  INV_X1 NOT_2746( .ZN(II17100), .A(g6098) );
  INV_X1 NOT_2747( .ZN(g10126), .A(II17100) );
  INV_X1 NOT_2748( .ZN(II17103), .A(g3494) );
  INV_X1 NOT_2749( .ZN(g10127), .A(II17103) );
  INV_X1 NOT_2750( .ZN(II17106), .A(g6945) );
  INV_X1 NOT_2751( .ZN(g10130), .A(II17106) );
  INV_X1 NOT_2752( .ZN(II17122), .A(g7195) );
  INV_X1 NOT_2753( .ZN(g10158), .A(II17122) );
  INV_X1 NOT_2754( .ZN(II17125), .A(g7053) );
  INV_X1 NOT_2755( .ZN(g10161), .A(II17125) );
  INV_X1 NOT_2756( .ZN(II17140), .A(g3806) );
  INV_X1 NOT_2757( .ZN(g10176), .A(II17140) );
  INV_X1 NOT_2758( .ZN(II17143), .A(g7303) );
  INV_X1 NOT_2759( .ZN(g10179), .A(II17143) );
  INV_X1 NOT_2760( .ZN(II17159), .A(g3900) );
  INV_X1 NOT_2761( .ZN(g10189), .A(II17159) );
  INV_X1 NOT_2762( .ZN(II17184), .A(g3494) );
  INV_X1 NOT_2763( .ZN(g10214), .A(II17184) );
  INV_X1 NOT_2764( .ZN(g10229), .A(g5349) );
  INV_X1 NOT_2765( .ZN(II17200), .A(g7936) );
  INV_X1 NOT_2766( .ZN(g10230), .A(II17200) );
  INV_X1 NOT_2767( .ZN(II17203), .A(g6115) );
  INV_X1 NOT_2768( .ZN(g10231), .A(II17203) );
  INV_X1 NOT_2769( .ZN(II17206), .A(g3650) );
  INV_X1 NOT_2770( .ZN(g10232), .A(II17206) );
  INV_X1 NOT_2771( .ZN(II17209), .A(g7195) );
  INV_X1 NOT_2772( .ZN(g10235), .A(II17209) );
  INV_X1 NOT_2773( .ZN(II17225), .A(g7391) );
  INV_X1 NOT_2774( .ZN(g10263), .A(II17225) );
  INV_X1 NOT_2775( .ZN(II17228), .A(g7303) );
  INV_X1 NOT_2776( .ZN(g10266), .A(II17228) );
  INV_X1 NOT_2777( .ZN(II17235), .A(g3900) );
  INV_X1 NOT_2778( .ZN(g10273), .A(II17235) );
  INV_X1 NOT_2779( .ZN(II17238), .A(g3900) );
  INV_X1 NOT_2780( .ZN(g10276), .A(II17238) );
  INV_X1 NOT_2781( .ZN(II17278), .A(g3650) );
  INV_X1 NOT_2782( .ZN(g10316), .A(II17278) );
  INV_X1 NOT_2783( .ZN(g10331), .A(g5366) );
  INV_X1 NOT_2784( .ZN(II17294), .A(g7936) );
  INV_X1 NOT_2785( .ZN(g10332), .A(II17294) );
  INV_X1 NOT_2786( .ZN(II17297), .A(g6130) );
  INV_X1 NOT_2787( .ZN(g10333), .A(II17297) );
  INV_X1 NOT_2788( .ZN(II17300), .A(g3806) );
  INV_X1 NOT_2789( .ZN(g10334), .A(II17300) );
  INV_X1 NOT_2790( .ZN(II17303), .A(g7391) );
  INV_X1 NOT_2791( .ZN(g10337), .A(II17303) );
  INV_X1 NOT_2792( .ZN(II17311), .A(g3900) );
  INV_X1 NOT_2793( .ZN(g10357), .A(II17311) );
  INV_X1 NOT_2794( .ZN(II17363), .A(g3806) );
  INV_X1 NOT_2795( .ZN(g10409), .A(II17363) );
  INV_X1 NOT_2796( .ZN(II17370), .A(g3900) );
  INV_X1 NOT_2797( .ZN(g10416), .A(II17370) );
  INV_X1 NOT_2798( .ZN(II17373), .A(g3900) );
  INV_X1 NOT_2799( .ZN(g10419), .A(II17373) );
  INV_X1 NOT_2800( .ZN(g10424), .A(g7910) );
  INV_X1 NOT_2801( .ZN(g10481), .A(g7826) );
  INV_X1 NOT_2802( .ZN(II17433), .A(g3900) );
  INV_X1 NOT_2803( .ZN(g10482), .A(II17433) );
  INV_X1 NOT_2804( .ZN(g10486), .A(g7957) );
  INV_X1 NOT_2805( .ZN(g10500), .A(g7962) );
  INV_X1 NOT_2806( .ZN(II17483), .A(g3900) );
  INV_X1 NOT_2807( .ZN(g10542), .A(II17483) );
  INV_X1 NOT_2808( .ZN(II17486), .A(g3900) );
  INV_X1 NOT_2809( .ZN(g10545), .A(II17486) );
  INV_X1 NOT_2810( .ZN(g10549), .A(g7999) );
  INV_X1 NOT_2811( .ZN(g10560), .A(g8008) );
  INV_X1 NOT_2812( .ZN(g10574), .A(g8013) );
  INV_X1 NOT_2813( .ZN(II17527), .A(g3900) );
  INV_X1 NOT_2814( .ZN(g10601), .A(II17527) );
  INV_X1 NOT_2815( .ZN(g10606), .A(g8074) );
  INV_X1 NOT_2816( .ZN(g10617), .A(g8083) );
  INV_X1 NOT_2817( .ZN(g10631), .A(g8088) );
  INV_X1 NOT_2818( .ZN(II17557), .A(g3900) );
  INV_X1 NOT_2819( .ZN(g10646), .A(II17557) );
  INV_X1 NOT_2820( .ZN(g10653), .A(g8159) );
  INV_X1 NOT_2821( .ZN(g10664), .A(g8168) );
  INV_X1 NOT_2822( .ZN(g10683), .A(g8245) );
  INV_X1 NOT_2823( .ZN(g10694), .A(g4326) );
  INV_X1 NOT_2824( .ZN(g10714), .A(g4495) );
  INV_X1 NOT_2825( .ZN(g10730), .A(g6173) );
  INV_X1 NOT_2826( .ZN(g10735), .A(g4671) );
  INV_X1 NOT_2827( .ZN(g10749), .A(g6205) );
  INV_X1 NOT_2828( .ZN(g10754), .A(g4848) );
  INV_X1 NOT_2829( .ZN(g10765), .A(g6048) );
  INV_X1 NOT_2830( .ZN(g10766), .A(g6676) );
  INV_X1 NOT_2831( .ZN(g10767), .A(g6294) );
  INV_X1 NOT_2832( .ZN(g10772), .A(g6978) );
  INV_X1 NOT_2833( .ZN(g10773), .A(g6431) );
  INV_X1 NOT_2834( .ZN(II17627), .A(g7575) );
  INV_X1 NOT_2835( .ZN(g10779), .A(II17627) );
  INV_X1 NOT_2836( .ZN(g10783), .A(g7228) );
  INV_X1 NOT_2837( .ZN(II17632), .A(g6183) );
  INV_X1 NOT_2838( .ZN(g10787), .A(II17632) );
  INV_X1 NOT_2839( .ZN(g10788), .A(g7424) );
  INV_X1 NOT_2840( .ZN(II17637), .A(g6204) );
  INV_X1 NOT_2841( .ZN(g10792), .A(II17637) );
  INV_X1 NOT_2842( .ZN(II17641), .A(g6215) );
  INV_X1 NOT_2843( .ZN(g10796), .A(II17641) );
  INV_X1 NOT_2844( .ZN(II17645), .A(g6288) );
  INV_X1 NOT_2845( .ZN(g10800), .A(II17645) );
  INV_X1 NOT_2846( .ZN(II17649), .A(g6293) );
  INV_X1 NOT_2847( .ZN(g10804), .A(II17649) );
  INV_X1 NOT_2848( .ZN(II17653), .A(g6304) );
  INV_X1 NOT_2849( .ZN(g10808), .A(II17653) );
  INV_X1 NOT_2850( .ZN(g10809), .A(g5701) );
  INV_X1 NOT_2851( .ZN(II17658), .A(g6367) );
  INV_X1 NOT_2852( .ZN(g10813), .A(II17658) );
  INV_X1 NOT_2853( .ZN(II17662), .A(g6425) );
  INV_X1 NOT_2854( .ZN(g10817), .A(II17662) );
  INV_X1 NOT_2855( .ZN(II17666), .A(g6430) );
  INV_X1 NOT_2856( .ZN(g10821), .A(II17666) );
  INV_X1 NOT_2857( .ZN(II17670), .A(g6441) );
  INV_X1 NOT_2858( .ZN(g10825), .A(II17670) );
  INV_X1 NOT_2859( .ZN(II17673), .A(g8107) );
  INV_X1 NOT_2860( .ZN(g10826), .A(II17673) );
  INV_X1 NOT_2861( .ZN(g10829), .A(g5749) );
  INV_X1 NOT_2862( .ZN(II17677), .A(g6517) );
  INV_X1 NOT_2863( .ZN(g10830), .A(II17677) );
  INV_X1 NOT_2864( .ZN(II17681), .A(g6572) );
  INV_X1 NOT_2865( .ZN(g10834), .A(II17681) );
  INV_X1 NOT_2866( .ZN(II17685), .A(g6630) );
  INV_X4 NOT_2867( .ZN(g10838), .A(II17685) );
  INV_X4 NOT_2868( .ZN(II17689), .A(g6635) );
  INV_X4 NOT_2869( .ZN(g10842), .A(II17689) );
  INV_X4 NOT_2870( .ZN(II17692), .A(g8107) );
  INV_X1 NOT_2871( .ZN(g10843), .A(II17692) );
  INV_X1 NOT_2872( .ZN(g10846), .A(g5799) );
  INV_X1 NOT_2873( .ZN(g10847), .A(g5800) );
  INV_X1 NOT_2874( .ZN(g10848), .A(g5801) );
  INV_X1 NOT_2875( .ZN(II17698), .A(g6711) );
  INV_X1 NOT_2876( .ZN(g10849), .A(II17698) );
  INV_X1 NOT_2877( .ZN(II17701), .A(g6781) );
  INV_X1 NOT_2878( .ZN(g10850), .A(II17701) );
  INV_X1 NOT_2879( .ZN(II17705), .A(g6836) );
  INV_X1 NOT_2880( .ZN(g10854), .A(II17705) );
  INV_X1 NOT_2881( .ZN(II17709), .A(g6894) );
  INV_X1 NOT_2882( .ZN(g10858), .A(II17709) );
  INV_X1 NOT_2883( .ZN(II17712), .A(g8031) );
  INV_X1 NOT_2884( .ZN(g10859), .A(II17712) );
  INV_X1 NOT_2885( .ZN(II17715), .A(g8107) );
  INV_X1 NOT_2886( .ZN(g10862), .A(II17715) );
  INV_X1 NOT_2887( .ZN(g10865), .A(g6131) );
  INV_X1 NOT_2888( .ZN(g10866), .A(g5849) );
  INV_X1 NOT_2889( .ZN(g10867), .A(g5850) );
  INV_X1 NOT_2890( .ZN(II17721), .A(g6641) );
  INV_X1 NOT_2891( .ZN(g10868), .A(II17721) );
  INV_X1 NOT_2892( .ZN(II17724), .A(g6942) );
  INV_X1 NOT_2893( .ZN(g10869), .A(II17724) );
  INV_X1 NOT_2894( .ZN(II17727), .A(g7013) );
  INV_X1 NOT_2895( .ZN(g10870), .A(II17727) );
  INV_X1 NOT_2896( .ZN(II17730), .A(g7083) );
  INV_X1 NOT_2897( .ZN(g10871), .A(II17730) );
  INV_X1 NOT_2898( .ZN(II17734), .A(g7138) );
  INV_X1 NOT_2899( .ZN(g10875), .A(II17734) );
  INV_X1 NOT_2900( .ZN(II17737), .A(g6000) );
  INV_X1 NOT_2901( .ZN(g10876), .A(II17737) );
  INV_X1 NOT_2902( .ZN(II17740), .A(g8031) );
  INV_X1 NOT_2903( .ZN(g10877), .A(II17740) );
  INV_X1 NOT_2904( .ZN(II17743), .A(g8107) );
  INV_X1 NOT_2905( .ZN(g10880), .A(II17743) );
  INV_X1 NOT_2906( .ZN(II17746), .A(g8107) );
  INV_X1 NOT_2907( .ZN(g10883), .A(II17746) );
  INV_X1 NOT_2908( .ZN(g10886), .A(g5889) );
  INV_X1 NOT_2909( .ZN(II17750), .A(g7157) );
  INV_X1 NOT_2910( .ZN(g10887), .A(II17750) );
  INV_X1 NOT_2911( .ZN(II17753), .A(g6943) );
  INV_X1 NOT_2912( .ZN(g10888), .A(II17753) );
  INV_X1 NOT_2913( .ZN(II17756), .A(g7192) );
  INV_X1 NOT_2914( .ZN(g10889), .A(II17756) );
  INV_X1 NOT_2915( .ZN(II17759), .A(g7263) );
  INV_X1 NOT_2916( .ZN(g10890), .A(II17759) );
  INV_X1 NOT_2917( .ZN(II17762), .A(g7333) );
  INV_X1 NOT_2918( .ZN(g10891), .A(II17762) );
  INV_X1 NOT_2919( .ZN(II17765), .A(g7976) );
  INV_X1 NOT_2920( .ZN(g10892), .A(II17765) );
  INV_X1 NOT_2921( .ZN(II17768), .A(g8031) );
  INV_X1 NOT_2922( .ZN(g10895), .A(II17768) );
  INV_X1 NOT_2923( .ZN(II17771), .A(g8107) );
  INV_X1 NOT_2924( .ZN(g10898), .A(II17771) );
  INV_X1 NOT_2925( .ZN(II17774), .A(g8107) );
  INV_X1 NOT_2926( .ZN(g10901), .A(II17774) );
  INV_X1 NOT_2927( .ZN(g10904), .A(g5922) );
  INV_X1 NOT_2928( .ZN(g10905), .A(g5923) );
  INV_X1 NOT_2929( .ZN(g10906), .A(g5924) );
  INV_X1 NOT_2930( .ZN(II17780), .A(g7348) );
  INV_X1 NOT_2931( .ZN(g10907), .A(II17780) );
  INV_X1 NOT_2932( .ZN(II17783), .A(g7353) );
  INV_X1 NOT_2933( .ZN(g10908), .A(II17783) );
  INV_X1 NOT_2934( .ZN(II17786), .A(g7193) );
  INV_X1 NOT_2935( .ZN(g10909), .A(II17786) );
  INV_X1 NOT_2936( .ZN(II17789), .A(g7388) );
  INV_X1 NOT_2937( .ZN(g10910), .A(II17789) );
  INV_X1 NOT_2938( .ZN(II17792), .A(g7459) );
  INV_X1 NOT_2939( .ZN(g10911), .A(II17792) );
  INV_X1 NOT_2940( .ZN(II17795), .A(g7976) );
  INV_X1 NOT_2941( .ZN(g10912), .A(II17795) );
  INV_X1 NOT_2942( .ZN(II17798), .A(g8031) );
  INV_X1 NOT_2943( .ZN(g10915), .A(II17798) );
  INV_X1 NOT_2944( .ZN(II17801), .A(g8107) );
  INV_X1 NOT_2945( .ZN(g10918), .A(II17801) );
  INV_X1 NOT_2946( .ZN(II17804), .A(g8031) );
  INV_X1 NOT_2947( .ZN(g10921), .A(II17804) );
  INV_X1 NOT_2948( .ZN(II17807), .A(g8107) );
  INV_X1 NOT_2949( .ZN(g10924), .A(II17807) );
  INV_X1 NOT_2950( .ZN(g10927), .A(g6153) );
  INV_X1 NOT_2951( .ZN(g10928), .A(g5951) );
  INV_X1 NOT_2952( .ZN(g10929), .A(g5952) );
  INV_X1 NOT_2953( .ZN(II17813), .A(g5707) );
  INV_X1 NOT_2954( .ZN(g10930), .A(II17813) );
  INV_X1 NOT_2955( .ZN(II17816), .A(g7346) );
  INV_X1 NOT_2956( .ZN(g10931), .A(II17816) );
  INV_X1 NOT_2957( .ZN(II17819), .A(g6448) );
  INV_X1 NOT_2958( .ZN(g10932), .A(II17819) );
  INV_X1 NOT_2959( .ZN(II17822), .A(g7478) );
  INV_X1 NOT_2960( .ZN(g10933), .A(II17822) );
  INV_X1 NOT_2961( .ZN(II17825), .A(g7483) );
  INV_X1 NOT_2962( .ZN(g10934), .A(II17825) );
  INV_X1 NOT_2963( .ZN(II17828), .A(g7389) );
  INV_X1 NOT_2964( .ZN(g10935), .A(II17828) );
  INV_X1 NOT_2965( .ZN(II17831), .A(g7518) );
  INV_X1 NOT_2966( .ZN(g10936), .A(II17831) );
  INV_X1 NOT_2967( .ZN(II17834), .A(g7976) );
  INV_X1 NOT_2968( .ZN(g10937), .A(II17834) );
  INV_X1 NOT_2969( .ZN(II17837), .A(g8031) );
  INV_X1 NOT_2970( .ZN(g10940), .A(II17837) );
  INV_X1 NOT_2971( .ZN(II17840), .A(g8107) );
  INV_X1 NOT_2972( .ZN(g10943), .A(II17840) );
  INV_X1 NOT_2973( .ZN(II17843), .A(g8031) );
  INV_X1 NOT_2974( .ZN(g10946), .A(II17843) );
  INV_X1 NOT_2975( .ZN(II17846), .A(g8107) );
  INV_X1 NOT_2976( .ZN(g10949), .A(II17846) );
  INV_X1 NOT_2977( .ZN(II17849), .A(g8103) );
  INV_X1 NOT_2978( .ZN(g10952), .A(II17849) );
  INV_X1 NOT_2979( .ZN(g10961), .A(g5978) );
  INV_X1 NOT_2980( .ZN(g10962), .A(g5979) );
  INV_X1 NOT_2981( .ZN(II17854), .A(g6232) );
  INV_X1 NOT_2982( .ZN(g10963), .A(II17854) );
  INV_X1 NOT_2983( .ZN(II17857), .A(g6448) );
  INV_X1 NOT_2984( .ZN(g10966), .A(II17857) );
  INV_X1 NOT_2985( .ZN(II17860), .A(g5765) );
  INV_X1 NOT_2986( .ZN(g10967), .A(II17860) );
  INV_X1 NOT_2987( .ZN(II17863), .A(g7476) );
  INV_X1 NOT_2988( .ZN(g10968), .A(II17863) );
  INV_X1 NOT_2989( .ZN(II17866), .A(g6713) );
  INV_X1 NOT_2990( .ZN(g10969), .A(II17866) );
  INV_X1 NOT_2991( .ZN(II17869), .A(g7534) );
  INV_X1 NOT_2992( .ZN(g10972), .A(II17869) );
  INV_X1 NOT_2993( .ZN(II17872), .A(g7539) );
  INV_X1 NOT_2994( .ZN(g10973), .A(II17872) );
  INV_X1 NOT_2995( .ZN(II17875), .A(g7976) );
  INV_X1 NOT_2996( .ZN(g10974), .A(II17875) );
  INV_X1 NOT_2997( .ZN(II17878), .A(g8031) );
  INV_X1 NOT_2998( .ZN(g10977), .A(II17878) );
  INV_X1 NOT_2999( .ZN(II17881), .A(g7976) );
  INV_X1 NOT_3000( .ZN(g10980), .A(II17881) );
  INV_X1 NOT_3001( .ZN(II17884), .A(g8031) );
  INV_X1 NOT_3002( .ZN(g10983), .A(II17884) );
  INV_X1 NOT_3003( .ZN(g10986), .A(g6014) );
  INV_X1 NOT_3004( .ZN(g10987), .A(g6015) );
  INV_X1 NOT_3005( .ZN(II17889), .A(g6314) );
  INV_X1 NOT_3006( .ZN(g10988), .A(II17889) );
  INV_X1 NOT_3007( .ZN(II17892), .A(g6232) );
  INV_X1 NOT_3008( .ZN(g10991), .A(II17892) );
  INV_X1 NOT_3009( .ZN(II17895), .A(g6448) );
  INV_X1 NOT_3010( .ZN(g10994), .A(II17895) );
  INV_X1 NOT_3011( .ZN(II17898), .A(g6643) );
  INV_X1 NOT_3012( .ZN(g10995), .A(II17898) );
  INV_X1 NOT_3013( .ZN(II17901), .A(g6369) );
  INV_X1 NOT_3014( .ZN(g10996), .A(II17901) );
  INV_X1 NOT_3015( .ZN(II17904), .A(g6713) );
  INV_X1 NOT_3016( .ZN(g10999), .A(II17904) );
  INV_X1 NOT_3017( .ZN(II17907), .A(g5824) );
  INV_X1 NOT_3018( .ZN(g11002), .A(II17907) );
  INV_X1 NOT_3019( .ZN(II17910), .A(g7532) );
  INV_X1 NOT_3020( .ZN(g11003), .A(II17910) );
  INV_X1 NOT_3021( .ZN(II17913), .A(g7015) );
  INV_X1 NOT_3022( .ZN(g11004), .A(II17913) );
  INV_X1 NOT_3023( .ZN(II17916), .A(g7560) );
  INV_X1 NOT_3024( .ZN(g11007), .A(II17916) );
  INV_X1 NOT_3025( .ZN(II17919), .A(g7976) );
  INV_X1 NOT_3026( .ZN(g11008), .A(II17919) );
  INV_X1 NOT_3027( .ZN(II17922), .A(g8031) );
  INV_X1 NOT_3028( .ZN(g11011), .A(II17922) );
  INV_X1 NOT_3029( .ZN(II17925), .A(g7976) );
  INV_X1 NOT_3030( .ZN(g11014), .A(II17925) );
  INV_X1 NOT_3031( .ZN(II17928), .A(g8031) );
  INV_X1 NOT_3032( .ZN(g11017), .A(II17928) );
  INV_X1 NOT_3033( .ZN(g11020), .A(g6029) );
  INV_X1 NOT_3034( .ZN(g11021), .A(g6030) );
  INV_X1 NOT_3035( .ZN(II17933), .A(g3254) );
  INV_X1 NOT_3036( .ZN(g11022), .A(II17933) );
  INV_X1 NOT_3037( .ZN(II17936), .A(g6314) );
  INV_X1 NOT_3038( .ZN(g11025), .A(II17936) );
  INV_X1 NOT_3039( .ZN(II17939), .A(g6232) );
  INV_X1 NOT_3040( .ZN(g11028), .A(II17939) );
  INV_X1 NOT_3041( .ZN(II17942), .A(g5548) );
  INV_X1 NOT_3042( .ZN(g11031), .A(II17942) );
  INV_X1 NOT_3043( .ZN(II17945), .A(g5668) );
  INV_X1 NOT_3044( .ZN(g11032), .A(II17945) );
  INV_X1 NOT_3045( .ZN(II17948), .A(g6643) );
  INV_X1 NOT_3046( .ZN(g11035), .A(II17948) );
  INV_X1 NOT_3047( .ZN(II17951), .A(g6519) );
  INV_X1 NOT_3048( .ZN(g11036), .A(II17951) );
  INV_X1 NOT_3049( .ZN(II17954), .A(g6369) );
  INV_X1 NOT_3050( .ZN(g11039), .A(II17954) );
  INV_X1 NOT_3051( .ZN(II17957), .A(g6713) );
  INV_X1 NOT_3052( .ZN(g11042), .A(II17957) );
  INV_X1 NOT_3053( .ZN(II17960), .A(g6945) );
  INV_X1 NOT_3054( .ZN(g11045), .A(II17960) );
  INV_X1 NOT_3055( .ZN(II17963), .A(g6574) );
  INV_X1 NOT_3056( .ZN(g11048), .A(II17963) );
  INV_X1 NOT_3057( .ZN(II17966), .A(g7015) );
  INV_X1 NOT_3058( .ZN(g11051), .A(II17966) );
  INV_X1 NOT_3059( .ZN(II17969), .A(g5880) );
  INV_X1 NOT_3060( .ZN(g11054), .A(II17969) );
  INV_X1 NOT_3061( .ZN(II17972), .A(g7558) );
  INV_X1 NOT_3062( .ZN(g11055), .A(II17972) );
  INV_X1 NOT_3063( .ZN(II17975), .A(g7265) );
  INV_X1 NOT_3064( .ZN(g11056), .A(II17975) );
  INV_X1 NOT_3065( .ZN(II17978), .A(g7795) );
  INV_X1 NOT_3066( .ZN(g11059), .A(II17978) );
  INV_X1 NOT_3067( .ZN(II17981), .A(g7976) );
  INV_X1 NOT_3068( .ZN(g11063), .A(II17981) );
  INV_X1 NOT_3069( .ZN(II17984), .A(g7976) );
  INV_X1 NOT_3070( .ZN(g11066), .A(II17984) );
  INV_X1 NOT_3071( .ZN(g11069), .A(g8257) );
  INV_X1 NOT_3072( .ZN(g11078), .A(g6041) );
  INV_X1 NOT_3073( .ZN(II17989), .A(g3254) );
  INV_X1 NOT_3074( .ZN(g11079), .A(II17989) );
  INV_X1 NOT_3075( .ZN(II17992), .A(g6314) );
  INV_X1 NOT_3076( .ZN(g11082), .A(II17992) );
  INV_X1 NOT_3077( .ZN(II17995), .A(g6232) );
  INV_X1 NOT_3078( .ZN(g11085), .A(II17995) );
  INV_X1 NOT_3079( .ZN(II17998), .A(g5668) );
  INV_X1 NOT_3080( .ZN(g11088), .A(II17998) );
  INV_X1 NOT_3081( .ZN(II18001), .A(g6643) );
  INV_X1 NOT_3082( .ZN(g11091), .A(II18001) );
  INV_X1 NOT_3083( .ZN(II18004), .A(g3410) );
  INV_X1 NOT_3084( .ZN(g11092), .A(II18004) );
  INV_X1 NOT_3085( .ZN(II18007), .A(g6519) );
  INV_X1 NOT_3086( .ZN(g11095), .A(II18007) );
  INV_X1 NOT_3087( .ZN(II18010), .A(g6369) );
  INV_X1 NOT_3088( .ZN(g11098), .A(II18010) );
  INV_X1 NOT_3089( .ZN(II18013), .A(g5594) );
  INV_X1 NOT_3090( .ZN(g11101), .A(II18013) );
  INV_X1 NOT_3091( .ZN(II18016), .A(g5720) );
  INV_X1 NOT_3092( .ZN(g11102), .A(II18016) );
  INV_X1 NOT_3093( .ZN(II18019), .A(g6945) );
  INV_X1 NOT_3094( .ZN(g11105), .A(II18019) );
  INV_X1 NOT_3095( .ZN(II18022), .A(g6783) );
  INV_X1 NOT_3096( .ZN(g11108), .A(II18022) );
  INV_X1 NOT_3097( .ZN(II18025), .A(g6574) );
  INV_X1 NOT_3098( .ZN(g11111), .A(II18025) );
  INV_X1 NOT_3099( .ZN(II18028), .A(g7015) );
  INV_X4 NOT_3100( .ZN(g11114), .A(II18028) );
  INV_X4 NOT_3101( .ZN(II18031), .A(g7195) );
  INV_X4 NOT_3102( .ZN(g11117), .A(II18031) );
  INV_X1 NOT_3103( .ZN(II18034), .A(g6838) );
  INV_X1 NOT_3104( .ZN(g11120), .A(II18034) );
  INV_X1 NOT_3105( .ZN(II18037), .A(g7265) );
  INV_X1 NOT_3106( .ZN(g11123), .A(II18037) );
  INV_X1 NOT_3107( .ZN(II18040), .A(g7976) );
  INV_X1 NOT_3108( .ZN(g11126), .A(II18040) );
  INV_X1 NOT_3109( .ZN(II18043), .A(g7976) );
  INV_X1 NOT_3110( .ZN(g11129), .A(II18043) );
  INV_X1 NOT_3111( .ZN(II18046), .A(g3254) );
  INV_X1 NOT_3112( .ZN(g11132), .A(II18046) );
  INV_X1 NOT_3113( .ZN(II18049), .A(g6314) );
  INV_X1 NOT_3114( .ZN(g11135), .A(II18049) );
  INV_X1 NOT_3115( .ZN(II18052), .A(g6232) );
  INV_X1 NOT_3116( .ZN(g11138), .A(II18052) );
  INV_X1 NOT_3117( .ZN(II18055), .A(g5668) );
  INV_X1 NOT_3118( .ZN(g11141), .A(II18055) );
  INV_X1 NOT_3119( .ZN(II18058), .A(g6643) );
  INV_X1 NOT_3120( .ZN(g11144), .A(II18058) );
  INV_X1 NOT_3121( .ZN(II18061), .A(g3410) );
  INV_X1 NOT_3122( .ZN(g11145), .A(II18061) );
  INV_X1 NOT_3123( .ZN(II18064), .A(g6519) );
  INV_X1 NOT_3124( .ZN(g11148), .A(II18064) );
  INV_X1 NOT_3125( .ZN(II18067), .A(g6369) );
  INV_X1 NOT_3126( .ZN(g11151), .A(II18067) );
  INV_X1 NOT_3127( .ZN(II18070), .A(g5720) );
  INV_X1 NOT_3128( .ZN(g11154), .A(II18070) );
  INV_X1 NOT_3129( .ZN(II18073), .A(g6945) );
  INV_X1 NOT_3130( .ZN(g11157), .A(II18073) );
  INV_X1 NOT_3131( .ZN(II18076), .A(g3566) );
  INV_X1 NOT_3132( .ZN(g11160), .A(II18076) );
  INV_X1 NOT_3133( .ZN(II18079), .A(g6783) );
  INV_X1 NOT_3134( .ZN(g11163), .A(II18079) );
  INV_X1 NOT_3135( .ZN(II18082), .A(g6574) );
  INV_X1 NOT_3136( .ZN(g11166), .A(II18082) );
  INV_X1 NOT_3137( .ZN(II18085), .A(g5611) );
  INV_X1 NOT_3138( .ZN(g11169), .A(II18085) );
  INV_X1 NOT_3139( .ZN(II18088), .A(g5778) );
  INV_X1 NOT_3140( .ZN(g11170), .A(II18088) );
  INV_X1 NOT_3141( .ZN(II18091), .A(g7195) );
  INV_X1 NOT_3142( .ZN(g11173), .A(II18091) );
  INV_X1 NOT_3143( .ZN(II18094), .A(g7085) );
  INV_X1 NOT_3144( .ZN(g11176), .A(II18094) );
  INV_X1 NOT_3145( .ZN(II18097), .A(g6838) );
  INV_X1 NOT_3146( .ZN(g11179), .A(II18097) );
  INV_X1 NOT_3147( .ZN(II18100), .A(g7265) );
  INV_X1 NOT_3148( .ZN(g11182), .A(II18100) );
  INV_X1 NOT_3149( .ZN(II18103), .A(g7391) );
  INV_X1 NOT_3150( .ZN(g11185), .A(II18103) );
  INV_X1 NOT_3151( .ZN(g11190), .A(g3999) );
  INV_X1 NOT_3152( .ZN(II18121), .A(g3254) );
  INV_X1 NOT_3153( .ZN(g11199), .A(II18121) );
  INV_X1 NOT_3154( .ZN(II18124), .A(g6314) );
  INV_X1 NOT_3155( .ZN(g11202), .A(II18124) );
  INV_X1 NOT_3156( .ZN(II18127), .A(g6232) );
  INV_X1 NOT_3157( .ZN(g11205), .A(II18127) );
  INV_X1 NOT_3158( .ZN(II18130), .A(g5547) );
  INV_X1 NOT_3159( .ZN(g11208), .A(II18130) );
  INV_X1 NOT_3160( .ZN(II18133), .A(g6448) );
  INV_X1 NOT_3161( .ZN(g11209), .A(II18133) );
  INV_X1 NOT_3162( .ZN(II18136), .A(g5668) );
  INV_X1 NOT_3163( .ZN(g11210), .A(II18136) );
  INV_X1 NOT_3164( .ZN(II18139), .A(g6643) );
  INV_X1 NOT_3165( .ZN(g11213), .A(II18139) );
  INV_X1 NOT_3166( .ZN(II18142), .A(g3410) );
  INV_X1 NOT_3167( .ZN(g11216), .A(II18142) );
  INV_X1 NOT_3168( .ZN(II18145), .A(g6519) );
  INV_X1 NOT_3169( .ZN(g11219), .A(II18145) );
  INV_X1 NOT_3170( .ZN(II18148), .A(g6369) );
  INV_X1 NOT_3171( .ZN(g11222), .A(II18148) );
  INV_X1 NOT_3172( .ZN(II18151), .A(g5720) );
  INV_X1 NOT_3173( .ZN(g11225), .A(II18151) );
  INV_X1 NOT_3174( .ZN(II18154), .A(g6945) );
  INV_X1 NOT_3175( .ZN(g11228), .A(II18154) );
  INV_X1 NOT_3176( .ZN(II18157), .A(g3566) );
  INV_X1 NOT_3177( .ZN(g11231), .A(II18157) );
  INV_X1 NOT_3178( .ZN(II18160), .A(g6783) );
  INV_X1 NOT_3179( .ZN(g11234), .A(II18160) );
  INV_X1 NOT_3180( .ZN(II18163), .A(g6574) );
  INV_X1 NOT_3181( .ZN(g11237), .A(II18163) );
  INV_X1 NOT_3182( .ZN(II18166), .A(g5778) );
  INV_X1 NOT_3183( .ZN(g11240), .A(II18166) );
  INV_X1 NOT_3184( .ZN(II18169), .A(g7195) );
  INV_X1 NOT_3185( .ZN(g11243), .A(II18169) );
  INV_X1 NOT_3186( .ZN(II18172), .A(g3722) );
  INV_X1 NOT_3187( .ZN(g11246), .A(II18172) );
  INV_X1 NOT_3188( .ZN(II18175), .A(g7085) );
  INV_X1 NOT_3189( .ZN(g11249), .A(II18175) );
  INV_X1 NOT_3190( .ZN(II18178), .A(g6838) );
  INV_X1 NOT_3191( .ZN(g11252), .A(II18178) );
  INV_X1 NOT_3192( .ZN(II18181), .A(g5636) );
  INV_X1 NOT_3193( .ZN(g11255), .A(II18181) );
  INV_X1 NOT_3194( .ZN(II18184), .A(g5837) );
  INV_X1 NOT_3195( .ZN(g11256), .A(II18184) );
  INV_X1 NOT_3196( .ZN(II18187), .A(g7391) );
  INV_X1 NOT_3197( .ZN(g11259), .A(II18187) );
  INV_X1 NOT_3198( .ZN(II18211), .A(g6232) );
  INV_X1 NOT_3199( .ZN(g11265), .A(II18211) );
  INV_X1 NOT_3200( .ZN(II18214), .A(g3254) );
  INV_X1 NOT_3201( .ZN(g11268), .A(II18214) );
  INV_X1 NOT_3202( .ZN(II18217), .A(g6314) );
  INV_X1 NOT_3203( .ZN(g11271), .A(II18217) );
  INV_X1 NOT_3204( .ZN(II18220), .A(g6232) );
  INV_X1 NOT_3205( .ZN(g11274), .A(II18220) );
  INV_X1 NOT_3206( .ZN(II18223), .A(g6448) );
  INV_X1 NOT_3207( .ZN(g11277), .A(II18223) );
  INV_X1 NOT_3208( .ZN(II18226), .A(g5668) );
  INV_X1 NOT_3209( .ZN(g11278), .A(II18226) );
  INV_X1 NOT_3210( .ZN(II18229), .A(g3410) );
  INV_X1 NOT_3211( .ZN(g11281), .A(II18229) );
  INV_X1 NOT_3212( .ZN(II18232), .A(g6519) );
  INV_X1 NOT_3213( .ZN(g11284), .A(II18232) );
  INV_X1 NOT_3214( .ZN(II18235), .A(g6369) );
  INV_X1 NOT_3215( .ZN(g11287), .A(II18235) );
  INV_X1 NOT_3216( .ZN(II18238), .A(g5593) );
  INV_X1 NOT_3217( .ZN(g11290), .A(II18238) );
  INV_X1 NOT_3218( .ZN(II18241), .A(g6713) );
  INV_X1 NOT_3219( .ZN(g11291), .A(II18241) );
  INV_X1 NOT_3220( .ZN(II18244), .A(g5720) );
  INV_X1 NOT_3221( .ZN(g11294), .A(II18244) );
  INV_X1 NOT_3222( .ZN(II18247), .A(g6945) );
  INV_X1 NOT_3223( .ZN(g11297), .A(II18247) );
  INV_X1 NOT_3224( .ZN(II18250), .A(g3566) );
  INV_X1 NOT_3225( .ZN(g11300), .A(II18250) );
  INV_X1 NOT_3226( .ZN(II18253), .A(g6783) );
  INV_X1 NOT_3227( .ZN(g11303), .A(II18253) );
  INV_X1 NOT_3228( .ZN(II18256), .A(g6574) );
  INV_X1 NOT_3229( .ZN(g11306), .A(II18256) );
  INV_X1 NOT_3230( .ZN(II18259), .A(g5778) );
  INV_X1 NOT_3231( .ZN(g11309), .A(II18259) );
  INV_X1 NOT_3232( .ZN(II18262), .A(g7195) );
  INV_X1 NOT_3233( .ZN(g11312), .A(II18262) );
  INV_X1 NOT_3234( .ZN(II18265), .A(g3722) );
  INV_X1 NOT_3235( .ZN(g11315), .A(II18265) );
  INV_X1 NOT_3236( .ZN(II18268), .A(g7085) );
  INV_X1 NOT_3237( .ZN(g11318), .A(II18268) );
  INV_X1 NOT_3238( .ZN(II18271), .A(g6838) );
  INV_X1 NOT_3239( .ZN(g11321), .A(II18271) );
  INV_X1 NOT_3240( .ZN(II18274), .A(g5837) );
  INV_X1 NOT_3241( .ZN(g11324), .A(II18274) );
  INV_X1 NOT_3242( .ZN(II18277), .A(g7391) );
  INV_X1 NOT_3243( .ZN(g11327), .A(II18277) );
  INV_X1 NOT_3244( .ZN(g11332), .A(g4094) );
  INV_X1 NOT_3245( .ZN(II18295), .A(g6314) );
  INV_X1 NOT_3246( .ZN(g11341), .A(II18295) );
  INV_X1 NOT_3247( .ZN(II18298), .A(g6232) );
  INV_X1 NOT_3248( .ZN(g11344), .A(II18298) );
  INV_X1 NOT_3249( .ZN(II18302), .A(g3254) );
  INV_X1 NOT_3250( .ZN(g11348), .A(II18302) );
  INV_X1 NOT_3251( .ZN(II18305), .A(g6314) );
  INV_X1 NOT_3252( .ZN(g11351), .A(II18305) );
  INV_X1 NOT_3253( .ZN(II18308), .A(g6448) );
  INV_X1 NOT_3254( .ZN(g11354), .A(II18308) );
  INV_X1 NOT_3255( .ZN(II18311), .A(g5668) );
  INV_X1 NOT_3256( .ZN(g11355), .A(II18311) );
  INV_X1 NOT_3257( .ZN(II18314), .A(g6369) );
  INV_X1 NOT_3258( .ZN(g11358), .A(II18314) );
  INV_X1 NOT_3259( .ZN(II18317), .A(g3410) );
  INV_X1 NOT_3260( .ZN(g11361), .A(II18317) );
  INV_X1 NOT_3261( .ZN(II18320), .A(g6519) );
  INV_X1 NOT_3262( .ZN(g11364), .A(II18320) );
  INV_X1 NOT_3263( .ZN(II18323), .A(g6369) );
  INV_X1 NOT_3264( .ZN(g11367), .A(II18323) );
  INV_X1 NOT_3265( .ZN(II18326), .A(g6713) );
  INV_X1 NOT_3266( .ZN(g11370), .A(II18326) );
  INV_X1 NOT_3267( .ZN(II18329), .A(g5720) );
  INV_X1 NOT_3268( .ZN(g11373), .A(II18329) );
  INV_X1 NOT_3269( .ZN(II18332), .A(g3566) );
  INV_X1 NOT_3270( .ZN(g11376), .A(II18332) );
  INV_X1 NOT_3271( .ZN(II18335), .A(g6783) );
  INV_X1 NOT_3272( .ZN(g11379), .A(II18335) );
  INV_X1 NOT_3273( .ZN(II18338), .A(g6574) );
  INV_X1 NOT_3274( .ZN(g11382), .A(II18338) );
  INV_X1 NOT_3275( .ZN(II18341), .A(g5610) );
  INV_X2 NOT_3276( .ZN(g11385), .A(II18341) );
  INV_X2 NOT_3277( .ZN(II18344), .A(g7015) );
  INV_X2 NOT_3278( .ZN(g11386), .A(II18344) );
  INV_X2 NOT_3279( .ZN(II18347), .A(g5778) );
  INV_X2 NOT_3280( .ZN(g11389), .A(II18347) );
  INV_X1 NOT_3281( .ZN(II18350), .A(g7195) );
  INV_X1 NOT_3282( .ZN(g11392), .A(II18350) );
  INV_X1 NOT_3283( .ZN(II18353), .A(g3722) );
  INV_X1 NOT_3284( .ZN(g11395), .A(II18353) );
  INV_X1 NOT_3285( .ZN(II18356), .A(g7085) );
  INV_X1 NOT_3286( .ZN(g11398), .A(II18356) );
  INV_X1 NOT_3287( .ZN(II18359), .A(g6838) );
  INV_X1 NOT_3288( .ZN(g11401), .A(II18359) );
  INV_X1 NOT_3289( .ZN(II18362), .A(g5837) );
  INV_X1 NOT_3290( .ZN(g11404), .A(II18362) );
  INV_X1 NOT_3291( .ZN(II18365), .A(g7391) );
  INV_X1 NOT_3292( .ZN(g11407), .A(II18365) );
  INV_X1 NOT_3293( .ZN(II18375), .A(g3254) );
  INV_X1 NOT_3294( .ZN(g11411), .A(II18375) );
  INV_X1 NOT_3295( .ZN(II18378), .A(g6314) );
  INV_X1 NOT_3296( .ZN(g11414), .A(II18378) );
  INV_X1 NOT_3297( .ZN(II18381), .A(g6232) );
  INV_X1 NOT_3298( .ZN(g11417), .A(II18381) );
  INV_X1 NOT_3299( .ZN(II18386), .A(g3254) );
  INV_X1 NOT_3300( .ZN(g11422), .A(II18386) );
  INV_X1 NOT_3301( .ZN(II18389), .A(g6519) );
  INV_X1 NOT_3302( .ZN(g11425), .A(II18389) );
  INV_X1 NOT_3303( .ZN(II18392), .A(g6369) );
  INV_X1 NOT_3304( .ZN(g11428), .A(II18392) );
  INV_X1 NOT_3305( .ZN(II18396), .A(g3410) );
  INV_X1 NOT_3306( .ZN(g11432), .A(II18396) );
  INV_X1 NOT_3307( .ZN(II18399), .A(g6519) );
  INV_X1 NOT_3308( .ZN(g11435), .A(II18399) );
  INV_X1 NOT_3309( .ZN(II18402), .A(g6713) );
  INV_X1 NOT_3310( .ZN(g11438), .A(II18402) );
  INV_X1 NOT_3311( .ZN(II18405), .A(g5720) );
  INV_X1 NOT_3312( .ZN(g11441), .A(II18405) );
  INV_X1 NOT_3313( .ZN(II18408), .A(g6574) );
  INV_X1 NOT_3314( .ZN(g11444), .A(II18408) );
  INV_X1 NOT_3315( .ZN(II18411), .A(g3566) );
  INV_X1 NOT_3316( .ZN(g11447), .A(II18411) );
  INV_X1 NOT_3317( .ZN(II18414), .A(g6783) );
  INV_X1 NOT_3318( .ZN(g11450), .A(II18414) );
  INV_X1 NOT_3319( .ZN(II18417), .A(g6574) );
  INV_X1 NOT_3320( .ZN(g11453), .A(II18417) );
  INV_X1 NOT_3321( .ZN(II18420), .A(g7015) );
  INV_X1 NOT_3322( .ZN(g11456), .A(II18420) );
  INV_X1 NOT_3323( .ZN(II18423), .A(g5778) );
  INV_X1 NOT_3324( .ZN(g11459), .A(II18423) );
  INV_X1 NOT_3325( .ZN(II18426), .A(g3722) );
  INV_X1 NOT_3326( .ZN(g11462), .A(II18426) );
  INV_X1 NOT_3327( .ZN(II18429), .A(g7085) );
  INV_X1 NOT_3328( .ZN(g11465), .A(II18429) );
  INV_X1 NOT_3329( .ZN(II18432), .A(g6838) );
  INV_X1 NOT_3330( .ZN(g11468), .A(II18432) );
  INV_X1 NOT_3331( .ZN(II18435), .A(g5635) );
  INV_X1 NOT_3332( .ZN(g11471), .A(II18435) );
  INV_X1 NOT_3333( .ZN(II18438), .A(g7265) );
  INV_X1 NOT_3334( .ZN(g11472), .A(II18438) );
  INV_X1 NOT_3335( .ZN(II18441), .A(g5837) );
  INV_X1 NOT_3336( .ZN(g11475), .A(II18441) );
  INV_X1 NOT_3337( .ZN(II18444), .A(g7391) );
  INV_X1 NOT_3338( .ZN(g11478), .A(II18444) );
  INV_X1 NOT_3339( .ZN(g11481), .A(g4204) );
  INV_X1 NOT_3340( .ZN(g11490), .A(g8276) );
  INV_X1 NOT_3341( .ZN(II18449), .A(g10868) );
  INV_X1 NOT_3342( .ZN(g11491), .A(II18449) );
  INV_X1 NOT_3343( .ZN(II18452), .A(g10930) );
  INV_X1 NOT_3344( .ZN(g11492), .A(II18452) );
  INV_X1 NOT_3345( .ZN(II18455), .A(g11031) );
  INV_X1 NOT_3346( .ZN(g11493), .A(II18455) );
  INV_X1 NOT_3347( .ZN(II18458), .A(g11208) );
  INV_X1 NOT_3348( .ZN(g11494), .A(II18458) );
  INV_X1 NOT_3349( .ZN(II18461), .A(g10931) );
  INV_X1 NOT_3350( .ZN(g11495), .A(II18461) );
  INV_X1 NOT_3351( .ZN(II18464), .A(g8620) );
  INV_X1 NOT_3352( .ZN(g11496), .A(II18464) );
  INV_X1 NOT_3353( .ZN(II18467), .A(g8769) );
  INV_X1 NOT_3354( .ZN(g11497), .A(II18467) );
  INV_X1 NOT_3355( .ZN(II18470), .A(g8808) );
  INV_X1 NOT_3356( .ZN(g11498), .A(II18470) );
  INV_X1 NOT_3357( .ZN(II18473), .A(g8839) );
  INV_X1 NOT_3358( .ZN(g11499), .A(II18473) );
  INV_X1 NOT_3359( .ZN(II18476), .A(g8791) );
  INV_X1 NOT_3360( .ZN(g11500), .A(II18476) );
  INV_X1 NOT_3361( .ZN(II18479), .A(g8820) );
  INV_X1 NOT_3362( .ZN(g11501), .A(II18479) );
  INV_X1 NOT_3363( .ZN(II18482), .A(g8859) );
  INV_X1 NOT_3364( .ZN(g11502), .A(II18482) );
  INV_X1 NOT_3365( .ZN(II18485), .A(g8809) );
  INV_X1 NOT_3366( .ZN(g11503), .A(II18485) );
  INV_X1 NOT_3367( .ZN(II18488), .A(g8840) );
  INV_X1 NOT_3368( .ZN(g11504), .A(II18488) );
  INV_X1 NOT_3369( .ZN(II18491), .A(g8891) );
  INV_X1 NOT_3370( .ZN(g11505), .A(II18491) );
  INV_X1 NOT_3371( .ZN(II18494), .A(g8821) );
  INV_X1 NOT_3372( .ZN(g11506), .A(II18494) );
  INV_X1 NOT_3373( .ZN(II18497), .A(g8860) );
  INV_X1 NOT_3374( .ZN(g11507), .A(II18497) );
  INV_X1 NOT_3375( .ZN(II18500), .A(g8924) );
  INV_X1 NOT_3376( .ZN(g11508), .A(II18500) );
  INV_X1 NOT_3377( .ZN(II18503), .A(g8658) );
  INV_X1 NOT_3378( .ZN(g11509), .A(II18503) );
  INV_X1 NOT_3379( .ZN(II18506), .A(g8699) );
  INV_X1 NOT_3380( .ZN(g11510), .A(II18506) );
  INV_X1 NOT_3381( .ZN(II18509), .A(g8770) );
  INV_X1 NOT_3382( .ZN(g11511), .A(II18509) );
  INV_X1 NOT_3383( .ZN(II18512), .A(g9309) );
  INV_X1 NOT_3384( .ZN(g11512), .A(II18512) );
  INV_X1 NOT_3385( .ZN(II18515), .A(g8843) );
  INV_X1 NOT_3386( .ZN(g11513), .A(II18515) );
  INV_X2 NOT_3387( .ZN(II18518), .A(g8893) );
  INV_X2 NOT_3388( .ZN(g11514), .A(II18518) );
  INV_X2 NOT_3389( .ZN(II18521), .A(g9449) );
  INV_X2 NOT_3390( .ZN(g11515), .A(II18521) );
  INV_X2 NOT_3391( .ZN(II18524), .A(g9640) );
  INV_X1 NOT_3392( .ZN(g11516), .A(II18524) );
  INV_X1 NOT_3393( .ZN(II18527), .A(g10017) );
  INV_X1 NOT_3394( .ZN(g11517), .A(II18527) );
  INV_X1 NOT_3395( .ZN(II18530), .A(g10888) );
  INV_X1 NOT_3396( .ZN(g11518), .A(II18530) );
  INV_X1 NOT_3397( .ZN(II18533), .A(g10967) );
  INV_X1 NOT_3398( .ZN(g11519), .A(II18533) );
  INV_X1 NOT_3399( .ZN(II18536), .A(g11101) );
  INV_X1 NOT_3400( .ZN(g11520), .A(II18536) );
  INV_X1 NOT_3401( .ZN(II18539), .A(g11290) );
  INV_X1 NOT_3402( .ZN(g11521), .A(II18539) );
  INV_X1 NOT_3403( .ZN(II18542), .A(g10968) );
  INV_X1 NOT_3404( .ZN(g11522), .A(II18542) );
  INV_X1 NOT_3405( .ZN(II18545), .A(g8630) );
  INV_X1 NOT_3406( .ZN(g11523), .A(II18545) );
  INV_X1 NOT_3407( .ZN(II18548), .A(g8792) );
  INV_X1 NOT_3408( .ZN(g11524), .A(II18548) );
  INV_X1 NOT_3409( .ZN(II18551), .A(g8824) );
  INV_X1 NOT_3410( .ZN(g11525), .A(II18551) );
  INV_X1 NOT_3411( .ZN(II18554), .A(g8866) );
  INV_X1 NOT_3412( .ZN(g11526), .A(II18554) );
  INV_X1 NOT_3413( .ZN(II18557), .A(g8810) );
  INV_X1 NOT_3414( .ZN(g11527), .A(II18557) );
  INV_X1 NOT_3415( .ZN(II18560), .A(g8844) );
  INV_X1 NOT_3416( .ZN(g11528), .A(II18560) );
  INV_X1 NOT_3417( .ZN(II18563), .A(g8897) );
  INV_X1 NOT_3418( .ZN(g11529), .A(II18563) );
  INV_X1 NOT_3419( .ZN(II18566), .A(g8825) );
  INV_X1 NOT_3420( .ZN(g11530), .A(II18566) );
  INV_X1 NOT_3421( .ZN(II18569), .A(g8867) );
  INV_X1 NOT_3422( .ZN(g11531), .A(II18569) );
  INV_X1 NOT_3423( .ZN(II18572), .A(g8931) );
  INV_X1 NOT_3424( .ZN(g11532), .A(II18572) );
  INV_X1 NOT_3425( .ZN(II18575), .A(g8845) );
  INV_X1 NOT_3426( .ZN(g11533), .A(II18575) );
  INV_X1 NOT_3427( .ZN(II18578), .A(g8898) );
  INV_X1 NOT_3428( .ZN(g11534), .A(II18578) );
  INV_X1 NOT_3429( .ZN(II18581), .A(g8964) );
  INV_X1 NOT_3430( .ZN(g11535), .A(II18581) );
  INV_X1 NOT_3431( .ZN(II18584), .A(g8677) );
  INV_X1 NOT_3432( .ZN(g11536), .A(II18584) );
  INV_X1 NOT_3433( .ZN(II18587), .A(g8718) );
  INV_X1 NOT_3434( .ZN(g11537), .A(II18587) );
  INV_X1 NOT_3435( .ZN(II18590), .A(g8793) );
  INV_X1 NOT_3436( .ZN(g11538), .A(II18590) );
  INV_X1 NOT_3437( .ZN(II18593), .A(g9390) );
  INV_X1 NOT_3438( .ZN(g11539), .A(II18593) );
  INV_X1 NOT_3439( .ZN(II18596), .A(g8870) );
  INV_X1 NOT_3440( .ZN(g11540), .A(II18596) );
  INV_X1 NOT_3441( .ZN(II18599), .A(g8933) );
  INV_X1 NOT_3442( .ZN(g11541), .A(II18599) );
  INV_X1 NOT_3443( .ZN(II18602), .A(g9591) );
  INV_X1 NOT_3444( .ZN(g11542), .A(II18602) );
  INV_X1 NOT_3445( .ZN(II18605), .A(g9786) );
  INV_X1 NOT_3446( .ZN(g11543), .A(II18605) );
  INV_X1 NOT_3447( .ZN(II18608), .A(g10126) );
  INV_X1 NOT_3448( .ZN(g11544), .A(II18608) );
  INV_X1 NOT_3449( .ZN(II18611), .A(g10909) );
  INV_X1 NOT_3450( .ZN(g11545), .A(II18611) );
  INV_X1 NOT_3451( .ZN(II18614), .A(g11002) );
  INV_X1 NOT_3452( .ZN(g11546), .A(II18614) );
  INV_X1 NOT_3453( .ZN(II18617), .A(g11169) );
  INV_X1 NOT_3454( .ZN(g11547), .A(II18617) );
  INV_X1 NOT_3455( .ZN(II18620), .A(g11385) );
  INV_X1 NOT_3456( .ZN(g11548), .A(II18620) );
  INV_X1 NOT_3457( .ZN(II18623), .A(g11003) );
  INV_X1 NOT_3458( .ZN(g11549), .A(II18623) );
  INV_X1 NOT_3459( .ZN(II18626), .A(g8649) );
  INV_X1 NOT_3460( .ZN(g11550), .A(II18626) );
  INV_X1 NOT_3461( .ZN(II18629), .A(g8811) );
  INV_X1 NOT_3462( .ZN(g11551), .A(II18629) );
  INV_X1 NOT_3463( .ZN(II18632), .A(g8850) );
  INV_X1 NOT_3464( .ZN(g11552), .A(II18632) );
  INV_X1 NOT_3465( .ZN(II18635), .A(g8904) );
  INV_X1 NOT_3466( .ZN(g11553), .A(II18635) );
  INV_X1 NOT_3467( .ZN(II18638), .A(g8826) );
  INV_X1 NOT_3468( .ZN(g11554), .A(II18638) );
  INV_X1 NOT_3469( .ZN(II18641), .A(g8871) );
  INV_X1 NOT_3470( .ZN(g11555), .A(II18641) );
  INV_X1 NOT_3471( .ZN(II18644), .A(g8937) );
  INV_X1 NOT_3472( .ZN(g11556), .A(II18644) );
  INV_X1 NOT_3473( .ZN(II18647), .A(g8851) );
  INV_X1 NOT_3474( .ZN(g11557), .A(II18647) );
  INV_X1 NOT_3475( .ZN(II18650), .A(g8905) );
  INV_X1 NOT_3476( .ZN(g11558), .A(II18650) );
  INV_X1 NOT_3477( .ZN(II18653), .A(g8971) );
  INV_X1 NOT_3478( .ZN(g11559), .A(II18653) );
  INV_X1 NOT_3479( .ZN(II18656), .A(g8872) );
  INV_X1 NOT_3480( .ZN(g11560), .A(II18656) );
  INV_X1 NOT_3481( .ZN(II18659), .A(g8938) );
  INV_X1 NOT_3482( .ZN(g11561), .A(II18659) );
  INV_X1 NOT_3483( .ZN(II18662), .A(g8996) );
  INV_X1 NOT_3484( .ZN(g11562), .A(II18662) );
  INV_X1 NOT_3485( .ZN(II18665), .A(g8689) );
  INV_X1 NOT_3486( .ZN(g11563), .A(II18665) );
  INV_X1 NOT_3487( .ZN(II18668), .A(g8756) );
  INV_X1 NOT_3488( .ZN(g11564), .A(II18668) );
  INV_X1 NOT_3489( .ZN(II18671), .A(g8812) );
  INV_X1 NOT_3490( .ZN(g11565), .A(II18671) );
  INV_X1 NOT_3491( .ZN(II18674), .A(g9487) );
  INV_X1 NOT_3492( .ZN(g11566), .A(II18674) );
  INV_X1 NOT_3493( .ZN(II18677), .A(g8908) );
  INV_X1 NOT_3494( .ZN(g11567), .A(II18677) );
  INV_X1 NOT_3495( .ZN(II18680), .A(g8973) );
  INV_X1 NOT_3496( .ZN(g11568), .A(II18680) );
  INV_X1 NOT_3497( .ZN(II18683), .A(g9733) );
  INV_X1 NOT_3498( .ZN(g11569), .A(II18683) );
  INV_X1 NOT_3499( .ZN(II18686), .A(g9932) );
  INV_X1 NOT_3500( .ZN(g11570), .A(II18686) );
  INV_X1 NOT_3501( .ZN(II18689), .A(g10231) );
  INV_X1 NOT_3502( .ZN(g11571), .A(II18689) );
  INV_X1 NOT_3503( .ZN(II18692), .A(g10935) );
  INV_X1 NOT_3504( .ZN(g11572), .A(II18692) );
  INV_X1 NOT_3505( .ZN(II18695), .A(g11054) );
  INV_X1 NOT_3506( .ZN(g11573), .A(II18695) );
  INV_X1 NOT_3507( .ZN(II18698), .A(g11255) );
  INV_X1 NOT_3508( .ZN(g11574), .A(II18698) );
  INV_X1 NOT_3509( .ZN(II18701), .A(g11471) );
  INV_X1 NOT_3510( .ZN(g11575), .A(II18701) );
  INV_X1 NOT_3511( .ZN(II18704), .A(g11055) );
  INV_X2 NOT_3512( .ZN(g11576), .A(II18704) );
  INV_X2 NOT_3513( .ZN(II18707), .A(g8665) );
  INV_X1 NOT_3514( .ZN(g11577), .A(II18707) );
  INV_X1 NOT_3515( .ZN(II18710), .A(g8827) );
  INV_X1 NOT_3516( .ZN(g11578), .A(II18710) );
  INV_X1 NOT_3517( .ZN(II18713), .A(g8877) );
  INV_X1 NOT_3518( .ZN(g11579), .A(II18713) );
  INV_X1 NOT_3519( .ZN(II18716), .A(g8944) );
  INV_X1 NOT_3520( .ZN(g11580), .A(II18716) );
  INV_X1 NOT_3521( .ZN(II18719), .A(g8852) );
  INV_X1 NOT_3522( .ZN(g11581), .A(II18719) );
  INV_X1 NOT_3523( .ZN(II18722), .A(g8909) );
  INV_X1 NOT_3524( .ZN(g11582), .A(II18722) );
  INV_X1 NOT_3525( .ZN(II18725), .A(g8977) );
  INV_X1 NOT_3526( .ZN(g11583), .A(II18725) );
  INV_X1 NOT_3527( .ZN(II18728), .A(g8878) );
  INV_X1 NOT_3528( .ZN(g11584), .A(II18728) );
  INV_X1 NOT_3529( .ZN(II18731), .A(g8945) );
  INV_X1 NOT_3530( .ZN(g11585), .A(II18731) );
  INV_X1 NOT_3531( .ZN(II18734), .A(g9003) );
  INV_X1 NOT_3532( .ZN(g11586), .A(II18734) );
  INV_X1 NOT_3533( .ZN(II18737), .A(g8910) );
  INV_X1 NOT_3534( .ZN(g11587), .A(II18737) );
  INV_X1 NOT_3535( .ZN(II18740), .A(g8978) );
  INV_X1 NOT_3536( .ZN(g11588), .A(II18740) );
  INV_X1 NOT_3537( .ZN(II18743), .A(g9025) );
  INV_X1 NOT_3538( .ZN(g11589), .A(II18743) );
  INV_X1 NOT_3539( .ZN(II18746), .A(g8707) );
  INV_X1 NOT_3540( .ZN(g11590), .A(II18746) );
  INV_X1 NOT_3541( .ZN(II18749), .A(g8779) );
  INV_X1 NOT_3542( .ZN(g11591), .A(II18749) );
  INV_X1 NOT_3543( .ZN(II18752), .A(g8828) );
  INV_X1 NOT_3544( .ZN(g11592), .A(II18752) );
  INV_X1 NOT_3545( .ZN(II18755), .A(g9629) );
  INV_X1 NOT_3546( .ZN(g11593), .A(II18755) );
  INV_X1 NOT_3547( .ZN(II18758), .A(g8948) );
  INV_X1 NOT_3548( .ZN(g11594), .A(II18758) );
  INV_X1 NOT_3549( .ZN(II18761), .A(g9005) );
  INV_X1 NOT_3550( .ZN(g11595), .A(II18761) );
  INV_X1 NOT_3551( .ZN(II18764), .A(g9879) );
  INV_X1 NOT_3552( .ZN(g11596), .A(II18764) );
  INV_X1 NOT_3553( .ZN(II18767), .A(g10086) );
  INV_X1 NOT_3554( .ZN(g11597), .A(II18767) );
  INV_X1 NOT_3555( .ZN(II18770), .A(g10333) );
  INV_X1 NOT_3556( .ZN(g11598), .A(II18770) );
  INV_X1 NOT_3557( .ZN(II18773), .A(g10830) );
  INV_X1 NOT_3558( .ZN(g11599), .A(II18773) );
  INV_X1 NOT_3559( .ZN(II18777), .A(g9050) );
  INV_X1 NOT_3560( .ZN(g11603), .A(II18777) );
  INV_X1 NOT_3561( .ZN(II18780), .A(g10870) );
  INV_X1 NOT_3562( .ZN(g11606), .A(II18780) );
  INV_X1 NOT_3563( .ZN(II18784), .A(g9067) );
  INV_X1 NOT_3564( .ZN(g11608), .A(II18784) );
  INV_X1 NOT_3565( .ZN(II18787), .A(g10910) );
  INV_X1 NOT_3566( .ZN(g11611), .A(II18787) );
  INV_X1 NOT_3567( .ZN(II18791), .A(g9084) );
  INV_X1 NOT_3568( .ZN(g11613), .A(II18791) );
  INV_X1 NOT_3569( .ZN(II18794), .A(g10973) );
  INV_X1 NOT_3570( .ZN(g11616), .A(II18794) );
  INV_X1 NOT_3571( .ZN(g11620), .A(g10601) );
  INV_X1 NOT_3572( .ZN(g11623), .A(g10961) );
  INV_X1 NOT_3573( .ZN(II18810), .A(g10813) );
  INV_X1 NOT_3574( .ZN(g11628), .A(II18810) );
  INV_X1 NOT_3575( .ZN(II18813), .A(g10850) );
  INV_X1 NOT_3576( .ZN(g11629), .A(II18813) );
  INV_X1 NOT_3577( .ZN(II18817), .A(g9067) );
  INV_X1 NOT_3578( .ZN(g11633), .A(II18817) );
  INV_X1 NOT_3579( .ZN(II18820), .A(g10890) );
  INV_X1 NOT_3580( .ZN(g11636), .A(II18820) );
  INV_X1 NOT_3581( .ZN(II18824), .A(g9084) );
  INV_X1 NOT_3582( .ZN(g11638), .A(II18824) );
  INV_X1 NOT_3583( .ZN(II18827), .A(g10936) );
  INV_X1 NOT_3584( .ZN(g11641), .A(II18827) );
  INV_X1 NOT_3585( .ZN(g11642), .A(g10646) );
  INV_X1 NOT_3586( .ZN(II18835), .A(g10834) );
  INV_X1 NOT_3587( .ZN(g11651), .A(II18835) );
  INV_X1 NOT_3588( .ZN(II18838), .A(g10871) );
  INV_X1 NOT_3589( .ZN(g11652), .A(II18838) );
  INV_X1 NOT_3590( .ZN(II18842), .A(g9084) );
  INV_X1 NOT_3591( .ZN(g11656), .A(II18842) );
  INV_X1 NOT_3592( .ZN(II18845), .A(g10911) );
  INV_X1 NOT_3593( .ZN(g11659), .A(II18845) );
  INV_X1 NOT_3594( .ZN(II18854), .A(g10854) );
  INV_X1 NOT_3595( .ZN(g11670), .A(II18854) );
  INV_X1 NOT_3596( .ZN(II18857), .A(g10891) );
  INV_X1 NOT_3597( .ZN(g11671), .A(II18857) );
  INV_X1 NOT_3598( .ZN(II18866), .A(g10875) );
  INV_X1 NOT_3599( .ZN(g11682), .A(II18866) );
  INV_X1 NOT_3600( .ZN(g11706), .A(g10928) );
  INV_X1 NOT_3601( .ZN(g11732), .A(g10826) );
  INV_X1 NOT_3602( .ZN(g11734), .A(g10843) );
  INV_X1 NOT_3603( .ZN(g11735), .A(g10859) );
  INV_X1 NOT_3604( .ZN(g11736), .A(g10862) );
  INV_X1 NOT_3605( .ZN(g11737), .A(g10809) );
  INV_X1 NOT_3606( .ZN(g11740), .A(g10877) );
  INV_X1 NOT_3607( .ZN(g11741), .A(g10880) );
  INV_X1 NOT_3608( .ZN(g11742), .A(g10883) );
  INV_X1 NOT_3609( .ZN(g11743), .A(g8530) );
  INV_X1 NOT_3610( .ZN(g11745), .A(g10892) );
  INV_X1 NOT_3611( .ZN(g11746), .A(g10895) );
  INV_X1 NOT_3612( .ZN(g11747), .A(g10898) );
  INV_X1 NOT_3613( .ZN(g11748), .A(g10901) );
  INV_X1 NOT_3614( .ZN(II18929), .A(g10711) );
  INV_X1 NOT_3615( .ZN(g11749), .A(II18929) );
  INV_X1 NOT_3616( .ZN(g11758), .A(g8514) );
  INV_X1 NOT_3617( .ZN(g11761), .A(g10912) );
  INV_X1 NOT_3618( .ZN(g11762), .A(g10915) );
  INV_X1 NOT_3619( .ZN(g11763), .A(g10918) );
  INV_X1 NOT_3620( .ZN(g11764), .A(g10921) );
  INV_X1 NOT_3621( .ZN(g11765), .A(g10924) );
  INV_X1 NOT_3622( .ZN(g11766), .A(g10886) );
  INV_X1 NOT_3623( .ZN(II18943), .A(g9149) );
  INV_X1 NOT_3624( .ZN(g11769), .A(II18943) );
  INV_X1 NOT_3625( .ZN(g11770), .A(g10932) );
  INV_X1 NOT_3626( .ZN(g11774), .A(g10937) );
  INV_X1 NOT_3627( .ZN(g11775), .A(g10940) );
  INV_X1 NOT_3628( .ZN(g11776), .A(g10943) );
  INV_X1 NOT_3629( .ZN(g11777), .A(g10946) );
  INV_X1 NOT_3630( .ZN(g11778), .A(g10949) );
  INV_X1 NOT_3631( .ZN(g11779), .A(g10906) );
  INV_X1 NOT_3632( .ZN(g11782), .A(g10963) );
  INV_X1 NOT_3633( .ZN(g11783), .A(g10966) );
  INV_X1 NOT_3634( .ZN(II18962), .A(g9159) );
  INV_X1 NOT_3635( .ZN(g11786), .A(II18962) );
  INV_X1 NOT_3636( .ZN(g11787), .A(g10969) );
  INV_X1 NOT_3637( .ZN(II18969), .A(g8726) );
  INV_X1 NOT_3638( .ZN(g11791), .A(II18969) );
  INV_X1 NOT_3639( .ZN(g11794), .A(g10974) );
  INV_X1 NOT_3640( .ZN(g11795), .A(g10977) );
  INV_X1 NOT_3641( .ZN(g11796), .A(g10980) );
  INV_X1 NOT_3642( .ZN(g11797), .A(g10983) );
  INV_X1 NOT_3643( .ZN(g11798), .A(g10867) );
  INV_X1 NOT_3644( .ZN(g11801), .A(g10988) );
  INV_X1 NOT_3645( .ZN(g11802), .A(g10991) );
  INV_X1 NOT_3646( .ZN(g11803), .A(g10994) );
  INV_X1 NOT_3647( .ZN(g11804), .A(g10995) );
  INV_X1 NOT_3648( .ZN(g11808), .A(g10996) );
  INV_X1 NOT_3649( .ZN(g11809), .A(g10999) );
  INV_X1 NOT_3650( .ZN(II18990), .A(g9183) );
  INV_X1 NOT_3651( .ZN(g11812), .A(II18990) );
  INV_X1 NOT_3652( .ZN(g11813), .A(g11004) );
  INV_X1 NOT_3653( .ZN(g11817), .A(g11008) );
  INV_X1 NOT_3654( .ZN(g11818), .A(g11011) );
  INV_X1 NOT_3655( .ZN(g11819), .A(g11014) );
  INV_X1 NOT_3656( .ZN(g11820), .A(g11017) );
  INV_X1 NOT_3657( .ZN(g11821), .A(g10848) );
  INV_X1 NOT_3658( .ZN(g11824), .A(g11022) );
  INV_X1 NOT_3659( .ZN(g11825), .A(g11025) );
  INV_X1 NOT_3660( .ZN(g11826), .A(g11028) );
  INV_X1 NOT_3661( .ZN(g11827), .A(g11032) );
  INV_X1 NOT_3662( .ZN(g11829), .A(g11035) );
  INV_X1 NOT_3663( .ZN(g11834), .A(g11036) );
  INV_X1 NOT_3664( .ZN(g11835), .A(g11039) );
  INV_X1 NOT_3665( .ZN(g11836), .A(g11042) );
  INV_X1 NOT_3666( .ZN(g11837), .A(g11045) );
  INV_X1 NOT_3667( .ZN(g11841), .A(g11048) );
  INV_X1 NOT_3668( .ZN(g11842), .A(g11051) );
  INV_X1 NOT_3669( .ZN(II19025), .A(g9225) );
  INV_X1 NOT_3670( .ZN(g11845), .A(II19025) );
  INV_X1 NOT_3671( .ZN(g11846), .A(g11056) );
  INV_X1 NOT_3672( .ZN(II19030), .A(g8726) );
  INV_X2 NOT_3673( .ZN(g11848), .A(II19030) );
  INV_X2 NOT_3674( .ZN(g11852), .A(g11063) );
  INV_X2 NOT_3675( .ZN(g11853), .A(g11066) );
  INV_X2 NOT_3676( .ZN(g11854), .A(g11078) );
  INV_X1 NOT_3677( .ZN(g11856), .A(g11079) );
  INV_X1 NOT_3678( .ZN(g11857), .A(g11082) );
  INV_X1 NOT_3679( .ZN(g11858), .A(g11085) );
  INV_X1 NOT_3680( .ZN(g11859), .A(g11088) );
  INV_X1 NOT_3681( .ZN(g11862), .A(g11091) );
  INV_X1 NOT_3682( .ZN(g11866), .A(g11092) );
  INV_X1 NOT_3683( .ZN(g11867), .A(g11095) );
  INV_X1 NOT_3684( .ZN(g11868), .A(g11098) );
  INV_X1 NOT_3685( .ZN(g11869), .A(g11102) );
  INV_X1 NOT_3686( .ZN(g11871), .A(g11105) );
  INV_X1 NOT_3687( .ZN(g11876), .A(g11108) );
  INV_X1 NOT_3688( .ZN(g11877), .A(g11111) );
  INV_X1 NOT_3689( .ZN(g11878), .A(g11114) );
  INV_X1 NOT_3690( .ZN(g11879), .A(g11117) );
  INV_X1 NOT_3691( .ZN(g11883), .A(g11120) );
  INV_X1 NOT_3692( .ZN(g11884), .A(g11123) );
  INV_X1 NOT_3693( .ZN(g11886), .A(g11126) );
  INV_X1 NOT_3694( .ZN(g11887), .A(g11129) );
  INV_X1 NOT_3695( .ZN(g11888), .A(g11021) );
  INV_X1 NOT_3696( .ZN(g11891), .A(g11132) );
  INV_X1 NOT_3697( .ZN(g11892), .A(g11135) );
  INV_X1 NOT_3698( .ZN(g11893), .A(g11138) );
  INV_X1 NOT_3699( .ZN(g11894), .A(g11141) );
  INV_X1 NOT_3700( .ZN(g11895), .A(g11144) );
  INV_X1 NOT_3701( .ZN(g11898), .A(g11145) );
  INV_X1 NOT_3702( .ZN(g11899), .A(g11148) );
  INV_X1 NOT_3703( .ZN(g11900), .A(g11151) );
  INV_X1 NOT_3704( .ZN(g11901), .A(g11154) );
  INV_X1 NOT_3705( .ZN(g11904), .A(g11157) );
  INV_X1 NOT_3706( .ZN(g11908), .A(g11160) );
  INV_X1 NOT_3707( .ZN(g11909), .A(g11163) );
  INV_X1 NOT_3708( .ZN(g11910), .A(g11166) );
  INV_X1 NOT_3709( .ZN(g11911), .A(g11170) );
  INV_X1 NOT_3710( .ZN(g11913), .A(g11173) );
  INV_X1 NOT_3711( .ZN(g11918), .A(g11176) );
  INV_X1 NOT_3712( .ZN(g11919), .A(g11179) );
  INV_X1 NOT_3713( .ZN(g11920), .A(g11182) );
  INV_X1 NOT_3714( .ZN(g11921), .A(g11185) );
  INV_X1 NOT_3715( .ZN(II19105), .A(g8726) );
  INV_X1 NOT_3716( .ZN(g11923), .A(II19105) );
  INV_X1 NOT_3717( .ZN(g11927), .A(g10987) );
  INV_X1 NOT_3718( .ZN(g11929), .A(g11199) );
  INV_X1 NOT_3719( .ZN(g11930), .A(g11202) );
  INV_X1 NOT_3720( .ZN(g11931), .A(g11205) );
  INV_X1 NOT_3721( .ZN(g11932), .A(g11209) );
  INV_X1 NOT_3722( .ZN(g11933), .A(g11210) );
  INV_X1 NOT_3723( .ZN(g11936), .A(g11213) );
  INV_X1 NOT_3724( .ZN(II19119), .A(g9202) );
  INV_X1 NOT_3725( .ZN(g11937), .A(II19119) );
  INV_X1 NOT_3726( .ZN(g11941), .A(g11216) );
  INV_X1 NOT_3727( .ZN(g11942), .A(g11219) );
  INV_X1 NOT_3728( .ZN(g11943), .A(g11222) );
  INV_X1 NOT_3729( .ZN(g11944), .A(g11225) );
  INV_X1 NOT_3730( .ZN(g11945), .A(g11228) );
  INV_X1 NOT_3731( .ZN(g11948), .A(g11231) );
  INV_X1 NOT_3732( .ZN(g11949), .A(g11234) );
  INV_X1 NOT_3733( .ZN(g11950), .A(g11237) );
  INV_X1 NOT_3734( .ZN(g11951), .A(g11240) );
  INV_X1 NOT_3735( .ZN(g11954), .A(g11243) );
  INV_X1 NOT_3736( .ZN(g11958), .A(g11246) );
  INV_X1 NOT_3737( .ZN(g11959), .A(g11249) );
  INV_X1 NOT_3738( .ZN(g11960), .A(g11252) );
  INV_X1 NOT_3739( .ZN(g11961), .A(g11256) );
  INV_X1 NOT_3740( .ZN(g11963), .A(g11259) );
  INV_X1 NOT_3741( .ZN(g11968), .A(g11265) );
  INV_X1 NOT_3742( .ZN(g11969), .A(g11268) );
  INV_X1 NOT_3743( .ZN(g11970), .A(g11271) );
  INV_X1 NOT_3744( .ZN(g11971), .A(g11274) );
  INV_X1 NOT_3745( .ZN(g11972), .A(g11277) );
  INV_X1 NOT_3746( .ZN(g11973), .A(g11278) );
  INV_X1 NOT_3747( .ZN(II19160), .A(g10549) );
  INV_X1 NOT_3748( .ZN(g11976), .A(II19160) );
  INV_X1 NOT_3749( .ZN(g11982), .A(g11281) );
  INV_X1 NOT_3750( .ZN(g11983), .A(g11284) );
  INV_X1 NOT_3751( .ZN(g11984), .A(g11287) );
  INV_X1 NOT_3752( .ZN(g11985), .A(g11291) );
  INV_X1 NOT_3753( .ZN(g11986), .A(g11294) );
  INV_X1 NOT_3754( .ZN(g11989), .A(g11297) );
  INV_X1 NOT_3755( .ZN(II19174), .A(g9263) );
  INV_X1 NOT_3756( .ZN(g11990), .A(II19174) );
  INV_X1 NOT_3757( .ZN(g11994), .A(g11300) );
  INV_X1 NOT_3758( .ZN(g11995), .A(g11303) );
  INV_X1 NOT_3759( .ZN(g11996), .A(g11306) );
  INV_X1 NOT_3760( .ZN(g11997), .A(g11309) );
  INV_X1 NOT_3761( .ZN(g11998), .A(g11312) );
  INV_X1 NOT_3762( .ZN(g12001), .A(g11315) );
  INV_X1 NOT_3763( .ZN(g12002), .A(g11318) );
  INV_X1 NOT_3764( .ZN(g12003), .A(g11321) );
  INV_X1 NOT_3765( .ZN(g12004), .A(g11324) );
  INV_X1 NOT_3766( .ZN(g12007), .A(g11327) );
  INV_X1 NOT_3767( .ZN(II19195), .A(g8726) );
  INV_X1 NOT_3768( .ZN(g12009), .A(II19195) );
  INV_X1 NOT_3769( .ZN(g12013), .A(g10772) );
  INV_X1 NOT_3770( .ZN(g12017), .A(g10100) );
  INV_X1 NOT_3771( .ZN(g12020), .A(g11341) );
  INV_X1 NOT_3772( .ZN(g12021), .A(g11344) );
  INV_X1 NOT_3773( .ZN(g12022), .A(g11348) );
  INV_X1 NOT_3774( .ZN(g12023), .A(g11351) );
  INV_X1 NOT_3775( .ZN(g12024), .A(g11354) );
  INV_X1 NOT_3776( .ZN(g12025), .A(g11355) );
  INV_X1 NOT_3777( .ZN(II19208), .A(g10424) );
  INV_X1 NOT_3778( .ZN(g12027), .A(II19208) );
  INV_X1 NOT_3779( .ZN(II19211), .A(g10486) );
  INV_X1 NOT_3780( .ZN(g12030), .A(II19211) );
  INV_X1 NOT_3781( .ZN(g12037), .A(g11358) );
  INV_X1 NOT_3782( .ZN(g12038), .A(g11361) );
  INV_X1 NOT_3783( .ZN(g12039), .A(g11364) );
  INV_X1 NOT_3784( .ZN(g12040), .A(g11367) );
  INV_X1 NOT_3785( .ZN(g12041), .A(g11370) );
  INV_X1 NOT_3786( .ZN(g12042), .A(g11373) );
  INV_X1 NOT_3787( .ZN(II19226), .A(g10606) );
  INV_X1 NOT_3788( .ZN(g12045), .A(II19226) );
  INV_X1 NOT_3789( .ZN(g12051), .A(g11376) );
  INV_X1 NOT_3790( .ZN(g12052), .A(g11379) );
  INV_X1 NOT_3791( .ZN(g12053), .A(g11382) );
  INV_X1 NOT_3792( .ZN(g12054), .A(g11386) );
  INV_X1 NOT_3793( .ZN(g12055), .A(g11389) );
  INV_X1 NOT_3794( .ZN(g12058), .A(g11392) );
  INV_X1 NOT_3795( .ZN(II19240), .A(g9341) );
  INV_X1 NOT_3796( .ZN(g12059), .A(II19240) );
  INV_X1 NOT_3797( .ZN(g12063), .A(g11395) );
  INV_X1 NOT_3798( .ZN(g12064), .A(g11398) );
  INV_X1 NOT_3799( .ZN(g12065), .A(g11401) );
  INV_X1 NOT_3800( .ZN(g12066), .A(g11404) );
  INV_X1 NOT_3801( .ZN(g12067), .A(g11407) );
  INV_X1 NOT_3802( .ZN(g12071), .A(g10783) );
  INV_X1 NOT_3803( .ZN(g12075), .A(g11411) );
  INV_X1 NOT_3804( .ZN(g12076), .A(g11414) );
  INV_X1 NOT_3805( .ZN(g12077), .A(g11417) );
  INV_X1 NOT_3806( .ZN(g12078), .A(g11422) );
  INV_X1 NOT_3807( .ZN(g12084), .A(g11425) );
  INV_X1 NOT_3808( .ZN(g12085), .A(g11428) );
  INV_X1 NOT_3809( .ZN(g12086), .A(g11432) );
  INV_X1 NOT_3810( .ZN(g12087), .A(g11435) );
  INV_X1 NOT_3811( .ZN(g12088), .A(g11438) );
  INV_X1 NOT_3812( .ZN(g12089), .A(g11441) );
  INV_X1 NOT_3813( .ZN(II19271), .A(g10500) );
  INV_X1 NOT_3814( .ZN(g12091), .A(II19271) );
  INV_X1 NOT_3815( .ZN(II19274), .A(g10560) );
  INV_X1 NOT_3816( .ZN(g12094), .A(II19274) );
  INV_X1 NOT_3817( .ZN(g12101), .A(g11444) );
  INV_X1 NOT_3818( .ZN(g12102), .A(g11447) );
  INV_X1 NOT_3819( .ZN(g12103), .A(g11450) );
  INV_X1 NOT_3820( .ZN(g12104), .A(g11453) );
  INV_X1 NOT_3821( .ZN(g12105), .A(g11456) );
  INV_X1 NOT_3822( .ZN(g12106), .A(g11459) );
  INV_X1 NOT_3823( .ZN(II19289), .A(g10653) );
  INV_X1 NOT_3824( .ZN(g12109), .A(II19289) );
  INV_X1 NOT_3825( .ZN(g12115), .A(g11462) );
  INV_X1 NOT_3826( .ZN(g12116), .A(g11465) );
  INV_X1 NOT_3827( .ZN(g12117), .A(g11468) );
  INV_X1 NOT_3828( .ZN(g12118), .A(g11472) );
  INV_X1 NOT_3829( .ZN(g12119), .A(g11475) );
  INV_X1 NOT_3830( .ZN(g12122), .A(g11478) );
  INV_X1 NOT_3831( .ZN(II19303), .A(g9422) );
  INV_X1 NOT_3832( .ZN(g12123), .A(II19303) );
  INV_X1 NOT_3833( .ZN(II19307), .A(g8726) );
  INV_X1 NOT_3834( .ZN(g12125), .A(II19307) );
  INV_X1 NOT_3835( .ZN(g12130), .A(g10788) );
  INV_X1 NOT_3836( .ZN(g12134), .A(g8321) );
  INV_X1 NOT_3837( .ZN(g12135), .A(g8324) );
  INV_X1 NOT_3838( .ZN(II19315), .A(g10424) );
  INV_X1 NOT_3839( .ZN(g12136), .A(II19315) );
  INV_X1 NOT_3840( .ZN(II19318), .A(g10486) );
  INV_X1 NOT_3841( .ZN(g12139), .A(II19318) );
  INV_X1 NOT_3842( .ZN(II19321), .A(g10549) );
  INV_X1 NOT_3843( .ZN(g12142), .A(II19321) );
  INV_X1 NOT_3844( .ZN(g12147), .A(g8330) );
  INV_X1 NOT_3845( .ZN(g12148), .A(g8333) );
  INV_X1 NOT_3846( .ZN(g12149), .A(g8336) );
  INV_X1 NOT_3847( .ZN(g12150), .A(g8341) );
  INV_X1 NOT_3848( .ZN(g12156), .A(g8344) );
  INV_X1 NOT_3849( .ZN(g12157), .A(g8347) );
  INV_X1 NOT_3850( .ZN(g12158), .A(g8351) );
  INV_X1 NOT_3851( .ZN(g12159), .A(g8354) );
  INV_X1 NOT_3852( .ZN(g12160), .A(g8357) );
  INV_X1 NOT_3853( .ZN(g12161), .A(g8360) );
  INV_X1 NOT_3854( .ZN(II19342), .A(g10574) );
  INV_X1 NOT_3855( .ZN(g12163), .A(II19342) );
  INV_X1 NOT_3856( .ZN(II19345), .A(g10617) );
  INV_X1 NOT_3857( .ZN(g12166), .A(II19345) );
  INV_X1 NOT_3858( .ZN(g12173), .A(g8363) );
  INV_X1 NOT_3859( .ZN(g12174), .A(g8366) );
  INV_X2 NOT_3860( .ZN(g12175), .A(g8369) );
  INV_X2 NOT_3861( .ZN(g12176), .A(g8372) );
  INV_X2 NOT_3862( .ZN(g12177), .A(g8375) );
  INV_X1 NOT_3863( .ZN(g12178), .A(g8378) );
  INV_X1 NOT_3864( .ZN(II19360), .A(g10683) );
  INV_X1 NOT_3865( .ZN(g12181), .A(II19360) );
  INV_X1 NOT_3866( .ZN(g12187), .A(g8285) );
  INV_X1 NOT_3867( .ZN(g12191), .A(g8382) );
  INV_X1 NOT_3868( .ZN(g12196), .A(g8388) );
  INV_X1 NOT_3869( .ZN(g12197), .A(g8391) );
  INV_X1 NOT_3870( .ZN(II19374), .A(g10500) );
  INV_X1 NOT_3871( .ZN(g12198), .A(II19374) );
  INV_X1 NOT_3872( .ZN(II19377), .A(g10560) );
  INV_X1 NOT_3873( .ZN(g12201), .A(II19377) );
  INV_X1 NOT_3874( .ZN(II19380), .A(g10606) );
  INV_X1 NOT_3875( .ZN(g12204), .A(II19380) );
  INV_X1 NOT_3876( .ZN(g12209), .A(g8397) );
  INV_X1 NOT_3877( .ZN(g12210), .A(g8400) );
  INV_X1 NOT_3878( .ZN(g12211), .A(g8403) );
  INV_X1 NOT_3879( .ZN(g12212), .A(g8408) );
  INV_X1 NOT_3880( .ZN(g12218), .A(g8411) );
  INV_X1 NOT_3881( .ZN(g12219), .A(g8414) );
  INV_X1 NOT_3882( .ZN(g12220), .A(g8418) );
  INV_X1 NOT_3883( .ZN(g12221), .A(g8421) );
  INV_X1 NOT_3884( .ZN(g12222), .A(g8424) );
  INV_X1 NOT_3885( .ZN(g12223), .A(g8427) );
  INV_X1 NOT_3886( .ZN(II19401), .A(g10631) );
  INV_X1 NOT_3887( .ZN(g12225), .A(II19401) );
  INV_X1 NOT_3888( .ZN(II19404), .A(g10664) );
  INV_X1 NOT_3889( .ZN(g12228), .A(II19404) );
  INV_X1 NOT_3890( .ZN(g12235), .A(g8294) );
  INV_X1 NOT_3891( .ZN(II19412), .A(g10486) );
  INV_X1 NOT_3892( .ZN(g12239), .A(II19412) );
  INV_X1 NOT_3893( .ZN(II19415), .A(g10549) );
  INV_X1 NOT_3894( .ZN(g12242), .A(II19415) );
  INV_X1 NOT_3895( .ZN(g12246), .A(g8434) );
  INV_X1 NOT_3896( .ZN(g12251), .A(g8440) );
  INV_X1 NOT_3897( .ZN(g12252), .A(g8443) );
  INV_X1 NOT_3898( .ZN(II19426), .A(g10574) );
  INV_X1 NOT_3899( .ZN(g12253), .A(II19426) );
  INV_X1 NOT_3900( .ZN(II19429), .A(g10617) );
  INV_X1 NOT_3901( .ZN(g12256), .A(II19429) );
  INV_X1 NOT_3902( .ZN(II19432), .A(g10653) );
  INV_X1 NOT_3903( .ZN(g12259), .A(II19432) );
  INV_X1 NOT_3904( .ZN(g12264), .A(g8449) );
  INV_X1 NOT_3905( .ZN(g12265), .A(g8452) );
  INV_X1 NOT_3906( .ZN(g12266), .A(g8455) );
  INV_X1 NOT_3907( .ZN(g12267), .A(g8460) );
  INV_X1 NOT_3908( .ZN(g12275), .A(g8303) );
  INV_X1 NOT_3909( .ZN(II19449), .A(g10424) );
  INV_X1 NOT_3910( .ZN(g12279), .A(II19449) );
  INV_X1 NOT_3911( .ZN(II19452), .A(g10560) );
  INV_X1 NOT_3912( .ZN(g12282), .A(II19452) );
  INV_X1 NOT_3913( .ZN(II19455), .A(g10606) );
  INV_X1 NOT_3914( .ZN(g12285), .A(II19455) );
  INV_X1 NOT_3915( .ZN(g12289), .A(g8469) );
  INV_X1 NOT_3916( .ZN(g12294), .A(g8475) );
  INV_X1 NOT_3917( .ZN(g12295), .A(g8478) );
  INV_X1 NOT_3918( .ZN(II19466), .A(g10631) );
  INV_X1 NOT_3919( .ZN(g12296), .A(II19466) );
  INV_X1 NOT_3920( .ZN(II19469), .A(g10664) );
  INV_X1 NOT_3921( .ZN(g12299), .A(II19469) );
  INV_X1 NOT_3922( .ZN(II19472), .A(g10683) );
  INV_X1 NOT_3923( .ZN(g12302), .A(II19472) );
  INV_X1 NOT_3924( .ZN(g12308), .A(g8312) );
  INV_X1 NOT_3925( .ZN(II19479), .A(g10549) );
  INV_X1 NOT_3926( .ZN(g12312), .A(II19479) );
  INV_X1 NOT_3927( .ZN(II19482), .A(g10500) );
  INV_X1 NOT_3928( .ZN(g12315), .A(II19482) );
  INV_X1 NOT_3929( .ZN(II19485), .A(g10617) );
  INV_X1 NOT_3930( .ZN(g12318), .A(II19485) );
  INV_X1 NOT_3931( .ZN(II19488), .A(g10653) );
  INV_X1 NOT_3932( .ZN(g12321), .A(II19488) );
  INV_X1 NOT_3933( .ZN(g12325), .A(g8494) );
  INV_X1 NOT_3934( .ZN(g12332), .A(g10829) );
  INV_X1 NOT_3935( .ZN(II19500), .A(g10424) );
  INV_X1 NOT_3936( .ZN(g12333), .A(II19500) );
  INV_X1 NOT_3937( .ZN(II19503), .A(g10486) );
  INV_X1 NOT_3938( .ZN(g12336), .A(II19503) );
  INV_X1 NOT_3939( .ZN(II19507), .A(g10606) );
  INV_X1 NOT_3940( .ZN(g12340), .A(II19507) );
  INV_X1 NOT_3941( .ZN(II19510), .A(g10574) );
  INV_X1 NOT_3942( .ZN(g12343), .A(II19510) );
  INV_X1 NOT_3943( .ZN(II19513), .A(g10664) );
  INV_X1 NOT_3944( .ZN(g12346), .A(II19513) );
  INV_X1 NOT_3945( .ZN(II19516), .A(g10683) );
  INV_X1 NOT_3946( .ZN(g12349), .A(II19516) );
  INV_X1 NOT_3947( .ZN(g12354), .A(g8381) );
  INV_X1 NOT_3948( .ZN(g12362), .A(g10866) );
  INV_X1 NOT_3949( .ZN(II19523), .A(g10500) );
  INV_X1 NOT_3950( .ZN(g12363), .A(II19523) );
  INV_X1 NOT_3951( .ZN(II19526), .A(g10560) );
  INV_X1 NOT_3952( .ZN(g12366), .A(II19526) );
  INV_X1 NOT_3953( .ZN(II19530), .A(g10653) );
  INV_X1 NOT_3954( .ZN(g12370), .A(II19530) );
  INV_X1 NOT_3955( .ZN(II19533), .A(g10631) );
  INV_X1 NOT_3956( .ZN(g12373), .A(II19533) );
  INV_X1 NOT_3957( .ZN(g12378), .A(g10847) );
  INV_X1 NOT_3958( .ZN(II19539), .A(g10549) );
  INV_X1 NOT_3959( .ZN(g12379), .A(II19539) );
  INV_X1 NOT_3960( .ZN(II19542), .A(g10574) );
  INV_X1 NOT_3961( .ZN(g12382), .A(II19542) );
  INV_X1 NOT_3962( .ZN(II19545), .A(g10617) );
  INV_X1 NOT_3963( .ZN(g12385), .A(II19545) );
  INV_X1 NOT_3964( .ZN(II19549), .A(g10683) );
  INV_X1 NOT_3965( .ZN(g12389), .A(II19549) );
  INV_X1 NOT_3966( .ZN(II19552), .A(g8430) );
  INV_X1 NOT_3967( .ZN(g12392), .A(II19552) );
  INV_X1 NOT_3968( .ZN(g12408), .A(g11020) );
  INV_X1 NOT_3969( .ZN(II19557), .A(g10606) );
  INV_X1 NOT_3970( .ZN(g12409), .A(II19557) );
  INV_X1 NOT_3971( .ZN(II19560), .A(g10631) );
  INV_X1 NOT_3972( .ZN(g12412), .A(II19560) );
  INV_X1 NOT_3973( .ZN(II19563), .A(g10664) );
  INV_X1 NOT_3974( .ZN(g12415), .A(II19563) );
  INV_X1 NOT_3975( .ZN(g12420), .A(g10986) );
  INV_X1 NOT_3976( .ZN(II19569), .A(g10653) );
  INV_X1 NOT_3977( .ZN(g12421), .A(II19569) );
  INV_X1 NOT_3978( .ZN(g12424), .A(g10962) );
  INV_X1 NOT_3979( .ZN(II19573), .A(g8835) );
  INV_X1 NOT_3980( .ZN(g12425), .A(II19573) );
  INV_X1 NOT_3981( .ZN(II19576), .A(g10683) );
  INV_X1 NOT_3982( .ZN(g12426), .A(II19576) );
  INV_X1 NOT_3983( .ZN(g12430), .A(g10905) );
  INV_X1 NOT_3984( .ZN(II19582), .A(g8862) );
  INV_X1 NOT_3985( .ZN(g12432), .A(II19582) );
  INV_X1 NOT_3986( .ZN(g12434), .A(g10929) );
  INV_X1 NOT_3987( .ZN(II19587), .A(g9173) );
  INV_X1 NOT_3988( .ZN(g12435), .A(II19587) );
  INV_X1 NOT_3989( .ZN(II19591), .A(g8900) );
  INV_X1 NOT_3990( .ZN(g12437), .A(II19591) );
  INV_X1 NOT_3991( .ZN(g12438), .A(g10846) );
  INV_X1 NOT_3992( .ZN(II19595), .A(g10810) );
  INV_X1 NOT_3993( .ZN(g12439), .A(II19595) );
  INV_X1 NOT_3994( .ZN(II19598), .A(g9215) );
  INV_X1 NOT_3995( .ZN(g12440), .A(II19598) );
  INV_X1 NOT_3996( .ZN(II19602), .A(g8940) );
  INV_X1 NOT_3997( .ZN(g12442), .A(II19602) );
  INV_X1 NOT_3998( .ZN(II19605), .A(g10797) );
  INV_X1 NOT_3999( .ZN(g12443), .A(II19605) );
  INV_X1 NOT_4000( .ZN(II19608), .A(g10831) );
  INV_X1 NOT_4001( .ZN(g12444), .A(II19608) );
  INV_X1 NOT_4002( .ZN(II19611), .A(g9276) );
  INV_X1 NOT_4003( .ZN(g12445), .A(II19611) );
  INV_X1 NOT_4004( .ZN(II19615), .A(g10789) );
  INV_X1 NOT_4005( .ZN(g12447), .A(II19615) );
  INV_X1 NOT_4006( .ZN(II19618), .A(g10814) );
  INV_X1 NOT_4007( .ZN(g12448), .A(II19618) );
  INV_X1 NOT_4008( .ZN(II19621), .A(g10851) );
  INV_X1 NOT_4009( .ZN(g12449), .A(II19621) );
  INV_X1 NOT_4010( .ZN(II19624), .A(g9354) );
  INV_X1 NOT_4011( .ZN(g12450), .A(II19624) );
  INV_X1 NOT_4012( .ZN(II19628), .A(g10784) );
  INV_X1 NOT_4013( .ZN(g12452), .A(II19628) );
  INV_X1 NOT_4014( .ZN(II19631), .A(g10801) );
  INV_X1 NOT_4015( .ZN(g12453), .A(II19631) );
  INV_X1 NOT_4016( .ZN(II19634), .A(g10835) );
  INV_X1 NOT_4017( .ZN(g12454), .A(II19634) );
  INV_X1 NOT_4018( .ZN(II19637), .A(g10872) );
  INV_X1 NOT_4019( .ZN(g12455), .A(II19637) );
  INV_X1 NOT_4020( .ZN(g12456), .A(g8602) );
  INV_X1 NOT_4021( .ZN(II19642), .A(g10793) );
  INV_X1 NOT_4022( .ZN(g12460), .A(II19642) );
  INV_X1 NOT_4023( .ZN(II19645), .A(g10818) );
  INV_X1 NOT_4024( .ZN(g12461), .A(II19645) );
  INV_X1 NOT_4025( .ZN(II19648), .A(g10855) );
  INV_X2 NOT_4026( .ZN(g12462), .A(II19648) );
  INV_X2 NOT_4027( .ZN(g12463), .A(g10730) );
  INV_X2 NOT_4028( .ZN(g12466), .A(g8614) );
  INV_X2 NOT_4029( .ZN(II19654), .A(g10805) );
  INV_X1 NOT_4030( .ZN(g12470), .A(II19654) );
  INV_X1 NOT_4031( .ZN(II19657), .A(g10839) );
  INV_X1 NOT_4032( .ZN(g12471), .A(II19657) );
  INV_X1 NOT_4033( .ZN(g12472), .A(g8617) );
  INV_X1 NOT_4034( .ZN(g12473), .A(g8580) );
  INV_X1 NOT_4035( .ZN(g12476), .A(g8622) );
  INV_X1 NOT_4036( .ZN(g12478), .A(g10749) );
  INV_X1 NOT_4037( .ZN(g12481), .A(g8627) );
  INV_X1 NOT_4038( .ZN(II19667), .A(g10822) );
  INV_X1 NOT_4039( .ZN(g12485), .A(II19667) );
  INV_X1 NOT_4040( .ZN(g12490), .A(g8587) );
  INV_X1 NOT_4041( .ZN(g12493), .A(g8632) );
  INV_X1 NOT_4042( .ZN(g12495), .A(g10767) );
  INV_X1 NOT_4043( .ZN(g12498), .A(g8637) );
  INV_X1 NOT_4044( .ZN(g12502), .A(g8640) );
  INV_X1 NOT_4045( .ZN(g12504), .A(g8643) );
  INV_X1 NOT_4046( .ZN(g12505), .A(g8646) );
  INV_X1 NOT_4047( .ZN(g12510), .A(g8594) );
  INV_X1 NOT_4048( .ZN(g12513), .A(g8651) );
  INV_X1 NOT_4049( .ZN(g12515), .A(g10773) );
  INV_X1 NOT_4050( .ZN(g12518), .A(g8655) );
  INV_X1 NOT_4051( .ZN(II19689), .A(g10016) );
  INV_X1 NOT_4052( .ZN(g12519), .A(II19689) );
  INV_X1 NOT_4053( .ZN(g12521), .A(g8659) );
  INV_X1 NOT_4054( .ZN(g12522), .A(g8662) );
  INV_X1 NOT_4055( .ZN(g12527), .A(g8605) );
  INV_X1 NOT_4056( .ZN(g12530), .A(g8667) );
  INV_X1 NOT_4057( .ZN(g12532), .A(g8670) );
  INV_X1 NOT_4058( .ZN(g12533), .A(g8673) );
  INV_X1 NOT_4059( .ZN(II19702), .A(g10125) );
  INV_X1 NOT_4060( .ZN(g12534), .A(II19702) );
  INV_X1 NOT_4061( .ZN(g12536), .A(g8678) );
  INV_X1 NOT_4062( .ZN(g12537), .A(g8681) );
  INV_X1 NOT_4063( .ZN(g12542), .A(g8684) );
  INV_X1 NOT_4064( .ZN(II19711), .A(g10230) );
  INV_X1 NOT_4065( .ZN(g12543), .A(II19711) );
  INV_X1 NOT_4066( .ZN(g12545), .A(g8690) );
  INV_X1 NOT_4067( .ZN(g12546), .A(g8693) );
  INV_X1 NOT_4068( .ZN(g12547), .A(g8696) );
  INV_X1 NOT_4069( .ZN(II19718), .A(g8726) );
  INV_X1 NOT_4070( .ZN(g12548), .A(II19718) );
  INV_X1 NOT_4071( .ZN(g12551), .A(g8700) );
  INV_X1 NOT_4072( .ZN(II19722), .A(g10332) );
  INV_X1 NOT_4073( .ZN(g12552), .A(II19722) );
  INV_X1 NOT_4074( .ZN(g12553), .A(g8708) );
  INV_X1 NOT_4075( .ZN(g12554), .A(g8711) );
  INV_X1 NOT_4076( .ZN(II19727), .A(g8726) );
  INV_X1 NOT_4077( .ZN(g12555), .A(II19727) );
  INV_X1 NOT_4078( .ZN(g12558), .A(g8714) );
  INV_X1 NOT_4079( .ZN(g12559), .A(g8719) );
  INV_X1 NOT_4080( .ZN(g12560), .A(g8745) );
  INV_X1 NOT_4081( .ZN(II19733), .A(g8726) );
  INV_X1 NOT_4082( .ZN(g12561), .A(II19733) );
  INV_X1 NOT_4083( .ZN(II19736), .A(g9184) );
  INV_X1 NOT_4084( .ZN(g12564), .A(II19736) );
  INV_X1 NOT_4085( .ZN(II19739), .A(g10694) );
  INV_X1 NOT_4086( .ZN(g12565), .A(II19739) );
  INV_X1 NOT_4087( .ZN(g12596), .A(g8748) );
  INV_X1 NOT_4088( .ZN(g12597), .A(g8752) );
  INV_X1 NOT_4089( .ZN(g12598), .A(g8757) );
  INV_X1 NOT_4090( .ZN(g12599), .A(g8763) );
  INV_X1 NOT_4091( .ZN(g12600), .A(g8766) );
  INV_X1 NOT_4092( .ZN(II19747), .A(g8726) );
  INV_X1 NOT_4093( .ZN(g12601), .A(II19747) );
  INV_X1 NOT_4094( .ZN(II19750), .A(g8726) );
  INV_X1 NOT_4095( .ZN(g12604), .A(II19750) );
  INV_X1 NOT_4096( .ZN(II19753), .A(g9229) );
  INV_X1 NOT_4097( .ZN(g12607), .A(II19753) );
  INV_X1 NOT_4098( .ZN(II19756), .A(g10424) );
  INV_X1 NOT_4099( .ZN(g12608), .A(II19756) );
  INV_X1 NOT_4100( .ZN(II19759), .A(g10714) );
  INV_X1 NOT_4101( .ZN(g12611), .A(II19759) );
  INV_X1 NOT_4102( .ZN(g12642), .A(g8771) );
  INV_X1 NOT_4103( .ZN(g12643), .A(g8775) );
  INV_X1 NOT_4104( .ZN(g12644), .A(g8780) );
  INV_X1 NOT_4105( .ZN(g12645), .A(g8785) );
  INV_X1 NOT_4106( .ZN(g12646), .A(g8788) );
  INV_X1 NOT_4107( .ZN(II19767), .A(g8726) );
  INV_X1 NOT_4108( .ZN(g12647), .A(II19767) );
  INV_X1 NOT_4109( .ZN(II19771), .A(g10038) );
  INV_X1 NOT_4110( .ZN(g12651), .A(II19771) );
  INV_X1 NOT_4111( .ZN(II19774), .A(g10500) );
  INV_X1 NOT_4112( .ZN(g12654), .A(II19774) );
  INV_X1 NOT_4113( .ZN(II19777), .A(g10735) );
  INV_X1 NOT_4114( .ZN(g12657), .A(II19777) );
  INV_X1 NOT_4115( .ZN(g12688), .A(g8794) );
  INV_X1 NOT_4116( .ZN(g12689), .A(g8798) );
  INV_X1 NOT_4117( .ZN(g12690), .A(g8802) );
  INV_X1 NOT_4118( .ZN(g12691), .A(g8805) );
  INV_X1 NOT_4119( .ZN(II19784), .A(g8726) );
  INV_X1 NOT_4120( .ZN(g12692), .A(II19784) );
  INV_X1 NOT_4121( .ZN(II19787), .A(g8726) );
  INV_X1 NOT_4122( .ZN(g12695), .A(II19787) );
  INV_X1 NOT_4123( .ZN(II19791), .A(g10486) );
  INV_X1 NOT_4124( .ZN(g12699), .A(II19791) );
  INV_X1 NOT_4125( .ZN(II19794), .A(g10676) );
  INV_X1 NOT_4126( .ZN(g12702), .A(II19794) );
  INV_X1 NOT_4127( .ZN(II19797), .A(g10147) );
  INV_X1 NOT_4128( .ZN(g12705), .A(II19797) );
  INV_X1 NOT_4129( .ZN(II19800), .A(g10574) );
  INV_X1 NOT_4130( .ZN(g12708), .A(II19800) );
  INV_X1 NOT_4131( .ZN(II19803), .A(g10754) );
  INV_X1 NOT_4132( .ZN(g12711), .A(II19803) );
  INV_X1 NOT_4133( .ZN(g12742), .A(g8813) );
  INV_X1 NOT_4134( .ZN(g12743), .A(g8817) );
  INV_X1 NOT_4135( .ZN(II19808), .A(g8726) );
  INV_X1 NOT_4136( .ZN(g12744), .A(II19808) );
  INV_X1 NOT_4137( .ZN(g12748), .A(g8823) );
  INV_X1 NOT_4138( .ZN(II19813), .A(g10649) );
  INV_X1 NOT_4139( .ZN(g12749), .A(II19813) );
  INV_X1 NOT_4140( .ZN(II19816), .A(g10703) );
  INV_X1 NOT_4141( .ZN(g12752), .A(II19816) );
  INV_X1 NOT_4142( .ZN(II19820), .A(g10560) );
  INV_X1 NOT_4143( .ZN(g12756), .A(II19820) );
  INV_X1 NOT_4144( .ZN(II19823), .A(g10705) );
  INV_X1 NOT_4145( .ZN(g12759), .A(II19823) );
  INV_X1 NOT_4146( .ZN(II19826), .A(g10252) );
  INV_X1 NOT_4147( .ZN(g12762), .A(II19826) );
  INV_X1 NOT_4148( .ZN(II19829), .A(g10631) );
  INV_X1 NOT_4149( .ZN(g12765), .A(II19829) );
  INV_X1 NOT_4150( .ZN(g12768), .A(g8829) );
  INV_X1 NOT_4151( .ZN(II19833), .A(g8726) );
  INV_X1 NOT_4152( .ZN(g12769), .A(II19833) );
  INV_X1 NOT_4153( .ZN(II19836), .A(g8726) );
  INV_X1 NOT_4154( .ZN(g12772), .A(II19836) );
  INV_X1 NOT_4155( .ZN(g12775), .A(g8832) );
  INV_X1 NOT_4156( .ZN(g12776), .A(g10766) );
  INV_X1 NOT_4157( .ZN(g12782), .A(g8836) );
  INV_X1 NOT_4158( .ZN(II19844), .A(g8533) );
  INV_X1 NOT_4159( .ZN(g12783), .A(II19844) );
  INV_X1 NOT_4160( .ZN(II19847), .A(g10677) );
  INV_X1 NOT_4161( .ZN(g12786), .A(II19847) );
  INV_X1 NOT_4162( .ZN(g12790), .A(g8847) );
  INV_X1 NOT_4163( .ZN(II19852), .A(g10679) );
  INV_X1 NOT_4164( .ZN(g12791), .A(II19852) );
  INV_X1 NOT_4165( .ZN(II19855), .A(g10723) );
  INV_X1 NOT_4166( .ZN(g12794), .A(II19855) );
  INV_X1 NOT_4167( .ZN(II19859), .A(g10617) );
  INV_X1 NOT_4168( .ZN(g12798), .A(II19859) );
  INV_X1 NOT_4169( .ZN(II19862), .A(g10725) );
  INV_X1 NOT_4170( .ZN(g12801), .A(II19862) );
  INV_X1 NOT_4171( .ZN(II19865), .A(g10354) );
  INV_X1 NOT_4172( .ZN(g12804), .A(II19865) );
  INV_X1 NOT_4173( .ZN(g12807), .A(g8853) );
  INV_X1 NOT_4174( .ZN(II19869), .A(g8726) );
  INV_X1 NOT_4175( .ZN(g12808), .A(II19869) );
  INV_X1 NOT_4176( .ZN(II19872), .A(g8317) );
  INV_X1 NOT_4177( .ZN(g12811), .A(II19872) );
  INV_X1 NOT_4178( .ZN(g12815), .A(g8856) );
  INV_X1 NOT_4179( .ZN(II19877), .A(g8547) );
  INV_X1 NOT_4180( .ZN(g12816), .A(II19877) );
  INV_X1 NOT_4181( .ZN(g12821), .A(g8863) );
  INV_X1 NOT_4182( .ZN(II19883), .A(g8550) );
  INV_X1 NOT_4183( .ZN(g12822), .A(II19883) );
  INV_X1 NOT_4184( .ZN(II19886), .A(g10706) );
  INV_X1 NOT_4185( .ZN(g12825), .A(II19886) );
  INV_X1 NOT_4186( .ZN(g12829), .A(g8874) );
  INV_X1 NOT_4187( .ZN(II19891), .A(g10708) );
  INV_X1 NOT_4188( .ZN(g12830), .A(II19891) );
  INV_X1 NOT_4189( .ZN(II19894), .A(g10744) );
  INV_X1 NOT_4190( .ZN(g12833), .A(II19894) );
  INV_X1 NOT_4191( .ZN(II19898), .A(g10664) );
  INV_X1 NOT_4192( .ZN(g12837), .A(II19898) );
  INV_X1 NOT_4193( .ZN(II19901), .A(g10746) );
  INV_X1 NOT_4194( .ZN(g12840), .A(II19901) );
  INV_X1 NOT_4195( .ZN(g12843), .A(g8879) );
  INV_X1 NOT_4196( .ZN(II19905), .A(g8726) );
  INV_X1 NOT_4197( .ZN(g12844), .A(II19905) );
  INV_X1 NOT_4198( .ZN(g12847), .A(g8882) );
  INV_X1 NOT_4199( .ZN(g12848), .A(g11059) );
  INV_X1 NOT_4200( .ZN(g12850), .A(g8885) );
  INV_X1 NOT_4201( .ZN(g12851), .A(g8888) );
  INV_X1 NOT_4202( .ZN(g12853), .A(g8894) );
  INV_X1 NOT_4203( .ZN(II19915), .A(g8560) );
  INV_X1 NOT_4204( .ZN(g12854), .A(II19915) );
  INV_X2 NOT_4205( .ZN(g12859), .A(g8901) );
  INV_X2 NOT_4206( .ZN(II19921), .A(g8563) );
  INV_X2 NOT_4207( .ZN(g12860), .A(II19921) );
  INV_X2 NOT_4208( .ZN(II19924), .A(g10726) );
  INV_X1 NOT_4209( .ZN(g12863), .A(II19924) );
  INV_X1 NOT_4210( .ZN(g12867), .A(g8912) );
  INV_X1 NOT_4211( .ZN(II19929), .A(g10728) );
  INV_X1 NOT_4212( .ZN(g12868), .A(II19929) );
  INV_X1 NOT_4213( .ZN(II19932), .A(g10763) );
  INV_X1 NOT_4214( .ZN(g12871), .A(II19932) );
  INV_X1 NOT_4215( .ZN(g12874), .A(g8915) );
  INV_X1 NOT_4216( .ZN(g12875), .A(g10779) );
  INV_X1 NOT_4217( .ZN(g12881), .A(g8918) );
  INV_X1 NOT_4218( .ZN(g12882), .A(g8921) );
  INV_X1 NOT_4219( .ZN(g12891), .A(g8925) );
  INV_X1 NOT_4220( .ZN(g12892), .A(g8928) );
  INV_X1 NOT_4221( .ZN(g12894), .A(g8934) );
  INV_X1 NOT_4222( .ZN(II19952), .A(g8571) );
  INV_X1 NOT_4223( .ZN(g12895), .A(II19952) );
  INV_X1 NOT_4224( .ZN(g12900), .A(g8941) );
  INV_X1 NOT_4225( .ZN(II19958), .A(g8574) );
  INV_X1 NOT_4226( .ZN(g12901), .A(II19958) );
  INV_X1 NOT_4227( .ZN(II19961), .A(g10747) );
  INV_X1 NOT_4228( .ZN(g12904), .A(II19961) );
  INV_X1 NOT_4229( .ZN(g12907), .A(g8949) );
  INV_X1 NOT_4230( .ZN(g12909), .A(g10904) );
  INV_X1 NOT_4231( .ZN(g12914), .A(g8952) );
  INV_X1 NOT_4232( .ZN(g12915), .A(g8955) );
  INV_X1 NOT_4233( .ZN(g12921), .A(g8958) );
  INV_X1 NOT_4234( .ZN(g12922), .A(g8961) );
  INV_X1 NOT_4235( .ZN(g12931), .A(g8965) );
  INV_X1 NOT_4236( .ZN(g12932), .A(g8968) );
  INV_X1 NOT_4237( .ZN(g12934), .A(g8974) );
  INV_X1 NOT_4238( .ZN(II19986), .A(g8577) );
  INV_X1 NOT_4239( .ZN(g12935), .A(II19986) );
  INV_X1 NOT_4240( .ZN(g12940), .A(g8980) );
  INV_X1 NOT_4241( .ZN(g12943), .A(g8984) );
  INV_X1 NOT_4242( .ZN(g12944), .A(g8987) );
  INV_X1 NOT_4243( .ZN(g12950), .A(g8990) );
  INV_X1 NOT_4244( .ZN(g12951), .A(g8993) );
  INV_X1 NOT_4245( .ZN(g12960), .A(g8997) );
  INV_X1 NOT_4246( .ZN(g12961), .A(g9000) );
  INV_X1 NOT_4247( .ZN(II20009), .A(g8313) );
  INV_X1 NOT_4248( .ZN(g12962), .A(II20009) );
  INV_X1 NOT_4249( .ZN(g12965), .A(g9006) );
  INV_X1 NOT_4250( .ZN(g12969), .A(g9010) );
  INV_X1 NOT_4251( .ZN(g12972), .A(g9013) );
  INV_X1 NOT_4252( .ZN(g12973), .A(g9016) );
  INV_X1 NOT_4253( .ZN(g12979), .A(g9019) );
  INV_X1 NOT_4254( .ZN(g12980), .A(g9022) );
  INV_X1 NOT_4255( .ZN(g12993), .A(g9035) );
  INV_X1 NOT_4256( .ZN(g12996), .A(g9038) );
  INV_X1 NOT_4257( .ZN(g12997), .A(g9041) );
  INV_X1 NOT_4258( .ZN(g12998), .A(g9044) );
  INV_X1 NOT_4259( .ZN(g13003), .A(g9058) );
  INV_X1 NOT_4260( .ZN(II20062), .A(g10480) );
  INV_X1 NOT_4261( .ZN(g13011), .A(II20062) );
  INV_X1 NOT_4262( .ZN(g13025), .A(g10810) );
  INV_X1 NOT_4263( .ZN(g13033), .A(g10797) );
  INV_X1 NOT_4264( .ZN(g13036), .A(g10831) );
  INV_X1 NOT_4265( .ZN(g13043), .A(g10789) );
  INV_X1 NOT_4266( .ZN(g13046), .A(g10814) );
  INV_X1 NOT_4267( .ZN(g13049), .A(g10851) );
  INV_X1 NOT_4268( .ZN(g13057), .A(g10784) );
  INV_X1 NOT_4269( .ZN(g13060), .A(g10801) );
  INV_X1 NOT_4270( .ZN(g13063), .A(g10835) );
  INV_X1 NOT_4271( .ZN(g13066), .A(g10872) );
  INV_X1 NOT_4272( .ZN(II20117), .A(g10876) );
  INV_X1 NOT_4273( .ZN(g13070), .A(II20117) );
  INV_X1 NOT_4274( .ZN(g13073), .A(g10793) );
  INV_X1 NOT_4275( .ZN(g13076), .A(g10818) );
  INV_X1 NOT_4276( .ZN(g13079), .A(g10855) );
  INV_X1 NOT_4277( .ZN(g13092), .A(g10805) );
  INV_X1 NOT_4278( .ZN(g13095), .A(g10839) );
  INV_X1 NOT_4279( .ZN(g13101), .A(g9128) );
  INV_X1 NOT_4280( .ZN(g13107), .A(g10822) );
  INV_X1 NOT_4281( .ZN(g13117), .A(g9134) );
  INV_X1 NOT_4282( .ZN(g13130), .A(g9140) );
  INV_X1 NOT_4283( .ZN(g13141), .A(g9146) );
  INV_X1 NOT_4284( .ZN(g13148), .A(g9170) );
  INV_X1 NOT_4285( .ZN(g13151), .A(g9184) );
  INV_X1 NOT_4286( .ZN(g13152), .A(g9196) );
  INV_X1 NOT_4287( .ZN(g13153), .A(g9199) );
  INV_X1 NOT_4288( .ZN(g13154), .A(g9212) );
  INV_X1 NOT_4289( .ZN(g13157), .A(g9229) );
  INV_X1 NOT_4290( .ZN(g13158), .A(g9242) );
  INV_X1 NOT_4291( .ZN(g13159), .A(g9245) );
  INV_X1 NOT_4292( .ZN(g13161), .A(g9257) );
  INV_X1 NOT_4293( .ZN(g13162), .A(g9260) );
  INV_X1 NOT_4294( .ZN(g13163), .A(g9273) );
  INV_X1 NOT_4295( .ZN(g13166), .A(g9290) );
  INV_X1 NOT_4296( .ZN(g13167), .A(g9303) );
  INV_X1 NOT_4297( .ZN(g13168), .A(g9306) );
  INV_X1 NOT_4298( .ZN(g13169), .A(g9320) );
  INV_X1 NOT_4299( .ZN(g13170), .A(g9323) );
  INV_X1 NOT_4300( .ZN(g13172), .A(g9335) );
  INV_X1 NOT_4301( .ZN(g13173), .A(g9338) );
  INV_X1 NOT_4302( .ZN(g13174), .A(g9351) );
  INV_X1 NOT_4303( .ZN(g13176), .A(g9368) );
  INV_X1 NOT_4304( .ZN(g13177), .A(g9371) );
  INV_X1 NOT_4305( .ZN(g13178), .A(g9384) );
  INV_X1 NOT_4306( .ZN(g13179), .A(g9387) );
  INV_X1 NOT_4307( .ZN(g13180), .A(g9401) );
  INV_X1 NOT_4308( .ZN(g13181), .A(g9404) );
  INV_X1 NOT_4309( .ZN(g13183), .A(g9416) );
  INV_X1 NOT_4310( .ZN(g13184), .A(g9419) );
  INV_X1 NOT_4311( .ZN(g13185), .A(g9443) );
  INV_X1 NOT_4312( .ZN(g13186), .A(g9446) );
  INV_X1 NOT_4313( .ZN(g13187), .A(g9450) );
  INV_X1 NOT_4314( .ZN(g13188), .A(g9465) );
  INV_X1 NOT_4315( .ZN(g13189), .A(g9468) );
  INV_X1 NOT_4316( .ZN(g13190), .A(g9481) );
  INV_X1 NOT_4317( .ZN(g13191), .A(g9484) );
  INV_X1 NOT_4318( .ZN(g13192), .A(g9498) );
  INV_X1 NOT_4319( .ZN(g13193), .A(g9501) );
  INV_X1 NOT_4320( .ZN(g13195), .A(g9524) );
  INV_X1 NOT_4321( .ZN(g13196), .A(g9528) );
  INV_X1 NOT_4322( .ZN(g13197), .A(g9531) );
  INV_X1 NOT_4323( .ZN(g13198), .A(g9585) );
  INV_X1 NOT_4324( .ZN(g13199), .A(g9588) );
  INV_X1 NOT_4325( .ZN(g13200), .A(g9592) );
  INV_X1 NOT_4326( .ZN(g13201), .A(g9607) );
  INV_X1 NOT_4327( .ZN(g13202), .A(g9610) );
  INV_X1 NOT_4328( .ZN(g13203), .A(g9623) );
  INV_X1 NOT_4329( .ZN(g13204), .A(g9626) );
  INV_X1 NOT_4330( .ZN(g13205), .A(g9641) );
  INV_X1 NOT_4331( .ZN(g13206), .A(g9644) );
  INV_X1 NOT_4332( .ZN(g13207), .A(g9666) );
  INV_X1 NOT_4333( .ZN(g13208), .A(g9670) );
  INV_X1 NOT_4334( .ZN(g13209), .A(g9673) );
  INV_X1 NOT_4335( .ZN(g13210), .A(g9727) );
  INV_X1 NOT_4336( .ZN(g13211), .A(g9730) );
  INV_X1 NOT_4337( .ZN(g13212), .A(g9734) );
  INV_X1 NOT_4338( .ZN(g13213), .A(g9749) );
  INV_X1 NOT_4339( .ZN(g13214), .A(g9752) );
  INV_X1 NOT_4340( .ZN(II20264), .A(g9027) );
  INV_X1 NOT_4341( .ZN(g13215), .A(II20264) );
  INV_X1 NOT_4342( .ZN(g13218), .A(g9767) );
  INV_X1 NOT_4343( .ZN(g13219), .A(g9770) );
  INV_X1 NOT_4344( .ZN(g13220), .A(g9787) );
  INV_X1 NOT_4345( .ZN(g13221), .A(g9790) );
  INV_X1 NOT_4346( .ZN(g13222), .A(g9812) );
  INV_X1 NOT_4347( .ZN(g13223), .A(g9816) );
  INV_X1 NOT_4348( .ZN(g13224), .A(g9819) );
  INV_X1 NOT_4349( .ZN(g13225), .A(g9873) );
  INV_X1 NOT_4350( .ZN(g13226), .A(g9876) );
  INV_X1 NOT_4351( .ZN(g13227), .A(g9880) );
  INV_X1 NOT_4352( .ZN(II20278), .A(g9027) );
  INV_X1 NOT_4353( .ZN(g13229), .A(II20278) );
  INV_X1 NOT_4354( .ZN(g13232), .A(g9895) );
  INV_X1 NOT_4355( .ZN(g13233), .A(g9898) );
  INV_X1 NOT_4356( .ZN(II20283), .A(g9050) );
  INV_X1 NOT_4357( .ZN(g13234), .A(II20283) );
  INV_X1 NOT_4358( .ZN(g13237), .A(g9913) );
  INV_X1 NOT_4359( .ZN(g13238), .A(g9916) );
  INV_X1 NOT_4360( .ZN(g13239), .A(g9933) );
  INV_X1 NOT_4361( .ZN(g13240), .A(g9936) );
  INV_X1 NOT_4362( .ZN(g13241), .A(g9958) );
  INV_X1 NOT_4363( .ZN(g13242), .A(g9962) );
  INV_X1 NOT_4364( .ZN(g13243), .A(g9965) );
  INV_X1 NOT_4365( .ZN(g13244), .A(g10004) );
  INV_X1 NOT_4366( .ZN(II20295), .A(g10015) );
  INV_X1 NOT_4367( .ZN(g13246), .A(II20295) );
  INV_X1 NOT_4368( .ZN(II20299), .A(g10800) );
  INV_X1 NOT_4369( .ZN(g13248), .A(II20299) );
  INV_X1 NOT_4370( .ZN(g13249), .A(g10018) );
  INV_X1 NOT_4371( .ZN(g13250), .A(g10021) );
  INV_X1 NOT_4372( .ZN(II20305), .A(g9050) );
  INV_X1 NOT_4373( .ZN(g13252), .A(II20305) );
  INV_X1 NOT_4374( .ZN(g13255), .A(g10049) );
  INV_X1 NOT_4375( .ZN(g13256), .A(g10052) );
  INV_X1 NOT_4376( .ZN(II20310), .A(g9067) );
  INV_X1 NOT_4377( .ZN(g13257), .A(II20310) );
  INV_X2 NOT_4378( .ZN(g13260), .A(g10067) );
  INV_X2 NOT_4379( .ZN(g13261), .A(g10070) );
  INV_X2 NOT_4380( .ZN(g13262), .A(g10087) );
  INV_X1 NOT_4381( .ZN(g13263), .A(g10090) );
  INV_X1 NOT_4382( .ZN(g13264), .A(g10096) );
  INV_X1 NOT_4383( .ZN(g13265), .A(g8568) );
  INV_X1 NOT_4384( .ZN(II20320), .A(g10792) );
  INV_X1 NOT_4385( .ZN(g13267), .A(II20320) );
  INV_X1 NOT_4386( .ZN(g13268), .A(g10109) );
  INV_X1 NOT_4387( .ZN(II20324), .A(g10124) );
  INV_X1 NOT_4388( .ZN(g13269), .A(II20324) );
  INV_X1 NOT_4389( .ZN(II20328), .A(g10817) );
  INV_X1 NOT_4390( .ZN(g13271), .A(II20328) );
  INV_X1 NOT_4391( .ZN(g13272), .A(g10127) );
  INV_X1 NOT_4392( .ZN(g13273), .A(g10130) );
  INV_X1 NOT_4393( .ZN(II20334), .A(g9067) );
  INV_X1 NOT_4394( .ZN(g13275), .A(II20334) );
  INV_X1 NOT_4395( .ZN(g13278), .A(g10158) );
  INV_X1 NOT_4396( .ZN(g13279), .A(g10161) );
  INV_X1 NOT_4397( .ZN(II20339), .A(g9084) );
  INV_X1 NOT_4398( .ZN(g13280), .A(II20339) );
  INV_X1 NOT_4399( .ZN(g13283), .A(g10176) );
  INV_X1 NOT_4400( .ZN(g13284), .A(g10179) );
  INV_X1 NOT_4401( .ZN(g13285), .A(g10189) );
  INV_X1 NOT_4402( .ZN(II20347), .A(g10787) );
  INV_X1 NOT_4403( .ZN(g13290), .A(II20347) );
  INV_X1 NOT_4404( .ZN(II20351), .A(g10804) );
  INV_X1 NOT_4405( .ZN(g13292), .A(II20351) );
  INV_X1 NOT_4406( .ZN(g13293), .A(g10214) );
  INV_X1 NOT_4407( .ZN(II20355), .A(g10229) );
  INV_X1 NOT_4408( .ZN(g13294), .A(II20355) );
  INV_X1 NOT_4409( .ZN(II20359), .A(g10838) );
  INV_X1 NOT_4410( .ZN(g13296), .A(II20359) );
  INV_X1 NOT_4411( .ZN(g13297), .A(g10232) );
  INV_X1 NOT_4412( .ZN(g13298), .A(g10235) );
  INV_X1 NOT_4413( .ZN(II20365), .A(g9084) );
  INV_X1 NOT_4414( .ZN(g13300), .A(II20365) );
  INV_X1 NOT_4415( .ZN(g13303), .A(g10263) );
  INV_X1 NOT_4416( .ZN(g13304), .A(g10266) );
  INV_X1 NOT_4417( .ZN(g13308), .A(g10273) );
  INV_X1 NOT_4418( .ZN(g13309), .A(g10276) );
  INV_X1 NOT_4419( .ZN(II20376), .A(g8569) );
  INV_X1 NOT_4420( .ZN(g13317), .A(II20376) );
  INV_X1 NOT_4421( .ZN(II20379), .A(g11213) );
  INV_X1 NOT_4422( .ZN(g13318), .A(II20379) );
  INV_X1 NOT_4423( .ZN(II20382), .A(g10907) );
  INV_X1 NOT_4424( .ZN(g13319), .A(II20382) );
  INV_X1 NOT_4425( .ZN(II20386), .A(g10796) );
  INV_X1 NOT_4426( .ZN(g13321), .A(II20386) );
  INV_X1 NOT_4427( .ZN(II20390), .A(g10821) );
  INV_X1 NOT_4428( .ZN(g13323), .A(II20390) );
  INV_X1 NOT_4429( .ZN(g13324), .A(g10316) );
  INV_X1 NOT_4430( .ZN(II20394), .A(g10331) );
  INV_X1 NOT_4431( .ZN(g13325), .A(II20394) );
  INV_X1 NOT_4432( .ZN(II20398), .A(g10858) );
  INV_X1 NOT_4433( .ZN(g13327), .A(II20398) );
  INV_X1 NOT_4434( .ZN(g13328), .A(g10334) );
  INV_X1 NOT_4435( .ZN(g13329), .A(g10337) );
  INV_X1 NOT_4436( .ZN(g13330), .A(g10357) );
  INV_X1 NOT_4437( .ZN(II20407), .A(g9027) );
  INV_X1 NOT_4438( .ZN(g13336), .A(II20407) );
  INV_X1 NOT_4439( .ZN(II20410), .A(g10887) );
  INV_X1 NOT_4440( .ZN(g13339), .A(II20410) );
  INV_X1 NOT_4441( .ZN(II20414), .A(g8575) );
  INV_X1 NOT_4442( .ZN(g13341), .A(II20414) );
  INV_X1 NOT_4443( .ZN(II20417), .A(g10933) );
  INV_X1 NOT_4444( .ZN(g13342), .A(II20417) );
  INV_X1 NOT_4445( .ZN(II20421), .A(g10808) );
  INV_X1 NOT_4446( .ZN(g13344), .A(II20421) );
  INV_X1 NOT_4447( .ZN(II20425), .A(g10842) );
  INV_X1 NOT_4448( .ZN(g13346), .A(II20425) );
  INV_X1 NOT_4449( .ZN(g13347), .A(g10409) );
  INV_X1 NOT_4450( .ZN(g13351), .A(g10416) );
  INV_X1 NOT_4451( .ZN(g13352), .A(g10419) );
  INV_X1 NOT_4452( .ZN(II20441), .A(g9027) );
  INV_X1 NOT_4453( .ZN(g13356), .A(II20441) );
  INV_X1 NOT_4454( .ZN(II20444), .A(g10869) );
  INV_X1 NOT_4455( .ZN(g13359), .A(II20444) );
  INV_X1 NOT_4456( .ZN(II20448), .A(g9050) );
  INV_X1 NOT_4457( .ZN(g13361), .A(II20448) );
  INV_X1 NOT_4458( .ZN(II20451), .A(g10908) );
  INV_X1 NOT_4459( .ZN(g13364), .A(II20451) );
  INV_X1 NOT_4460( .ZN(II20455), .A(g8578) );
  INV_X1 NOT_4461( .ZN(g13366), .A(II20455) );
  INV_X1 NOT_4462( .ZN(II20458), .A(g10972) );
  INV_X1 NOT_4463( .ZN(g13367), .A(II20458) );
  INV_X1 NOT_4464( .ZN(II20462), .A(g10825) );
  INV_X1 NOT_4465( .ZN(g13369), .A(II20462) );
  INV_X1 NOT_4466( .ZN(g13373), .A(g10482) );
  INV_X1 NOT_4467( .ZN(II20476), .A(g9027) );
  INV_X1 NOT_4468( .ZN(g13381), .A(II20476) );
  INV_X1 NOT_4469( .ZN(II20479), .A(g10849) );
  INV_X1 NOT_4470( .ZN(g13384), .A(II20479) );
  INV_X1 NOT_4471( .ZN(II20483), .A(g9050) );
  INV_X1 NOT_4472( .ZN(g13386), .A(II20483) );
  INV_X1 NOT_4473( .ZN(II20486), .A(g10889) );
  INV_X1 NOT_4474( .ZN(g13389), .A(II20486) );
  INV_X1 NOT_4475( .ZN(II20490), .A(g9067) );
  INV_X1 NOT_4476( .ZN(g13391), .A(II20490) );
  INV_X1 NOT_4477( .ZN(II20493), .A(g10934) );
  INV_X1 NOT_4478( .ZN(g13394), .A(II20493) );
  INV_X1 NOT_4479( .ZN(II20497), .A(g8579) );
  INV_X1 NOT_4480( .ZN(g13396), .A(II20497) );
  INV_X1 NOT_4481( .ZN(II20500), .A(g11007) );
  INV_X1 NOT_4482( .ZN(g13397), .A(II20500) );
  INV_X1 NOT_4483( .ZN(g13398), .A(g10542) );
  INV_X1 NOT_4484( .ZN(g13400), .A(g10545) );
  INV_X1 NOT_4485( .ZN(II20514), .A(g11769) );
  INV_X1 NOT_4486( .ZN(g13405), .A(II20514) );
  INV_X1 NOT_4487( .ZN(II20517), .A(g12425) );
  INV_X1 NOT_4488( .ZN(g13406), .A(II20517) );
  INV_X1 NOT_4489( .ZN(II20520), .A(g13246) );
  INV_X1 NOT_4490( .ZN(g13407), .A(II20520) );
  INV_X1 NOT_4491( .ZN(II20523), .A(g13317) );
  INV_X1 NOT_4492( .ZN(g13408), .A(II20523) );
  INV_X1 NOT_4493( .ZN(II20526), .A(g12519) );
  INV_X1 NOT_4494( .ZN(g13409), .A(II20526) );
  INV_X1 NOT_4495( .ZN(II20529), .A(g13319) );
  INV_X1 NOT_4496( .ZN(g13410), .A(II20529) );
  INV_X1 NOT_4497( .ZN(II20532), .A(g13339) );
  INV_X1 NOT_4498( .ZN(g13411), .A(II20532) );
  INV_X1 NOT_4499( .ZN(II20535), .A(g13359) );
  INV_X1 NOT_4500( .ZN(g13412), .A(II20535) );
  INV_X1 NOT_4501( .ZN(II20538), .A(g13384) );
  INV_X1 NOT_4502( .ZN(g13413), .A(II20538) );
  INV_X1 NOT_4503( .ZN(II20541), .A(g11599) );
  INV_X1 NOT_4504( .ZN(g13414), .A(II20541) );
  INV_X1 NOT_4505( .ZN(II20544), .A(g11628) );
  INV_X1 NOT_4506( .ZN(g13415), .A(II20544) );
  INV_X1 NOT_4507( .ZN(II20547), .A(g13248) );
  INV_X1 NOT_4508( .ZN(g13416), .A(II20547) );
  INV_X1 NOT_4509( .ZN(II20550), .A(g13267) );
  INV_X1 NOT_4510( .ZN(g13417), .A(II20550) );
  INV_X1 NOT_4511( .ZN(II20553), .A(g13290) );
  INV_X1 NOT_4512( .ZN(g13418), .A(II20553) );
  INV_X1 NOT_4513( .ZN(II20556), .A(g12435) );
  INV_X1 NOT_4514( .ZN(g13419), .A(II20556) );
  INV_X1 NOT_4515( .ZN(II20559), .A(g11937) );
  INV_X1 NOT_4516( .ZN(g13420), .A(II20559) );
  INV_X1 NOT_4517( .ZN(II20562), .A(g11786) );
  INV_X1 NOT_4518( .ZN(g13421), .A(II20562) );
  INV_X1 NOT_4519( .ZN(II20565), .A(g12432) );
  INV_X1 NOT_4520( .ZN(g13422), .A(II20565) );
  INV_X1 NOT_4521( .ZN(II20568), .A(g13269) );
  INV_X1 NOT_4522( .ZN(g13423), .A(II20568) );
  INV_X1 NOT_4523( .ZN(II20571), .A(g13341) );
  INV_X1 NOT_4524( .ZN(g13424), .A(II20571) );
  INV_X1 NOT_4525( .ZN(II20574), .A(g12534) );
  INV_X1 NOT_4526( .ZN(g13425), .A(II20574) );
  INV_X1 NOT_4527( .ZN(II20577), .A(g13342) );
  INV_X1 NOT_4528( .ZN(g13426), .A(II20577) );
  INV_X1 NOT_4529( .ZN(II20580), .A(g13364) );
  INV_X1 NOT_4530( .ZN(g13427), .A(II20580) );
  INV_X1 NOT_4531( .ZN(II20583), .A(g13389) );
  INV_X1 NOT_4532( .ZN(g13428), .A(II20583) );
  INV_X1 NOT_4533( .ZN(II20586), .A(g11606) );
  INV_X1 NOT_4534( .ZN(g13429), .A(II20586) );
  INV_X1 NOT_4535( .ZN(II20589), .A(g11629) );
  INV_X1 NOT_4536( .ZN(g13430), .A(II20589) );
  INV_X1 NOT_4537( .ZN(II20592), .A(g11651) );
  INV_X1 NOT_4538( .ZN(g13431), .A(II20592) );
  INV_X1 NOT_4539( .ZN(II20595), .A(g13271) );
  INV_X1 NOT_4540( .ZN(g13432), .A(II20595) );
  INV_X1 NOT_4541( .ZN(II20598), .A(g13292) );
  INV_X1 NOT_4542( .ZN(g13433), .A(II20598) );
  INV_X1 NOT_4543( .ZN(II20601), .A(g13321) );
  INV_X1 NOT_4544( .ZN(g13434), .A(II20601) );
  INV_X1 NOT_4545( .ZN(II20604), .A(g12440) );
  INV_X1 NOT_4546( .ZN(g13435), .A(II20604) );
  INV_X1 NOT_4547( .ZN(II20607), .A(g11990) );
  INV_X1 NOT_4548( .ZN(g13436), .A(II20607) );
  INV_X1 NOT_4549( .ZN(II20610), .A(g11812) );
  INV_X1 NOT_4550( .ZN(g13437), .A(II20610) );
  INV_X1 NOT_4551( .ZN(II20613), .A(g12437) );
  INV_X1 NOT_4552( .ZN(g13438), .A(II20613) );
  INV_X1 NOT_4553( .ZN(II20616), .A(g13294) );
  INV_X1 NOT_4554( .ZN(g13439), .A(II20616) );
  INV_X1 NOT_4555( .ZN(II20619), .A(g13366) );
  INV_X1 NOT_4556( .ZN(g13440), .A(II20619) );
  INV_X1 NOT_4557( .ZN(II20622), .A(g12543) );
  INV_X1 NOT_4558( .ZN(g13441), .A(II20622) );
  INV_X1 NOT_4559( .ZN(II20625), .A(g13367) );
  INV_X1 NOT_4560( .ZN(g13442), .A(II20625) );
  INV_X1 NOT_4561( .ZN(II20628), .A(g13394) );
  INV_X1 NOT_4562( .ZN(g13443), .A(II20628) );
  INV_X1 NOT_4563( .ZN(II20631), .A(g11611) );
  INV_X1 NOT_4564( .ZN(g13444), .A(II20631) );
  INV_X1 NOT_4565( .ZN(II20634), .A(g11636) );
  INV_X1 NOT_4566( .ZN(g13445), .A(II20634) );
  INV_X1 NOT_4567( .ZN(II20637), .A(g11652) );
  INV_X1 NOT_4568( .ZN(g13446), .A(II20637) );
  INV_X1 NOT_4569( .ZN(II20640), .A(g11670) );
  INV_X1 NOT_4570( .ZN(g13447), .A(II20640) );
  INV_X1 NOT_4571( .ZN(II20643), .A(g13296) );
  INV_X1 NOT_4572( .ZN(g13448), .A(II20643) );
  INV_X1 NOT_4573( .ZN(II20646), .A(g13323) );
  INV_X1 NOT_4574( .ZN(g13449), .A(II20646) );
  INV_X1 NOT_4575( .ZN(II20649), .A(g13344) );
  INV_X1 NOT_4576( .ZN(g13450), .A(II20649) );
  INV_X1 NOT_4577( .ZN(II20652), .A(g12445) );
  INV_X1 NOT_4578( .ZN(g13451), .A(II20652) );
  INV_X1 NOT_4579( .ZN(II20655), .A(g12059) );
  INV_X1 NOT_4580( .ZN(g13452), .A(II20655) );
  INV_X1 NOT_4581( .ZN(II20658), .A(g11845) );
  INV_X1 NOT_4582( .ZN(g13453), .A(II20658) );
  INV_X1 NOT_4583( .ZN(II20661), .A(g12442) );
  INV_X1 NOT_4584( .ZN(g13454), .A(II20661) );
  INV_X1 NOT_4585( .ZN(II20664), .A(g13325) );
  INV_X1 NOT_4586( .ZN(g13455), .A(II20664) );
  INV_X1 NOT_4587( .ZN(II20667), .A(g13396) );
  INV_X1 NOT_4588( .ZN(g13456), .A(II20667) );
  INV_X1 NOT_4589( .ZN(II20670), .A(g12552) );
  INV_X1 NOT_4590( .ZN(g13457), .A(II20670) );
  INV_X1 NOT_4591( .ZN(II20673), .A(g13397) );
  INV_X1 NOT_4592( .ZN(g13458), .A(II20673) );
  INV_X1 NOT_4593( .ZN(II20676), .A(g11616) );
  INV_X1 NOT_4594( .ZN(g13459), .A(II20676) );
  INV_X1 NOT_4595( .ZN(II20679), .A(g11641) );
  INV_X1 NOT_4596( .ZN(g13460), .A(II20679) );
  INV_X1 NOT_4597( .ZN(II20682), .A(g11659) );
  INV_X1 NOT_4598( .ZN(g13461), .A(II20682) );
  INV_X1 NOT_4599( .ZN(II20685), .A(g11671) );
  INV_X1 NOT_4600( .ZN(g13462), .A(II20685) );
  INV_X1 NOT_4601( .ZN(II20688), .A(g11682) );
  INV_X1 NOT_4602( .ZN(g13463), .A(II20688) );
  INV_X1 NOT_4603( .ZN(II20691), .A(g13327) );
  INV_X1 NOT_4604( .ZN(g13464), .A(II20691) );
  INV_X1 NOT_4605( .ZN(II20694), .A(g13346) );
  INV_X1 NOT_4606( .ZN(g13465), .A(II20694) );
  INV_X1 NOT_4607( .ZN(II20697), .A(g13369) );
  INV_X1 NOT_4608( .ZN(g13466), .A(II20697) );
  INV_X1 NOT_4609( .ZN(II20700), .A(g12450) );
  INV_X1 NOT_4610( .ZN(g13467), .A(II20700) );
  INV_X1 NOT_4611( .ZN(II20703), .A(g12123) );
  INV_X1 NOT_4612( .ZN(g13468), .A(II20703) );
  INV_X1 NOT_4613( .ZN(II20706), .A(g11490) );
  INV_X2 NOT_4614( .ZN(g13469), .A(II20706) );
  INV_X2 NOT_4615( .ZN(II20709), .A(g13070) );
  INV_X1 NOT_4616( .ZN(g13475), .A(II20709) );
  INV_X1 NOT_4617( .ZN(g13519), .A(g13228) );
  INV_X1 NOT_4618( .ZN(g13530), .A(g13251) );
  INV_X1 NOT_4619( .ZN(g13541), .A(g13274) );
  INV_X1 NOT_4620( .ZN(g13552), .A(g13299) );
  INV_X1 NOT_4621( .ZN(g13565), .A(g12192) );
  INV_X1 NOT_4622( .ZN(g13568), .A(g11627) );
  INV_X1 NOT_4623( .ZN(II20791), .A(g13149) );
  INV_X1 NOT_4624( .ZN(g13571), .A(II20791) );
  INV_X1 NOT_4625( .ZN(II20794), .A(g13111) );
  INV_X1 NOT_4626( .ZN(g13572), .A(II20794) );
  INV_X1 NOT_4627( .ZN(g13573), .A(g12247) );
  INV_X1 NOT_4628( .ZN(g13576), .A(g11650) );
  INV_X1 NOT_4629( .ZN(II20799), .A(g13155) );
  INV_X1 NOT_4630( .ZN(g13579), .A(II20799) );
  INV_X1 NOT_4631( .ZN(II20802), .A(g13160) );
  INV_X1 NOT_4632( .ZN(g13580), .A(II20802) );
  INV_X1 NOT_4633( .ZN(II20805), .A(g13124) );
  INV_X1 NOT_4634( .ZN(g13581), .A(II20805) );
  INV_X1 NOT_4635( .ZN(g13582), .A(g12290) );
  INV_X1 NOT_4636( .ZN(g13585), .A(g11669) );
  INV_X1 NOT_4637( .ZN(II20810), .A(g13164) );
  INV_X1 NOT_4638( .ZN(g13588), .A(II20810) );
  INV_X1 NOT_4639( .ZN(II20813), .A(g13265) );
  INV_X1 NOT_4640( .ZN(g13589), .A(II20813) );
  INV_X1 NOT_4641( .ZN(II20816), .A(g12487) );
  INV_X1 NOT_4642( .ZN(g13598), .A(II20816) );
  INV_X1 NOT_4643( .ZN(II20820), .A(g13171) );
  INV_X1 NOT_4644( .ZN(g13600), .A(II20820) );
  INV_X1 NOT_4645( .ZN(II20823), .A(g13135) );
  INV_X1 NOT_4646( .ZN(g13601), .A(II20823) );
  INV_X1 NOT_4647( .ZN(g13602), .A(g12326) );
  INV_X1 NOT_4648( .ZN(g13605), .A(g11681) );
  INV_X1 NOT_4649( .ZN(II20828), .A(g13175) );
  INV_X1 NOT_4650( .ZN(g13608), .A(II20828) );
  INV_X1 NOT_4651( .ZN(II20832), .A(g12507) );
  INV_X1 NOT_4652( .ZN(g13610), .A(II20832) );
  INV_X1 NOT_4653( .ZN(II20836), .A(g13182) );
  INV_X1 NOT_4654( .ZN(g13612), .A(II20836) );
  INV_X1 NOT_4655( .ZN(II20839), .A(g13143) );
  INV_X1 NOT_4656( .ZN(g13613), .A(II20839) );
  INV_X1 NOT_4657( .ZN(g13614), .A(g11690) );
  INV_X1 NOT_4658( .ZN(II20844), .A(g12524) );
  INV_X1 NOT_4659( .ZN(g13620), .A(II20844) );
  INV_X1 NOT_4660( .ZN(II20848), .A(g13194) );
  INV_X1 NOT_4661( .ZN(g13622), .A(II20848) );
  INV_X1 NOT_4662( .ZN(II20852), .A(g12457) );
  INV_X1 NOT_4663( .ZN(g13624), .A(II20852) );
  INV_X1 NOT_4664( .ZN(g13626), .A(g11697) );
  INV_X1 NOT_4665( .ZN(II20858), .A(g12539) );
  INV_X1 NOT_4666( .ZN(g13632), .A(II20858) );
  INV_X1 NOT_4667( .ZN(II20863), .A(g12467) );
  INV_X1 NOT_4668( .ZN(g13635), .A(II20863) );
  INV_X1 NOT_4669( .ZN(g13637), .A(g11703) );
  INV_X1 NOT_4670( .ZN(g13644), .A(g13215) );
  INV_X1 NOT_4671( .ZN(II20873), .A(g12482) );
  INV_X1 NOT_4672( .ZN(g13647), .A(II20873) );
  INV_X1 NOT_4673( .ZN(g13649), .A(g11711) );
  INV_X1 NOT_4674( .ZN(g13657), .A(g12452) );
  INV_X1 NOT_4675( .ZN(g13669), .A(g13229) );
  INV_X1 NOT_4676( .ZN(g13670), .A(g13234) );
  INV_X1 NOT_4677( .ZN(II20886), .A(g12499) );
  INV_X1 NOT_4678( .ZN(g13673), .A(II20886) );
  INV_X1 NOT_4679( .ZN(g13677), .A(g12447) );
  INV_X1 NOT_4680( .ZN(g13687), .A(g12460) );
  INV_X1 NOT_4681( .ZN(g13699), .A(g13252) );
  INV_X1 NOT_4682( .ZN(g13700), .A(g13257) );
  INV_X1 NOT_4683( .ZN(g13706), .A(g12443) );
  INV_X1 NOT_4684( .ZN(g13714), .A(g12453) );
  INV_X1 NOT_4685( .ZN(g13724), .A(g12470) );
  INV_X1 NOT_4686( .ZN(g13736), .A(g13275) );
  INV_X1 NOT_4687( .ZN(g13737), .A(g13280) );
  INV_X1 NOT_4688( .ZN(II20909), .A(g13055) );
  INV_X1 NOT_4689( .ZN(g13741), .A(II20909) );
  INV_X1 NOT_4690( .ZN(g13750), .A(g12439) );
  INV_X1 NOT_4691( .ZN(g13756), .A(g12448) );
  INV_X1 NOT_4692( .ZN(g13764), .A(g12461) );
  INV_X1 NOT_4693( .ZN(g13774), .A(g12485) );
  INV_X1 NOT_4694( .ZN(g13786), .A(g13300) );
  INV_X1 NOT_4695( .ZN(g13791), .A(g12444) );
  INV_X1 NOT_4696( .ZN(g13797), .A(g12454) );
  INV_X1 NOT_4697( .ZN(g13805), .A(g12471) );
  INV_X1 NOT_4698( .ZN(g13817), .A(g13336) );
  INV_X1 NOT_4699( .ZN(g13819), .A(g12449) );
  INV_X1 NOT_4700( .ZN(g13825), .A(g12462) );
  INV_X1 NOT_4701( .ZN(g13836), .A(g13356) );
  INV_X1 NOT_4702( .ZN(g13838), .A(g13361) );
  INV_X1 NOT_4703( .ZN(g13840), .A(g12455) );
  INV_X1 NOT_4704( .ZN(g13848), .A(g11744) );
  INV_X1 NOT_4705( .ZN(g13849), .A(g13381) );
  INV_X1 NOT_4706( .ZN(g13850), .A(g13386) );
  INV_X1 NOT_4707( .ZN(g13852), .A(g13391) );
  INV_X1 NOT_4708( .ZN(g13856), .A(g11759) );
  INV_X1 NOT_4709( .ZN(g13857), .A(g11760) );
  INV_X1 NOT_4710( .ZN(g13858), .A(g11603) );
  INV_X1 NOT_4711( .ZN(g13859), .A(g11608) );
  INV_X1 NOT_4712( .ZN(g13861), .A(g11613) );
  INV_X1 NOT_4713( .ZN(II20959), .A(g11713) );
  INV_X1 NOT_4714( .ZN(g13863), .A(II20959) );
  INV_X1 NOT_4715( .ZN(g13864), .A(g11767) );
  INV_X1 NOT_4716( .ZN(g13866), .A(g11772) );
  INV_X1 NOT_4717( .ZN(g13867), .A(g11773) );
  INV_X1 NOT_4718( .ZN(g13868), .A(g11633) );
  INV_X1 NOT_4719( .ZN(g13869), .A(g11638) );
  INV_X1 NOT_4720( .ZN(g13872), .A(g11780) );
  INV_X1 NOT_4721( .ZN(g13873), .A(g12698) );
  INV_X1 NOT_4722( .ZN(g13879), .A(g11784) );
  INV_X1 NOT_4723( .ZN(g13881), .A(g11789) );
  INV_X1 NOT_4724( .ZN(g13882), .A(g11790) );
  INV_X1 NOT_4725( .ZN(g13883), .A(g11656) );
  INV_X1 NOT_4726( .ZN(g13885), .A(g11799) );
  INV_X1 NOT_4727( .ZN(g13886), .A(g12747) );
  INV_X1 NOT_4728( .ZN(g13894), .A(g11806) );
  INV_X1 NOT_4729( .ZN(g13895), .A(g12755) );
  INV_X1 NOT_4730( .ZN(g13901), .A(g11810) );
  INV_X1 NOT_4731( .ZN(g13903), .A(g11815) );
  INV_X1 NOT_4732( .ZN(g13906), .A(g11822) );
  INV_X1 NOT_4733( .ZN(g13907), .A(g12781) );
  INV_X1 NOT_4734( .ZN(g13918), .A(g11830) );
  INV_X1 NOT_4735( .ZN(g13922), .A(g11831) );
  INV_X1 NOT_4736( .ZN(g13926), .A(g11832) );
  INV_X1 NOT_4737( .ZN(g13927), .A(g12789) );
  INV_X1 NOT_4738( .ZN(g13935), .A(g11839) );
  INV_X1 NOT_4739( .ZN(g13936), .A(g12797) );
  INV_X1 NOT_4740( .ZN(g13942), .A(g11843) );
  INV_X1 NOT_4741( .ZN(g13945), .A(g11855) );
  INV_X1 NOT_4742( .ZN(g13946), .A(g12814) );
  INV_X1 NOT_4743( .ZN(II21012), .A(g12503) );
  INV_X1 NOT_4744( .ZN(g13954), .A(II21012) );
  INV_X1 NOT_4745( .ZN(g13958), .A(g11863) );
  INV_X1 NOT_4746( .ZN(g13962), .A(g11864) );
  INV_X1 NOT_4747( .ZN(g13963), .A(g12820) );
  INV_X1 NOT_4748( .ZN(g13974), .A(g11872) );
  INV_X1 NOT_4749( .ZN(g13978), .A(g11873) );
  INV_X1 NOT_4750( .ZN(g13982), .A(g11874) );
  INV_X1 NOT_4751( .ZN(g13983), .A(g12828) );
  INV_X1 NOT_4752( .ZN(g13991), .A(g11881) );
  INV_X1 NOT_4753( .ZN(g13992), .A(g12836) );
  INV_X1 NOT_4754( .ZN(g13999), .A(g11889) );
  INV_X1 NOT_4755( .ZN(g14000), .A(g11890) );
  INV_X1 NOT_4756( .ZN(g14001), .A(g12849) );
  INV_X1 NOT_4757( .ZN(II21037), .A(g12486) );
  INV_X1 NOT_4758( .ZN(g14008), .A(II21037) );
  INV_X1 NOT_4759( .ZN(g14011), .A(g11896) );
  INV_X1 NOT_4760( .ZN(g14015), .A(g11897) );
  INV_X1 NOT_4761( .ZN(g14016), .A(g12852) );
  INV_X1 NOT_4762( .ZN(II21045), .A(g12520) );
  INV_X1 NOT_4763( .ZN(g14024), .A(II21045) );
  INV_X1 NOT_4764( .ZN(g14028), .A(g11905) );
  INV_X1 NOT_4765( .ZN(g14032), .A(g11906) );
  INV_X1 NOT_4766( .ZN(g14033), .A(g12858) );
  INV_X1 NOT_4767( .ZN(g14044), .A(g11914) );
  INV_X1 NOT_4768( .ZN(g14048), .A(g11915) );
  INV_X1 NOT_4769( .ZN(g14052), .A(g11916) );
  INV_X1 NOT_4770( .ZN(g14053), .A(g12866) );
  INV_X1 NOT_4771( .ZN(g14061), .A(g11928) );
  INV_X1 NOT_4772( .ZN(g14062), .A(g12880) );
  INV_X1 NOT_4773( .ZN(II21064), .A(g13147) );
  INV_X1 NOT_4774( .ZN(g14068), .A(II21064) );
  INV_X1 NOT_4775( .ZN(g14071), .A(g11934) );
  INV_X1 NOT_4776( .ZN(g14079), .A(g11935) );
  INV_X1 NOT_4777( .ZN(g14086), .A(g11938) );
  INV_X1 NOT_4778( .ZN(g14090), .A(g11939) );
  INV_X1 NOT_4779( .ZN(g14091), .A(g11940) );
  INV_X1 NOT_4780( .ZN(g14092), .A(g12890) );
  INV_X1 NOT_4781( .ZN(II21075), .A(g12506) );
  INV_X1 NOT_4782( .ZN(g14099), .A(II21075) );
  INV_X1 NOT_4783( .ZN(g14102), .A(g11946) );
  INV_X1 NOT_4784( .ZN(g14106), .A(g11947) );
  INV_X1 NOT_4785( .ZN(g14107), .A(g12893) );
  INV_X1 NOT_4786( .ZN(II21083), .A(g12535) );
  INV_X1 NOT_4787( .ZN(g14115), .A(II21083) );
  INV_X1 NOT_4788( .ZN(g14119), .A(g11955) );
  INV_X1 NOT_4789( .ZN(g14123), .A(g11956) );
  INV_X1 NOT_4790( .ZN(g14124), .A(g12899) );
  INV_X1 NOT_4791( .ZN(g14135), .A(g11964) );
  INV_X1 NOT_4792( .ZN(g14139), .A(g11965) );
  INV_X1 NOT_4793( .ZN(II21096), .A(g11749) );
  INV_X1 NOT_4794( .ZN(g14144), .A(II21096) );
  INV_X1 NOT_4795( .ZN(g14148), .A(g12912) );
  INV_X1 NOT_4796( .ZN(g14153), .A(g12913) );
  INV_X1 NOT_4797( .ZN(g14158), .A(g11974) );
  INV_X1 NOT_4798( .ZN(g14165), .A(g11975) );
  INV_X1 NOT_4799( .ZN(g14171), .A(g11979) );
  INV_X1 NOT_4800( .ZN(g14175), .A(g11980) );
  INV_X1 NOT_4801( .ZN(g14176), .A(g11981) );
  INV_X1 NOT_4802( .ZN(g14177), .A(g12920) );
  INV_X1 NOT_4803( .ZN(II21108), .A(g13150) );
  INV_X1 NOT_4804( .ZN(g14183), .A(II21108) );
  INV_X1 NOT_4805( .ZN(g14186), .A(g11987) );
  INV_X1 NOT_4806( .ZN(g14194), .A(g11988) );
  INV_X1 NOT_4807( .ZN(g14201), .A(g11991) );
  INV_X1 NOT_4808( .ZN(g14205), .A(g11992) );
  INV_X1 NOT_4809( .ZN(g14206), .A(g11993) );
  INV_X1 NOT_4810( .ZN(g14207), .A(g12930) );
  INV_X1 NOT_4811( .ZN(II21119), .A(g12523) );
  INV_X1 NOT_4812( .ZN(g14214), .A(II21119) );
  INV_X1 NOT_4813( .ZN(g14217), .A(g11999) );
  INV_X1 NOT_4814( .ZN(g14221), .A(g12000) );
  INV_X1 NOT_4815( .ZN(g14222), .A(g12933) );
  INV_X1 NOT_4816( .ZN(II21127), .A(g12544) );
  INV_X1 NOT_4817( .ZN(g14230), .A(II21127) );
  INV_X1 NOT_4818( .ZN(g14234), .A(g12008) );
  INV_X1 NOT_4819( .ZN(g14238), .A(g12939) );
  INV_X1 NOT_4820( .ZN(g14244), .A(g12026) );
  INV_X1 NOT_4821( .ZN(g14249), .A(g12034) );
  INV_X1 NOT_4822( .ZN(g14252), .A(g12035) );
  INV_X1 NOT_4823( .ZN(g14256), .A(g12036) );
  INV_X1 NOT_4824( .ZN(II21137), .A(g11749) );
  INV_X1 NOT_4825( .ZN(g14259), .A(II21137) );
  INV_X1 NOT_4826( .ZN(g14263), .A(g12941) );
  INV_X1 NOT_4827( .ZN(g14268), .A(g12942) );
  INV_X1 NOT_4828( .ZN(g14273), .A(g12043) );
  INV_X1 NOT_4829( .ZN(g14280), .A(g12044) );
  INV_X1 NOT_4830( .ZN(g14286), .A(g12048) );
  INV_X1 NOT_4831( .ZN(g14290), .A(g12049) );
  INV_X1 NOT_4832( .ZN(g14291), .A(g12050) );
  INV_X1 NOT_4833( .ZN(g14292), .A(g12949) );
  INV_X1 NOT_4834( .ZN(II21149), .A(g13156) );
  INV_X1 NOT_4835( .ZN(g14298), .A(II21149) );
  INV_X1 NOT_4836( .ZN(g14301), .A(g12056) );
  INV_X1 NOT_4837( .ZN(g14309), .A(g12057) );
  INV_X1 NOT_4838( .ZN(g14316), .A(g12060) );
  INV_X1 NOT_4839( .ZN(g14320), .A(g12061) );
  INV_X1 NOT_4840( .ZN(g14321), .A(g12062) );
  INV_X1 NOT_4841( .ZN(g14322), .A(g12959) );
  INV_X1 NOT_4842( .ZN(II21160), .A(g12538) );
  INV_X1 NOT_4843( .ZN(g14329), .A(II21160) );
  INV_X1 NOT_4844( .ZN(g14332), .A(g12068) );
  INV_X1 NOT_4845( .ZN(II21165), .A(g13110) );
  INV_X1 NOT_4846( .ZN(g14337), .A(II21165) );
  INV_X1 NOT_4847( .ZN(g14342), .A(g12967) );
  INV_X1 NOT_4848( .ZN(g14347), .A(g12079) );
  INV_X1 NOT_4849( .ZN(g14352), .A(g12081) );
  INV_X1 NOT_4850( .ZN(g14355), .A(g12082) );
  INV_X1 NOT_4851( .ZN(g14359), .A(g12083) );
  INV_X1 NOT_4852( .ZN(g14360), .A(g12968) );
  INV_X1 NOT_4853( .ZN(g14366), .A(g12090) );
  INV_X1 NOT_4854( .ZN(g14371), .A(g12098) );
  INV_X1 NOT_4855( .ZN(g14374), .A(g12099) );
  INV_X1 NOT_4856( .ZN(g14378), .A(g12100) );
  INV_X1 NOT_4857( .ZN(II21178), .A(g11749) );
  INV_X1 NOT_4858( .ZN(g14381), .A(II21178) );
  INV_X1 NOT_4859( .ZN(g14385), .A(g12970) );
  INV_X1 NOT_4860( .ZN(g14390), .A(g12971) );
  INV_X1 NOT_4861( .ZN(g14395), .A(g12107) );
  INV_X1 NOT_4862( .ZN(g14402), .A(g12108) );
  INV_X1 NOT_4863( .ZN(g14408), .A(g12112) );
  INV_X1 NOT_4864( .ZN(g14412), .A(g12113) );
  INV_X1 NOT_4865( .ZN(g14413), .A(g12114) );
  INV_X1 NOT_4866( .ZN(g14414), .A(g12978) );
  INV_X1 NOT_4867( .ZN(II21190), .A(g13165) );
  INV_X1 NOT_4868( .ZN(g14420), .A(II21190) );
  INV_X1 NOT_4869( .ZN(g14423), .A(g12120) );
  INV_X1 NOT_4870( .ZN(g14431), .A(g12121) );
  INV_X1 NOT_4871( .ZN(g14438), .A(g12124) );
  INV_X1 NOT_4872( .ZN(g14442), .A(g11768) );
  INV_X1 NOT_4873( .ZN(g14450), .A(g12146) );
  INV_X1 NOT_4874( .ZN(g14454), .A(g12991) );
  INV_X1 NOT_4875( .ZN(g14459), .A(g12151) );
  INV_X1 NOT_4876( .ZN(g14464), .A(g12153) );
  INV_X1 NOT_4877( .ZN(g14467), .A(g12154) );
  INV_X1 NOT_4878( .ZN(g14471), .A(g12155) );
  INV_X1 NOT_4879( .ZN(g14472), .A(g12992) );
  INV_X1 NOT_4880( .ZN(g14478), .A(g12162) );
  INV_X1 NOT_4881( .ZN(g14483), .A(g12170) );
  INV_X1 NOT_4882( .ZN(g14486), .A(g12171) );
  INV_X1 NOT_4883( .ZN(g14490), .A(g12172) );
  INV_X1 NOT_4884( .ZN(II21208), .A(g11749) );
  INV_X1 NOT_4885( .ZN(g14493), .A(II21208) );
  INV_X1 NOT_4886( .ZN(g14497), .A(g12994) );
  INV_X1 NOT_4887( .ZN(g14502), .A(g12995) );
  INV_X1 NOT_4888( .ZN(g14507), .A(g12179) );
  INV_X1 NOT_4889( .ZN(g14514), .A(g12180) );
  INV_X1 NOT_4890( .ZN(g14520), .A(g12184) );
  INV_X1 NOT_4891( .ZN(g14524), .A(g12185) );
  INV_X1 NOT_4892( .ZN(g14525), .A(g12195) );
  INV_X1 NOT_4893( .ZN(g14529), .A(g11785) );
  INV_X1 NOT_4894( .ZN(g14537), .A(g12208) );
  INV_X1 NOT_4895( .ZN(g14541), .A(g13001) );
  INV_X1 NOT_4896( .ZN(g14546), .A(g12213) );
  INV_X1 NOT_4897( .ZN(g14551), .A(g12215) );
  INV_X1 NOT_4898( .ZN(g14554), .A(g12216) );
  INV_X1 NOT_4899( .ZN(g14558), .A(g12217) );
  INV_X1 NOT_4900( .ZN(g14559), .A(g13002) );
  INV_X1 NOT_4901( .ZN(g14565), .A(g12224) );
  INV_X1 NOT_4902( .ZN(g14570), .A(g12232) );
  INV_X1 NOT_4903( .ZN(g14573), .A(g12233) );
  INV_X1 NOT_4904( .ZN(g14577), .A(g12234) );
  INV_X1 NOT_4905( .ZN(g14580), .A(g12250) );
  INV_X1 NOT_4906( .ZN(g14584), .A(g11811) );
  INV_X1 NOT_4907( .ZN(g14592), .A(g12263) );
  INV_X1 NOT_4908( .ZN(g14596), .A(g13022) );
  INV_X1 NOT_4909( .ZN(g14601), .A(g12268) );
  INV_X1 NOT_4910( .ZN(g14606), .A(g12270) );
  INV_X1 NOT_4911( .ZN(g14609), .A(g12271) );
  INV_X1 NOT_4912( .ZN(g14613), .A(g12272) );
  INV_X1 NOT_4913( .ZN(g14614), .A(g12293) );
  INV_X1 NOT_4914( .ZN(g14618), .A(g11844) );
  INV_X1 NOT_4915( .ZN(g14626), .A(g12306) );
  INV_X1 NOT_4916( .ZN(II21241), .A(g13378) );
  INV_X1 NOT_4917( .ZN(g14630), .A(II21241) );
  INV_X1 NOT_4918( .ZN(g14637), .A(g12329) );
  INV_X1 NOT_4919( .ZN(g14641), .A(g11823) );
  INV_X1 NOT_4920( .ZN(II21246), .A(g11624) );
  INV_X1 NOT_4921( .ZN(g14642), .A(II21246) );
  INV_X1 NOT_4922( .ZN(II21249), .A(g11600) );
  INV_X1 NOT_4923( .ZN(g14650), .A(II21249) );
  INV_X1 NOT_4924( .ZN(II21252), .A(g11644) );
  INV_X1 NOT_4925( .ZN(g14657), .A(II21252) );
  INV_X1 NOT_4926( .ZN(g14668), .A(g11865) );
  INV_X1 NOT_4927( .ZN(II21256), .A(g11647) );
  INV_X1 NOT_4928( .ZN(g14669), .A(II21256) );
  INV_X1 NOT_4929( .ZN(II21259), .A(g11630) );
  INV_X1 NOT_4930( .ZN(g14677), .A(II21259) );
  INV_X1 NOT_4931( .ZN(II21262), .A(g11713) );
  INV_X1 NOT_4932( .ZN(g14684), .A(II21262) );
  INV_X1 NOT_4933( .ZN(g14685), .A(g12245) );
  INV_X1 NOT_4934( .ZN(II21267), .A(g11663) );
  INV_X1 NOT_4935( .ZN(g14691), .A(II21267) );
  INV_X1 NOT_4936( .ZN(g14702), .A(g11907) );
  INV_X1 NOT_4937( .ZN(II21271), .A(g11666) );
  INV_X1 NOT_4938( .ZN(g14703), .A(II21271) );
  INV_X1 NOT_4939( .ZN(II21274), .A(g11653) );
  INV_X1 NOT_4940( .ZN(g14711), .A(II21274) );
  INV_X1 NOT_4941( .ZN(II21277), .A(g12430) );
  INV_X1 NOT_4942( .ZN(g14718), .A(II21277) );
  INV_X1 NOT_4943( .ZN(g14719), .A(g12288) );
  INV_X4 NOT_4944( .ZN(II21282), .A(g11675) );
  INV_X4 NOT_4945( .ZN(g14725), .A(II21282) );
  INV_X4 NOT_4946( .ZN(g14736), .A(g11957) );
  INV_X4 NOT_4947( .ZN(II21286), .A(g11678) );
  INV_X1 NOT_4948( .ZN(g14737), .A(II21286) );
  INV_X1 NOT_4949( .ZN(II21289), .A(g12434) );
  INV_X1 NOT_4950( .ZN(g14745), .A(II21289) );
  INV_X1 NOT_4951( .ZN(II21292), .A(g11888) );
  INV_X1 NOT_4952( .ZN(g14746), .A(II21292) );
  INV_X1 NOT_4953( .ZN(g14747), .A(g12324) );
  INV_X1 NOT_4954( .ZN(II21297), .A(g11687) );
  INV_X1 NOT_4955( .ZN(g14753), .A(II21297) );
  INV_X1 NOT_4956( .ZN(g14764), .A(g11791) );
  INV_X1 NOT_4957( .ZN(II21301), .A(g12438) );
  INV_X1 NOT_4958( .ZN(g14765), .A(II21301) );
  INV_X1 NOT_4959( .ZN(II21304), .A(g11927) );
  INV_X1 NOT_4960( .ZN(g14766), .A(II21304) );
  INV_X1 NOT_4961( .ZN(g14768), .A(g12352) );
  INV_X1 NOT_4962( .ZN(II21310), .A(g12332) );
  INV_X1 NOT_4963( .ZN(g14774), .A(II21310) );
  INV_X1 NOT_4964( .ZN(II21313), .A(g11743) );
  INV_X1 NOT_4965( .ZN(g14775), .A(II21313) );
  INV_X1 NOT_4966( .ZN(g14776), .A(g12033) );
  INV_X1 NOT_4967( .ZN(g14794), .A(g11848) );
  INV_X1 NOT_4968( .ZN(II21318), .A(g12362) );
  INV_X1 NOT_4969( .ZN(g14795), .A(II21318) );
  INV_X1 NOT_4970( .ZN(II21321), .A(g11758) );
  INV_X1 NOT_4971( .ZN(g14796), .A(II21321) );
  INV_X1 NOT_4972( .ZN(g14797), .A(g12080) );
  INV_X1 NOT_4973( .ZN(g14811), .A(g12097) );
  INV_X1 NOT_4974( .ZN(II21326), .A(g12378) );
  INV_X1 NOT_4975( .ZN(g14829), .A(II21326) );
  INV_X1 NOT_4976( .ZN(II21329), .A(g11766) );
  INV_X1 NOT_4977( .ZN(g14830), .A(II21329) );
  INV_X1 NOT_4978( .ZN(g14831), .A(g11828) );
  INV_X1 NOT_4979( .ZN(g14837), .A(g12145) );
  INV_X1 NOT_4980( .ZN(g14849), .A(g12152) );
  INV_X1 NOT_4981( .ZN(g14863), .A(g12169) );
  INV_X1 NOT_4982( .ZN(g14881), .A(g11923) );
  INV_X1 NOT_4983( .ZN(II21337), .A(g12408) );
  INV_X1 NOT_4984( .ZN(g14882), .A(II21337) );
  INV_X1 NOT_4985( .ZN(II21340), .A(g11779) );
  INV_X1 NOT_4986( .ZN(g14883), .A(II21340) );
  INV_X1 NOT_4987( .ZN(g14885), .A(g11860) );
  INV_X1 NOT_4988( .ZN(g14895), .A(g12193) );
  INV_X1 NOT_4989( .ZN(g14904), .A(g11870) );
  INV_X1 NOT_4990( .ZN(g14910), .A(g12207) );
  INV_X1 NOT_4991( .ZN(g14922), .A(g12214) );
  INV_X1 NOT_4992( .ZN(g14936), .A(g12231) );
  INV_X1 NOT_4993( .ZN(II21351), .A(g12420) );
  INV_X1 NOT_4994( .ZN(g14954), .A(II21351) );
  INV_X1 NOT_4995( .ZN(II21354), .A(g11798) );
  INV_X1 NOT_4996( .ZN(g14955), .A(II21354) );
  INV_X1 NOT_4997( .ZN(g14959), .A(g11976) );
  INV_X1 NOT_4998( .ZN(II21361), .A(g13026) );
  INV_X1 NOT_4999( .ZN(g14960), .A(II21361) );
  INV_X1 NOT_5000( .ZN(II21364), .A(g13028) );
  INV_X1 NOT_5001( .ZN(g14963), .A(II21364) );
  INV_X1 NOT_5002( .ZN(g14966), .A(g11902) );
  INV_X1 NOT_5003( .ZN(g14976), .A(g12248) );
  INV_X1 NOT_5004( .ZN(g14985), .A(g11912) );
  INV_X1 NOT_5005( .ZN(g14991), .A(g12262) );
  INV_X1 NOT_5006( .ZN(g15003), .A(g12269) );
  INV_X1 NOT_5007( .ZN(g15017), .A(g12009) );
  INV_X1 NOT_5008( .ZN(II21374), .A(g12424) );
  INV_X1 NOT_5009( .ZN(g15018), .A(II21374) );
  INV_X1 NOT_5010( .ZN(II21377), .A(g11821) );
  INV_X1 NOT_5011( .ZN(g15019), .A(II21377) );
  INV_X1 NOT_5012( .ZN(II21381), .A(g13157) );
  INV_X1 NOT_5013( .ZN(g15021), .A(II21381) );
  INV_X1 NOT_5014( .ZN(g15022), .A(g11781) );
  INV_X1 NOT_5015( .ZN(g15032), .A(g12027) );
  INV_X1 NOT_5016( .ZN(g15033), .A(g12030) );
  INV_X1 NOT_5017( .ZN(II21389), .A(g12883) );
  INV_X1 NOT_5018( .ZN(g15034), .A(II21389) );
  INV_X1 NOT_5019( .ZN(II21392), .A(g13020) );
  INV_X1 NOT_5020( .ZN(g15037), .A(II21392) );
  INV_X1 NOT_5021( .ZN(II21395), .A(g13034) );
  INV_X1 NOT_5022( .ZN(g15040), .A(II21395) );
  INV_X1 NOT_5023( .ZN(II21398), .A(g13021) );
  INV_X1 NOT_5024( .ZN(g15043), .A(II21398) );
  INV_X1 NOT_5025( .ZN(g15048), .A(g12045) );
  INV_X1 NOT_5026( .ZN(II21404), .A(g13037) );
  INV_X1 NOT_5027( .ZN(g15049), .A(II21404) );
  INV_X1 NOT_5028( .ZN(II21407), .A(g13039) );
  INV_X1 NOT_5029( .ZN(g15052), .A(II21407) );
  INV_X1 NOT_5030( .ZN(g15055), .A(g11952) );
  INV_X1 NOT_5031( .ZN(g15065), .A(g12291) );
  INV_X1 NOT_5032( .ZN(g15074), .A(g11962) );
  INV_X1 NOT_5033( .ZN(g15080), .A(g12305) );
  INV_X1 NOT_5034( .ZN(II21415), .A(g11854) );
  INV_X1 NOT_5035( .ZN(g15092), .A(II21415) );
  INV_X1 NOT_5036( .ZN(II21420), .A(g13166) );
  INV_X1 NOT_5037( .ZN(g15095), .A(II21420) );
  INV_X1 NOT_5038( .ZN(g15096), .A(g11800) );
  INV_X1 NOT_5039( .ZN(II21426), .A(g11661) );
  INV_X1 NOT_5040( .ZN(g15106), .A(II21426) );
  INV_X1 NOT_5041( .ZN(II21429), .A(g13027) );
  INV_X1 NOT_5042( .ZN(g15109), .A(II21429) );
  INV_X1 NOT_5043( .ZN(II21432), .A(g13044) );
  INV_X1 NOT_5044( .ZN(g15112), .A(II21432) );
  INV_X1 NOT_5045( .ZN(II21435), .A(g11662) );
  INV_X1 NOT_5046( .ZN(g15115), .A(II21435) );
  INV_X1 NOT_5047( .ZN(g15118), .A(g11807) );
  INV_X1 NOT_5048( .ZN(g15128), .A(g12091) );
  INV_X1 NOT_5049( .ZN(g15129), .A(g12094) );
  INV_X1 NOT_5050( .ZN(II21443), .A(g12923) );
  INV_X1 NOT_5051( .ZN(g15130), .A(II21443) );
  INV_X1 NOT_5052( .ZN(II21446), .A(g13029) );
  INV_X1 NOT_5053( .ZN(g15133), .A(II21446) );
  INV_X1 NOT_5054( .ZN(II21449), .A(g13047) );
  INV_X1 NOT_5055( .ZN(g15136), .A(II21449) );
  INV_X1 NOT_5056( .ZN(II21452), .A(g13030) );
  INV_X1 NOT_5057( .ZN(g15139), .A(II21452) );
  INV_X1 NOT_5058( .ZN(g15144), .A(g12109) );
  INV_X1 NOT_5059( .ZN(II21458), .A(g13050) );
  INV_X1 NOT_5060( .ZN(g15145), .A(II21458) );
  INV_X1 NOT_5061( .ZN(II21461), .A(g13052) );
  INV_X1 NOT_5062( .ZN(g15148), .A(II21461) );
  INV_X1 NOT_5063( .ZN(g15151), .A(g12005) );
  INV_X1 NOT_5064( .ZN(g15161), .A(g12327) );
  INV_X1 NOT_5065( .ZN(g15170), .A(g12125) );
  INV_X1 NOT_5066( .ZN(g15174), .A(g12136) );
  INV_X1 NOT_5067( .ZN(g15175), .A(g12139) );
  INV_X1 NOT_5068( .ZN(g15176), .A(g12142) );
  INV_X1 NOT_5069( .ZN(g15177), .A(g12339) );
  INV_X1 NOT_5070( .ZN(II21476), .A(g11672) );
  INV_X1 NOT_5071( .ZN(g15179), .A(II21476) );
  INV_X1 NOT_5072( .ZN(II21479), .A(g13035) );
  INV_X1 NOT_5073( .ZN(g15182), .A(II21479) );
  INV_X1 NOT_5074( .ZN(II21482), .A(g13058) );
  INV_X1 NOT_5075( .ZN(g15185), .A(II21482) );
  INV_X1 NOT_5076( .ZN(g15188), .A(g11833) );
  INV_X1 NOT_5077( .ZN(II21488), .A(g11673) );
  INV_X1 NOT_5078( .ZN(g15198), .A(II21488) );
  INV_X1 NOT_5079( .ZN(II21491), .A(g13038) );
  INV_X1 NOT_5080( .ZN(g15201), .A(II21491) );
  INV_X1 NOT_5081( .ZN(II21494), .A(g13061) );
  INV_X1 NOT_5082( .ZN(g15204), .A(II21494) );
  INV_X1 NOT_5083( .ZN(II21497), .A(g11674) );
  INV_X1 NOT_5084( .ZN(g15207), .A(II21497) );
  INV_X1 NOT_5085( .ZN(g15210), .A(g11840) );
  INV_X1 NOT_5086( .ZN(g15220), .A(g12163) );
  INV_X1 NOT_5087( .ZN(g15221), .A(g12166) );
  INV_X1 NOT_5088( .ZN(II21505), .A(g12952) );
  INV_X1 NOT_5089( .ZN(g15222), .A(II21505) );
  INV_X1 NOT_5090( .ZN(II21508), .A(g13040) );
  INV_X1 NOT_5091( .ZN(g15225), .A(II21508) );
  INV_X1 NOT_5092( .ZN(II21511), .A(g13064) );
  INV_X1 NOT_5093( .ZN(g15228), .A(II21511) );
  INV_X1 NOT_5094( .ZN(II21514), .A(g13041) );
  INV_X1 NOT_5095( .ZN(g15231), .A(II21514) );
  INV_X1 NOT_5096( .ZN(g15236), .A(g12181) );
  INV_X1 NOT_5097( .ZN(II21520), .A(g13067) );
  INV_X1 NOT_5098( .ZN(g15237), .A(II21520) );
  INV_X1 NOT_5099( .ZN(II21523), .A(g13069) );
  INV_X1 NOT_5100( .ZN(g15240), .A(II21523) );
  INV_X1 NOT_5101( .ZN(II21531), .A(g11683) );
  INV_X1 NOT_5102( .ZN(g15248), .A(II21531) );
  INV_X1 NOT_5103( .ZN(II21534), .A(g13045) );
  INV_X1 NOT_5104( .ZN(g15251), .A(II21534) );
  INV_X1 NOT_5105( .ZN(II21537), .A(g13071) );
  INV_X1 NOT_5106( .ZN(g15254), .A(II21537) );
  INV_X1 NOT_5107( .ZN(g15260), .A(g12198) );
  INV_X1 NOT_5108( .ZN(g15261), .A(g12201) );
  INV_X1 NOT_5109( .ZN(g15262), .A(g12204) );
  INV_X1 NOT_5110( .ZN(g15263), .A(g12369) );
  INV_X1 NOT_5111( .ZN(II21548), .A(g11684) );
  INV_X1 NOT_5112( .ZN(g15265), .A(II21548) );
  INV_X1 NOT_5113( .ZN(II21551), .A(g13048) );
  INV_X1 NOT_5114( .ZN(g15268), .A(II21551) );
  INV_X1 NOT_5115( .ZN(II21554), .A(g13074) );
  INV_X1 NOT_5116( .ZN(g15271), .A(II21554) );
  INV_X1 NOT_5117( .ZN(g15274), .A(g11875) );
  INV_X1 NOT_5118( .ZN(II21560), .A(g11685) );
  INV_X1 NOT_5119( .ZN(g15284), .A(II21560) );
  INV_X1 NOT_5120( .ZN(II21563), .A(g13051) );
  INV_X1 NOT_5121( .ZN(g15287), .A(II21563) );
  INV_X1 NOT_5122( .ZN(II21566), .A(g13077) );
  INV_X1 NOT_5123( .ZN(g15290), .A(II21566) );
  INV_X1 NOT_5124( .ZN(II21569), .A(g11686) );
  INV_X1 NOT_5125( .ZN(g15293), .A(II21569) );
  INV_X1 NOT_5126( .ZN(g15296), .A(g11882) );
  INV_X1 NOT_5127( .ZN(g15306), .A(g12225) );
  INV_X1 NOT_5128( .ZN(g15307), .A(g12228) );
  INV_X1 NOT_5129( .ZN(II21577), .A(g12981) );
  INV_X1 NOT_5130( .ZN(g15308), .A(II21577) );
  INV_X1 NOT_5131( .ZN(II21580), .A(g13053) );
  INV_X1 NOT_5132( .ZN(g15311), .A(II21580) );
  INV_X1 NOT_5133( .ZN(II21583), .A(g13080) );
  INV_X1 NOT_5134( .ZN(g15314), .A(II21583) );
  INV_X1 NOT_5135( .ZN(II21586), .A(g13054) );
  INV_X1 NOT_5136( .ZN(g15317), .A(II21586) );
  INV_X1 NOT_5137( .ZN(g15322), .A(g12239) );
  INV_X1 NOT_5138( .ZN(g15323), .A(g12242) );
  INV_X1 NOT_5139( .ZN(II21595), .A(g11691) );
  INV_X1 NOT_5140( .ZN(g15326), .A(II21595) );
  INV_X4 NOT_5141( .ZN(II21598), .A(g13059) );
  INV_X4 NOT_5142( .ZN(g15329), .A(II21598) );
  INV_X1 NOT_5143( .ZN(II21601), .A(g13087) );
  INV_X1 NOT_5144( .ZN(g15332), .A(II21601) );
  INV_X1 NOT_5145( .ZN(II21609), .A(g11692) );
  INV_X1 NOT_5146( .ZN(g15340), .A(II21609) );
  INV_X1 NOT_5147( .ZN(II21612), .A(g13062) );
  INV_X1 NOT_5148( .ZN(g15343), .A(II21612) );
  INV_X1 NOT_5149( .ZN(II21615), .A(g13090) );
  INV_X1 NOT_5150( .ZN(g15346), .A(II21615) );
  INV_X1 NOT_5151( .ZN(g15352), .A(g12253) );
  INV_X1 NOT_5152( .ZN(g15353), .A(g12256) );
  INV_X1 NOT_5153( .ZN(g15354), .A(g12259) );
  INV_X1 NOT_5154( .ZN(g15355), .A(g12388) );
  INV_X1 NOT_5155( .ZN(II21626), .A(g11693) );
  INV_X1 NOT_5156( .ZN(g15357), .A(II21626) );
  INV_X1 NOT_5157( .ZN(II21629), .A(g13065) );
  INV_X1 NOT_5158( .ZN(g15360), .A(II21629) );
  INV_X1 NOT_5159( .ZN(II21632), .A(g13093) );
  INV_X1 NOT_5160( .ZN(g15363), .A(II21632) );
  INV_X1 NOT_5161( .ZN(g15366), .A(g11917) );
  INV_X1 NOT_5162( .ZN(II21638), .A(g11694) );
  INV_X1 NOT_5163( .ZN(g15376), .A(II21638) );
  INV_X1 NOT_5164( .ZN(II21641), .A(g13068) );
  INV_X1 NOT_5165( .ZN(g15379), .A(II21641) );
  INV_X1 NOT_5166( .ZN(II21644), .A(g13096) );
  INV_X1 NOT_5167( .ZN(g15382), .A(II21644) );
  INV_X1 NOT_5168( .ZN(II21647), .A(g11695) );
  INV_X1 NOT_5169( .ZN(g15385), .A(II21647) );
  INV_X1 NOT_5170( .ZN(g15390), .A(g12279) );
  INV_X1 NOT_5171( .ZN(II21655), .A(g11696) );
  INV_X1 NOT_5172( .ZN(g15393), .A(II21655) );
  INV_X1 NOT_5173( .ZN(II21658), .A(g13072) );
  INV_X1 NOT_5174( .ZN(g15396), .A(II21658) );
  INV_X1 NOT_5175( .ZN(II21661), .A(g13098) );
  INV_X1 NOT_5176( .ZN(g15399), .A(II21661) );
  INV_X1 NOT_5177( .ZN(II21666), .A(g13100) );
  INV_X1 NOT_5178( .ZN(g15404), .A(II21666) );
  INV_X1 NOT_5179( .ZN(g15408), .A(g12282) );
  INV_X1 NOT_5180( .ZN(g15409), .A(g12285) );
  INV_X1 NOT_5181( .ZN(II21674), .A(g11698) );
  INV_X1 NOT_5182( .ZN(g15412), .A(II21674) );
  INV_X1 NOT_5183( .ZN(II21677), .A(g13075) );
  INV_X1 NOT_5184( .ZN(g15415), .A(II21677) );
  INV_X1 NOT_5185( .ZN(II21680), .A(g13102) );
  INV_X1 NOT_5186( .ZN(g15418), .A(II21680) );
  INV_X1 NOT_5187( .ZN(II21688), .A(g11699) );
  INV_X1 NOT_5188( .ZN(g15426), .A(II21688) );
  INV_X1 NOT_5189( .ZN(II21691), .A(g13078) );
  INV_X1 NOT_5190( .ZN(g15429), .A(II21691) );
  INV_X1 NOT_5191( .ZN(II21694), .A(g13105) );
  INV_X1 NOT_5192( .ZN(g15432), .A(II21694) );
  INV_X1 NOT_5193( .ZN(g15438), .A(g12296) );
  INV_X1 NOT_5194( .ZN(g15439), .A(g12299) );
  INV_X1 NOT_5195( .ZN(g15440), .A(g12302) );
  INV_X1 NOT_5196( .ZN(g15441), .A(g12418) );
  INV_X1 NOT_5197( .ZN(II21705), .A(g11700) );
  INV_X1 NOT_5198( .ZN(g15443), .A(II21705) );
  INV_X1 NOT_5199( .ZN(II21708), .A(g13081) );
  INV_X1 NOT_5200( .ZN(g15446), .A(II21708) );
  INV_X1 NOT_5201( .ZN(II21711), .A(g13108) );
  INV_X1 NOT_5202( .ZN(g15449), .A(II21711) );
  INV_X1 NOT_5203( .ZN(g15458), .A(g12312) );
  INV_X1 NOT_5204( .ZN(II21720), .A(g11701) );
  INV_X1 NOT_5205( .ZN(g15461), .A(II21720) );
  INV_X1 NOT_5206( .ZN(II21723), .A(g13088) );
  INV_X1 NOT_5207( .ZN(g15464), .A(II21723) );
  INV_X1 NOT_5208( .ZN(II21726), .A(g13112) );
  INV_X1 NOT_5209( .ZN(g15467), .A(II21726) );
  INV_X1 NOT_5210( .ZN(II21730), .A(g13089) );
  INV_X1 NOT_5211( .ZN(g15471), .A(II21730) );
  INV_X1 NOT_5212( .ZN(g15474), .A(g12315) );
  INV_X1 NOT_5213( .ZN(II21736), .A(g11702) );
  INV_X1 NOT_5214( .ZN(g15477), .A(II21736) );
  INV_X1 NOT_5215( .ZN(II21739), .A(g13091) );
  INV_X1 NOT_5216( .ZN(g15480), .A(II21739) );
  INV_X1 NOT_5217( .ZN(II21742), .A(g13114) );
  INV_X1 NOT_5218( .ZN(g15483), .A(II21742) );
  INV_X1 NOT_5219( .ZN(II21747), .A(g13116) );
  INV_X1 NOT_5220( .ZN(g15488), .A(II21747) );
  INV_X1 NOT_5221( .ZN(g15492), .A(g12318) );
  INV_X1 NOT_5222( .ZN(g15493), .A(g12321) );
  INV_X1 NOT_5223( .ZN(II21755), .A(g11704) );
  INV_X1 NOT_5224( .ZN(g15496), .A(II21755) );
  INV_X1 NOT_5225( .ZN(II21758), .A(g13094) );
  INV_X1 NOT_5226( .ZN(g15499), .A(II21758) );
  INV_X1 NOT_5227( .ZN(II21761), .A(g13118) );
  INV_X1 NOT_5228( .ZN(g15502), .A(II21761) );
  INV_X1 NOT_5229( .ZN(II21769), .A(g11705) );
  INV_X1 NOT_5230( .ZN(g15510), .A(II21769) );
  INV_X1 NOT_5231( .ZN(II21772), .A(g13097) );
  INV_X1 NOT_5232( .ZN(g15513), .A(II21772) );
  INV_X1 NOT_5233( .ZN(II21775), .A(g13121) );
  INV_X1 NOT_5234( .ZN(g15516), .A(II21775) );
  INV_X1 NOT_5235( .ZN(II21780), .A(g13305) );
  INV_X1 NOT_5236( .ZN(g15521), .A(II21780) );
  INV_X1 NOT_5237( .ZN(g15524), .A(g12333) );
  INV_X1 NOT_5238( .ZN(g15525), .A(g12336) );
  INV_X1 NOT_5239( .ZN(II21787), .A(g11707) );
  INV_X1 NOT_5240( .ZN(g15528), .A(II21787) );
  INV_X1 NOT_5241( .ZN(II21790), .A(g13099) );
  INV_X1 NOT_5242( .ZN(g15531), .A(II21790) );
  INV_X1 NOT_5243( .ZN(II21793), .A(g13123) );
  INV_X1 NOT_5244( .ZN(g15534), .A(II21793) );
  INV_X1 NOT_5245( .ZN(II21796), .A(g11708) );
  INV_X1 NOT_5246( .ZN(g15537), .A(II21796) );
  INV_X1 NOT_5247( .ZN(g15544), .A(g12340) );
  INV_X1 NOT_5248( .ZN(II21803), .A(g11709) );
  INV_X1 NOT_5249( .ZN(g15547), .A(II21803) );
  INV_X1 NOT_5250( .ZN(II21806), .A(g13103) );
  INV_X1 NOT_5251( .ZN(g15550), .A(II21806) );
  INV_X1 NOT_5252( .ZN(II21809), .A(g13125) );
  INV_X1 NOT_5253( .ZN(g15553), .A(II21809) );
  INV_X1 NOT_5254( .ZN(II21813), .A(g13104) );
  INV_X1 NOT_5255( .ZN(g15557), .A(II21813) );
  INV_X1 NOT_5256( .ZN(g15560), .A(g12343) );
  INV_X1 NOT_5257( .ZN(II21819), .A(g11710) );
  INV_X1 NOT_5258( .ZN(g15563), .A(II21819) );
  INV_X1 NOT_5259( .ZN(II21822), .A(g13106) );
  INV_X1 NOT_5260( .ZN(g15566), .A(II21822) );
  INV_X1 NOT_5261( .ZN(II21825), .A(g13127) );
  INV_X1 NOT_5262( .ZN(g15569), .A(II21825) );
  INV_X1 NOT_5263( .ZN(II21830), .A(g13129) );
  INV_X1 NOT_5264( .ZN(g15574), .A(II21830) );
  INV_X1 NOT_5265( .ZN(g15578), .A(g12346) );
  INV_X1 NOT_5266( .ZN(g15579), .A(g12349) );
  INV_X1 NOT_5267( .ZN(II21838), .A(g11712) );
  INV_X1 NOT_5268( .ZN(g15582), .A(II21838) );
  INV_X1 NOT_5269( .ZN(II21841), .A(g13109) );
  INV_X1 NOT_5270( .ZN(g15585), .A(II21841) );
  INV_X1 NOT_5271( .ZN(II21844), .A(g13131) );
  INV_X1 NOT_5272( .ZN(g15588), .A(II21844) );
  INV_X1 NOT_5273( .ZN(II21852), .A(g11716) );
  INV_X1 NOT_5274( .ZN(g15596), .A(II21852) );
  INV_X1 NOT_5275( .ZN(II21855), .A(g13113) );
  INV_X1 NOT_5276( .ZN(g15599), .A(II21855) );
  INV_X1 NOT_5277( .ZN(g15602), .A(g12363) );
  INV_X1 NOT_5278( .ZN(g15603), .A(g12366) );
  INV_X1 NOT_5279( .ZN(II21862), .A(g11717) );
  INV_X1 NOT_5280( .ZN(g15606), .A(II21862) );
  INV_X1 NOT_5281( .ZN(II21865), .A(g13115) );
  INV_X1 NOT_5282( .ZN(g15609), .A(II21865) );
  INV_X1 NOT_5283( .ZN(II21868), .A(g13134) );
  INV_X1 NOT_5284( .ZN(g15612), .A(II21868) );
  INV_X1 NOT_5285( .ZN(II21871), .A(g11718) );
  INV_X1 NOT_5286( .ZN(g15615), .A(II21871) );
  INV_X1 NOT_5287( .ZN(g15622), .A(g12370) );
  INV_X1 NOT_5288( .ZN(II21878), .A(g11719) );
  INV_X1 NOT_5289( .ZN(g15625), .A(II21878) );
  INV_X1 NOT_5290( .ZN(II21881), .A(g13119) );
  INV_X1 NOT_5291( .ZN(g15628), .A(II21881) );
  INV_X1 NOT_5292( .ZN(II21884), .A(g13136) );
  INV_X1 NOT_5293( .ZN(g15631), .A(II21884) );
  INV_X1 NOT_5294( .ZN(II21888), .A(g13120) );
  INV_X1 NOT_5295( .ZN(g15635), .A(II21888) );
  INV_X1 NOT_5296( .ZN(g15638), .A(g12373) );
  INV_X1 NOT_5297( .ZN(II21894), .A(g11720) );
  INV_X1 NOT_5298( .ZN(g15641), .A(II21894) );
  INV_X1 NOT_5299( .ZN(II21897), .A(g13122) );
  INV_X1 NOT_5300( .ZN(g15644), .A(II21897) );
  INV_X1 NOT_5301( .ZN(II21900), .A(g13138) );
  INV_X1 NOT_5302( .ZN(g15647), .A(II21900) );
  INV_X1 NOT_5303( .ZN(II21905), .A(g13140) );
  INV_X1 NOT_5304( .ZN(g15652), .A(II21905) );
  INV_X1 NOT_5305( .ZN(II21908), .A(g13082) );
  INV_X1 NOT_5306( .ZN(g15655), .A(II21908) );
  INV_X1 NOT_5307( .ZN(g15659), .A(g11706) );
  INV_X1 NOT_5308( .ZN(g15665), .A(g12379) );
  INV_X1 NOT_5309( .ZN(II21918), .A(g11721) );
  INV_X1 NOT_5310( .ZN(g15667), .A(II21918) );
  INV_X1 NOT_5311( .ZN(II21923), .A(g11722) );
  INV_X1 NOT_5312( .ZN(g15672), .A(II21923) );
  INV_X1 NOT_5313( .ZN(II21926), .A(g13126) );
  INV_X1 NOT_5314( .ZN(g15675), .A(II21926) );
  INV_X1 NOT_5315( .ZN(g15678), .A(g12382) );
  INV_X1 NOT_5316( .ZN(g15679), .A(g12385) );
  INV_X4 NOT_5317( .ZN(II21933), .A(g11723) );
  INV_X4 NOT_5318( .ZN(g15682), .A(II21933) );
  INV_X1 NOT_5319( .ZN(II21936), .A(g13128) );
  INV_X1 NOT_5320( .ZN(g15685), .A(II21936) );
  INV_X1 NOT_5321( .ZN(II21939), .A(g13142) );
  INV_X1 NOT_5322( .ZN(g15688), .A(II21939) );
  INV_X1 NOT_5323( .ZN(II21942), .A(g11724) );
  INV_X1 NOT_5324( .ZN(g15691), .A(II21942) );
  INV_X1 NOT_5325( .ZN(g15698), .A(g12389) );
  INV_X1 NOT_5326( .ZN(II21949), .A(g11725) );
  INV_X1 NOT_5327( .ZN(g15701), .A(II21949) );
  INV_X1 NOT_5328( .ZN(II21952), .A(g13132) );
  INV_X1 NOT_5329( .ZN(g15704), .A(II21952) );
  INV_X1 NOT_5330( .ZN(II21955), .A(g13144) );
  INV_X1 NOT_5331( .ZN(g15707), .A(II21955) );
  INV_X1 NOT_5332( .ZN(II21959), .A(g13133) );
  INV_X1 NOT_5333( .ZN(g15711), .A(II21959) );
  INV_X1 NOT_5334( .ZN(II21962), .A(g13004) );
  INV_X1 NOT_5335( .ZN(g15714), .A(II21962) );
  INV_X1 NOT_5336( .ZN(g15722), .A(g13011) );
  INV_X1 NOT_5337( .ZN(g15724), .A(g12409) );
  INV_X1 NOT_5338( .ZN(II21974), .A(g11726) );
  INV_X1 NOT_5339( .ZN(g15726), .A(II21974) );
  INV_X1 NOT_5340( .ZN(II21979), .A(g11727) );
  INV_X1 NOT_5341( .ZN(g15731), .A(II21979) );
  INV_X1 NOT_5342( .ZN(II21982), .A(g13137) );
  INV_X1 NOT_5343( .ZN(g15734), .A(II21982) );
  INV_X1 NOT_5344( .ZN(g15737), .A(g12412) );
  INV_X1 NOT_5345( .ZN(g15738), .A(g12415) );
  INV_X1 NOT_5346( .ZN(II21989), .A(g11728) );
  INV_X1 NOT_5347( .ZN(g15741), .A(II21989) );
  INV_X1 NOT_5348( .ZN(II21992), .A(g13139) );
  INV_X1 NOT_5349( .ZN(g15744), .A(II21992) );
  INV_X1 NOT_5350( .ZN(II21995), .A(g13146) );
  INV_X1 NOT_5351( .ZN(g15747), .A(II21995) );
  INV_X1 NOT_5352( .ZN(II21998), .A(g11729) );
  INV_X1 NOT_5353( .ZN(g15750), .A(II21998) );
  INV_X1 NOT_5354( .ZN(g15762), .A(g13011) );
  INV_X1 NOT_5355( .ZN(g15764), .A(g12421) );
  INV_X1 NOT_5356( .ZN(II22014), .A(g11730) );
  INV_X1 NOT_5357( .ZN(g15766), .A(II22014) );
  INV_X1 NOT_5358( .ZN(II22019), .A(g11731) );
  INV_X1 NOT_5359( .ZN(g15771), .A(II22019) );
  INV_X1 NOT_5360( .ZN(II22022), .A(g13145) );
  INV_X1 NOT_5361( .ZN(g15774), .A(II22022) );
  INV_X1 NOT_5362( .ZN(II22025), .A(g11617) );
  INV_X1 NOT_5363( .ZN(g15777), .A(II22025) );
  INV_X1 NOT_5364( .ZN(g15790), .A(g13011) );
  INV_X1 NOT_5365( .ZN(g15792), .A(g12426) );
  INV_X1 NOT_5366( .ZN(II22044), .A(g11733) );
  INV_X1 NOT_5367( .ZN(g15794), .A(II22044) );
  INV_X1 NOT_5368( .ZN(g15800), .A(g12909) );
  INV_X1 NOT_5369( .ZN(g15813), .A(g13011) );
  INV_X1 NOT_5370( .ZN(g15859), .A(g13378) );
  INV_X1 NOT_5371( .ZN(II22120), .A(g12909) );
  INV_X1 NOT_5372( .ZN(g15876), .A(II22120) );
  INV_X1 NOT_5373( .ZN(g15880), .A(g11624) );
  INV_X1 NOT_5374( .ZN(g15890), .A(g11600) );
  INV_X1 NOT_5375( .ZN(g15904), .A(g11644) );
  INV_X1 NOT_5376( .ZN(g15913), .A(g11647) );
  INV_X1 NOT_5377( .ZN(g15923), .A(g11630) );
  INV_X1 NOT_5378( .ZN(g15933), .A(g11663) );
  INV_X1 NOT_5379( .ZN(g15942), .A(g11666) );
  INV_X1 NOT_5380( .ZN(g15952), .A(g11653) );
  INV_X1 NOT_5381( .ZN(g15962), .A(g11675) );
  INV_X1 NOT_5382( .ZN(g15971), .A(g11678) );
  INV_X1 NOT_5383( .ZN(g15981), .A(g11687) );
  INV_X1 NOT_5384( .ZN(II22163), .A(g12433) );
  INV_X1 NOT_5385( .ZN(g15989), .A(II22163) );
  INV_X1 NOT_5386( .ZN(g15991), .A(g12548) );
  INV_X1 NOT_5387( .ZN(g15994), .A(g12555) );
  INV_X1 NOT_5388( .ZN(g15997), .A(g12561) );
  INV_X1 NOT_5389( .ZN(g16001), .A(g12601) );
  INV_X1 NOT_5390( .ZN(g16002), .A(g12604) );
  INV_X1 NOT_5391( .ZN(g16005), .A(g12608) );
  INV_X1 NOT_5392( .ZN(g16007), .A(g12647) );
  INV_X1 NOT_5393( .ZN(g16011), .A(g12651) );
  INV_X1 NOT_5394( .ZN(g16012), .A(g12654) );
  INV_X1 NOT_5395( .ZN(g16013), .A(g12692) );
  INV_X1 NOT_5396( .ZN(g16014), .A(g12695) );
  INV_X1 NOT_5397( .ZN(g16023), .A(g12699) );
  INV_X1 NOT_5398( .ZN(g16024), .A(g12702) );
  INV_X1 NOT_5399( .ZN(g16025), .A(g12705) );
  INV_X1 NOT_5400( .ZN(g16026), .A(g12708) );
  INV_X1 NOT_5401( .ZN(g16027), .A(g12744) );
  INV_X1 NOT_5402( .ZN(g16034), .A(g12749) );
  INV_X1 NOT_5403( .ZN(g16035), .A(g12752) );
  INV_X1 NOT_5404( .ZN(g16039), .A(g12756) );
  INV_X1 NOT_5405( .ZN(g16040), .A(g12759) );
  INV_X1 NOT_5406( .ZN(g16041), .A(g12762) );
  INV_X1 NOT_5407( .ZN(g16042), .A(g12765) );
  INV_X1 NOT_5408( .ZN(g16043), .A(g12769) );
  INV_X1 NOT_5409( .ZN(g16044), .A(g12772) );
  INV_X1 NOT_5410( .ZN(g16054), .A(g12783) );
  INV_X1 NOT_5411( .ZN(g16055), .A(g12786) );
  INV_X1 NOT_5412( .ZN(g16056), .A(g12791) );
  INV_X1 NOT_5413( .ZN(g16057), .A(g12794) );
  INV_X1 NOT_5414( .ZN(g16061), .A(g12798) );
  INV_X1 NOT_5415( .ZN(g16062), .A(g12801) );
  INV_X1 NOT_5416( .ZN(g16063), .A(g12804) );
  INV_X1 NOT_5417( .ZN(g16064), .A(g12808) );
  INV_X1 NOT_5418( .ZN(g16065), .A(g12811) );
  INV_X1 NOT_5419( .ZN(g16075), .A(g11861) );
  INV_X1 NOT_5420( .ZN(g16088), .A(g12816) );
  INV_X1 NOT_5421( .ZN(g16090), .A(g12822) );
  INV_X1 NOT_5422( .ZN(g16091), .A(g12825) );
  INV_X1 NOT_5423( .ZN(g16092), .A(g12830) );
  INV_X1 NOT_5424( .ZN(g16093), .A(g12833) );
  INV_X1 NOT_5425( .ZN(g16097), .A(g12837) );
  INV_X1 NOT_5426( .ZN(g16098), .A(g12840) );
  INV_X1 NOT_5427( .ZN(g16099), .A(g12844) );
  INV_X1 NOT_5428( .ZN(g16113), .A(g11903) );
  INV_X1 NOT_5429( .ZN(g16126), .A(g12854) );
  INV_X1 NOT_5430( .ZN(g16128), .A(g12860) );
  INV_X1 NOT_5431( .ZN(g16129), .A(g12863) );
  INV_X1 NOT_5432( .ZN(g16130), .A(g12868) );
  INV_X1 NOT_5433( .ZN(g16131), .A(g12871) );
  INV_X1 NOT_5434( .ZN(g16142), .A(g13057) );
  INV_X1 NOT_5435( .ZN(g16154), .A(g12194) );
  INV_X1 NOT_5436( .ZN(g16164), .A(g11953) );
  INV_X1 NOT_5437( .ZN(g16177), .A(g12895) );
  INV_X1 NOT_5438( .ZN(g16179), .A(g12901) );
  INV_X1 NOT_5439( .ZN(g16180), .A(g12904) );
  INV_X1 NOT_5440( .ZN(g16189), .A(g13043) );
  INV_X1 NOT_5441( .ZN(g16201), .A(g13073) );
  INV_X1 NOT_5442( .ZN(g16213), .A(g12249) );
  INV_X1 NOT_5443( .ZN(g16223), .A(g12006) );
  INV_X1 NOT_5444( .ZN(g16236), .A(g12935) );
  INV_X1 NOT_5445( .ZN(g16243), .A(g13033) );
  INV_X1 NOT_5446( .ZN(g16254), .A(g13060) );
  INV_X1 NOT_5447( .ZN(g16266), .A(g13092) );
  INV_X1 NOT_5448( .ZN(g16278), .A(g12292) );
  INV_X1 NOT_5449( .ZN(g16287), .A(g12962) );
  INV_X1 NOT_5450( .ZN(g16293), .A(g13025) );
  INV_X1 NOT_5451( .ZN(II22382), .A(g520) );
  INV_X1 NOT_5452( .ZN(g16297), .A(II22382) );
  INV_X1 NOT_5453( .ZN(g16302), .A(g13046) );
  INV_X1 NOT_5454( .ZN(g16313), .A(g13076) );
  INV_X1 NOT_5455( .ZN(g16325), .A(g13107) );
  INV_X1 NOT_5456( .ZN(g16337), .A(g12328) );
  INV_X1 NOT_5457( .ZN(g16351), .A(g13036) );
  INV_X1 NOT_5458( .ZN(II22414), .A(g1206) );
  INV_X1 NOT_5459( .ZN(g16355), .A(II22414) );
  INV_X1 NOT_5460( .ZN(g16360), .A(g13063) );
  INV_X1 NOT_5461( .ZN(g16371), .A(g13095) );
  INV_X1 NOT_5462( .ZN(g16395), .A(g13049) );
  INV_X1 NOT_5463( .ZN(II22444), .A(g1900) );
  INV_X1 NOT_5464( .ZN(g16399), .A(II22444) );
  INV_X1 NOT_5465( .ZN(g16404), .A(g13079) );
  INV_X1 NOT_5466( .ZN(g16433), .A(g13066) );
  INV_X1 NOT_5467( .ZN(II22475), .A(g2594) );
  INV_X1 NOT_5468( .ZN(g16437), .A(II22475) );
  INV_X1 NOT_5469( .ZN(g16466), .A(g12017) );
  INV_X1 NOT_5470( .ZN(II22503), .A(g13598) );
  INV_X1 NOT_5471( .ZN(g16467), .A(II22503) );
  INV_X1 NOT_5472( .ZN(II22506), .A(g13624) );
  INV_X1 NOT_5473( .ZN(g16468), .A(II22506) );
  INV_X1 NOT_5474( .ZN(II22509), .A(g13610) );
  INV_X1 NOT_5475( .ZN(g16469), .A(II22509) );
  INV_X1 NOT_5476( .ZN(II22512), .A(g13635) );
  INV_X1 NOT_5477( .ZN(g16470), .A(II22512) );
  INV_X1 NOT_5478( .ZN(II22515), .A(g13620) );
  INV_X1 NOT_5479( .ZN(g16471), .A(II22515) );
  INV_X1 NOT_5480( .ZN(II22518), .A(g13647) );
  INV_X1 NOT_5481( .ZN(g16472), .A(II22518) );
  INV_X1 NOT_5482( .ZN(II22521), .A(g13632) );
  INV_X1 NOT_5483( .ZN(g16473), .A(II22521) );
  INV_X1 NOT_5484( .ZN(II22524), .A(g13673) );
  INV_X1 NOT_5485( .ZN(g16474), .A(II22524) );
  INV_X1 NOT_5486( .ZN(II22527), .A(g13469) );
  INV_X1 NOT_5487( .ZN(g16475), .A(II22527) );
  INV_X1 NOT_5488( .ZN(II22530), .A(g14774) );
  INV_X1 NOT_5489( .ZN(g16476), .A(II22530) );
  INV_X1 NOT_5490( .ZN(II22533), .A(g14795) );
  INV_X1 NOT_5491( .ZN(g16477), .A(II22533) );
  INV_X1 NOT_5492( .ZN(II22536), .A(g14829) );
  INV_X1 NOT_5493( .ZN(g16478), .A(II22536) );
  INV_X1 NOT_5494( .ZN(II22539), .A(g14882) );
  INV_X1 NOT_5495( .ZN(g16479), .A(II22539) );
  INV_X1 NOT_5496( .ZN(II22542), .A(g14954) );
  INV_X1 NOT_5497( .ZN(g16480), .A(II22542) );
  INV_X1 NOT_5498( .ZN(II22545), .A(g15018) );
  INV_X1 NOT_5499( .ZN(g16481), .A(II22545) );
  INV_X1 NOT_5500( .ZN(II22548), .A(g14718) );
  INV_X1 NOT_5501( .ZN(g16482), .A(II22548) );
  INV_X1 NOT_5502( .ZN(II22551), .A(g14745) );
  INV_X1 NOT_5503( .ZN(g16483), .A(II22551) );
  INV_X1 NOT_5504( .ZN(II22554), .A(g14765) );
  INV_X1 NOT_5505( .ZN(g16484), .A(II22554) );
  INV_X1 NOT_5506( .ZN(II22557), .A(g14775) );
  INV_X1 NOT_5507( .ZN(g16485), .A(II22557) );
  INV_X1 NOT_5508( .ZN(II22560), .A(g14796) );
  INV_X1 NOT_5509( .ZN(g16486), .A(II22560) );
  INV_X1 NOT_5510( .ZN(II22563), .A(g14830) );
  INV_X1 NOT_5511( .ZN(g16487), .A(II22563) );
  INV_X1 NOT_5512( .ZN(II22566), .A(g14883) );
  INV_X1 NOT_5513( .ZN(g16488), .A(II22566) );
  INV_X1 NOT_5514( .ZN(II22569), .A(g14955) );
  INV_X1 NOT_5515( .ZN(g16489), .A(II22569) );
  INV_X1 NOT_5516( .ZN(II22572), .A(g15019) );
  INV_X1 NOT_5517( .ZN(g16490), .A(II22572) );
  INV_X1 NOT_5518( .ZN(II22575), .A(g15092) );
  INV_X1 NOT_5519( .ZN(g16491), .A(II22575) );
  INV_X1 NOT_5520( .ZN(II22578), .A(g14746) );
  INV_X1 NOT_5521( .ZN(g16492), .A(II22578) );
  INV_X1 NOT_5522( .ZN(II22581), .A(g14766) );
  INV_X1 NOT_5523( .ZN(g16493), .A(II22581) );
  INV_X1 NOT_5524( .ZN(II22584), .A(g15989) );
  INV_X1 NOT_5525( .ZN(g16494), .A(II22584) );
  INV_X1 NOT_5526( .ZN(II22587), .A(g14684) );
  INV_X1 NOT_5527( .ZN(g16495), .A(II22587) );
  INV_X1 NOT_5528( .ZN(II22590), .A(g13863) );
  INV_X1 NOT_5529( .ZN(g16496), .A(II22590) );
  INV_X1 NOT_5530( .ZN(II22593), .A(g15876) );
  INV_X1 NOT_5531( .ZN(g16497), .A(II22593) );
  INV_X1 NOT_5532( .ZN(g16501), .A(g14158) );
  INV_X1 NOT_5533( .ZN(II22599), .A(g14966) );
  INV_X1 NOT_5534( .ZN(g16506), .A(II22599) );
  INV_X1 NOT_5535( .ZN(g16507), .A(g14186) );
  INV_X1 NOT_5536( .ZN(II22604), .A(g15080) );
  INV_X1 NOT_5537( .ZN(g16514), .A(II22604) );
  INV_X4 NOT_5538( .ZN(g16515), .A(g14244) );
  INV_X4 NOT_5539( .ZN(g16523), .A(g14273) );
  INV_X1 NOT_5540( .ZN(II22611), .A(g15055) );
  INV_X1 NOT_5541( .ZN(g16528), .A(II22611) );
  INV_X1 NOT_5542( .ZN(g16529), .A(g14301) );
  INV_X1 NOT_5543( .ZN(II22618), .A(g14630) );
  INV_X1 NOT_5544( .ZN(g16540), .A(II22618) );
  INV_X1 NOT_5545( .ZN(g16543), .A(g14347) );
  INV_X1 NOT_5546( .ZN(g16546), .A(g14366) );
  INV_X1 NOT_5547( .ZN(g16554), .A(g14395) );
  INV_X1 NOT_5548( .ZN(II22626), .A(g15151) );
  INV_X1 NOT_5549( .ZN(g16559), .A(II22626) );
  INV_X1 NOT_5550( .ZN(g16560), .A(g14423) );
  INV_X1 NOT_5551( .ZN(II22640), .A(g14650) );
  INV_X1 NOT_5552( .ZN(g16572), .A(II22640) );
  INV_X1 NOT_5553( .ZN(g16575), .A(g14459) );
  INV_X1 NOT_5554( .ZN(g16578), .A(g14478) );
  INV_X1 NOT_5555( .ZN(g16586), .A(g14507) );
  INV_X1 NOT_5556( .ZN(II22651), .A(g14677) );
  INV_X1 NOT_5557( .ZN(g16596), .A(II22651) );
  INV_X1 NOT_5558( .ZN(g16599), .A(g14546) );
  INV_X1 NOT_5559( .ZN(g16602), .A(g14565) );
  INV_X1 NOT_5560( .ZN(II22657), .A(g14657) );
  INV_X1 NOT_5561( .ZN(g16608), .A(II22657) );
  INV_X1 NOT_5562( .ZN(II22663), .A(g14711) );
  INV_X1 NOT_5563( .ZN(g16616), .A(II22663) );
  INV_X1 NOT_5564( .ZN(g16619), .A(g14601) );
  INV_X1 NOT_5565( .ZN(II22667), .A(g14642) );
  INV_X1 NOT_5566( .ZN(g16622), .A(II22667) );
  INV_X1 NOT_5567( .ZN(II22671), .A(g14691) );
  INV_X1 NOT_5568( .ZN(g16626), .A(II22671) );
  INV_X1 NOT_5569( .ZN(II22676), .A(g14630) );
  INV_X1 NOT_5570( .ZN(g16633), .A(II22676) );
  INV_X1 NOT_5571( .ZN(II22679), .A(g14669) );
  INV_X1 NOT_5572( .ZN(g16636), .A(II22679) );
  INV_X1 NOT_5573( .ZN(II22683), .A(g14725) );
  INV_X1 NOT_5574( .ZN(g16640), .A(II22683) );
  INV_X1 NOT_5575( .ZN(II22687), .A(g14650) );
  INV_X1 NOT_5576( .ZN(g16644), .A(II22687) );
  INV_X1 NOT_5577( .ZN(II22690), .A(g14703) );
  INV_X1 NOT_5578( .ZN(g16647), .A(II22690) );
  INV_X1 NOT_5579( .ZN(II22694), .A(g14753) );
  INV_X1 NOT_5580( .ZN(g16651), .A(II22694) );
  INV_X1 NOT_5581( .ZN(II22699), .A(g14677) );
  INV_X1 NOT_5582( .ZN(g16656), .A(II22699) );
  INV_X1 NOT_5583( .ZN(II22702), .A(g14737) );
  INV_X1 NOT_5584( .ZN(g16659), .A(II22702) );
  INV_X1 NOT_5585( .ZN(g16665), .A(g14776) );
  INV_X1 NOT_5586( .ZN(II22715), .A(g14711) );
  INV_X1 NOT_5587( .ZN(g16673), .A(II22715) );
  INV_X1 NOT_5588( .ZN(II22718), .A(g14657) );
  INV_X1 NOT_5589( .ZN(g16676), .A(II22718) );
  INV_X1 NOT_5590( .ZN(g16682), .A(g14797) );
  INV_X1 NOT_5591( .ZN(g16686), .A(g14811) );
  INV_X1 NOT_5592( .ZN(II22726), .A(g14642) );
  INV_X1 NOT_5593( .ZN(g16694), .A(II22726) );
  INV_X1 NOT_5594( .ZN(g16697), .A(g14837) );
  INV_X1 NOT_5595( .ZN(II22730), .A(g14691) );
  INV_X1 NOT_5596( .ZN(g16702), .A(II22730) );
  INV_X1 NOT_5597( .ZN(g16708), .A(g14849) );
  INV_X1 NOT_5598( .ZN(g16712), .A(g14863) );
  INV_X1 NOT_5599( .ZN(II22737), .A(g14630) );
  INV_X1 NOT_5600( .ZN(g16719), .A(II22737) );
  INV_X1 NOT_5601( .ZN(g16722), .A(g14895) );
  INV_X1 NOT_5602( .ZN(II22741), .A(g14669) );
  INV_X1 NOT_5603( .ZN(g16725), .A(II22741) );
  INV_X1 NOT_5604( .ZN(g16728), .A(g14910) );
  INV_X1 NOT_5605( .ZN(II22745), .A(g14725) );
  INV_X1 NOT_5606( .ZN(g16733), .A(II22745) );
  INV_X1 NOT_5607( .ZN(g16739), .A(g14922) );
  INV_X1 NOT_5608( .ZN(g16743), .A(g14936) );
  INV_X1 NOT_5609( .ZN(g16749), .A(g15782) );
  INV_X1 NOT_5610( .ZN(II22752), .A(g14657) );
  INV_X1 NOT_5611( .ZN(g16758), .A(II22752) );
  INV_X1 NOT_5612( .ZN(II22755), .A(g14650) );
  INV_X1 NOT_5613( .ZN(g16761), .A(II22755) );
  INV_X1 NOT_5614( .ZN(g16764), .A(g14976) );
  INV_X1 NOT_5615( .ZN(II22759), .A(g14703) );
  INV_X1 NOT_5616( .ZN(g16767), .A(II22759) );
  INV_X1 NOT_5617( .ZN(g16770), .A(g14991) );
  INV_X1 NOT_5618( .ZN(II22763), .A(g14753) );
  INV_X1 NOT_5619( .ZN(g16775), .A(II22763) );
  INV_X1 NOT_5620( .ZN(g16781), .A(g15003) );
  INV_X1 NOT_5621( .ZN(II22768), .A(g14691) );
  INV_X1 NOT_5622( .ZN(g16785), .A(II22768) );
  INV_X1 NOT_5623( .ZN(II22771), .A(g14677) );
  INV_X1 NOT_5624( .ZN(g16788), .A(II22771) );
  INV_X1 NOT_5625( .ZN(g16791), .A(g15065) );
  INV_X1 NOT_5626( .ZN(II22775), .A(g14737) );
  INV_X1 NOT_5627( .ZN(g16794), .A(II22775) );
  INV_X1 NOT_5628( .ZN(g16797), .A(g15080) );
  INV_X1 NOT_5629( .ZN(g16804), .A(g15803) );
  INV_X1 NOT_5630( .ZN(g16809), .A(g15842) );
  INV_X1 NOT_5631( .ZN(II22783), .A(g13572) );
  INV_X1 NOT_5632( .ZN(g16813), .A(II22783) );
  INV_X1 NOT_5633( .ZN(II22786), .A(g14725) );
  INV_X1 NOT_5634( .ZN(g16814), .A(II22786) );
  INV_X1 NOT_5635( .ZN(II22789), .A(g14711) );
  INV_X1 NOT_5636( .ZN(g16817), .A(II22789) );
  INV_X1 NOT_5637( .ZN(g16820), .A(g15161) );
  INV_X1 NOT_5638( .ZN(g16825), .A(g15855) );
  INV_X1 NOT_5639( .ZN(II22797), .A(g14165) );
  INV_X1 NOT_5640( .ZN(g16830), .A(II22797) );
  INV_X1 NOT_5641( .ZN(II22800), .A(g13581) );
  INV_X1 NOT_5642( .ZN(g16831), .A(II22800) );
  INV_X1 NOT_5643( .ZN(II22803), .A(g14753) );
  INV_X1 NOT_5644( .ZN(g16832), .A(II22803) );
  INV_X1 NOT_5645( .ZN(g16836), .A(g15818) );
  INV_X1 NOT_5646( .ZN(g16840), .A(g15878) );
  INV_X1 NOT_5647( .ZN(II22810), .A(g14280) );
  INV_X1 NOT_5648( .ZN(g16842), .A(II22810) );
  INV_X1 NOT_5649( .ZN(II22813), .A(g13601) );
  INV_X1 NOT_5650( .ZN(g16843), .A(II22813) );
  INV_X1 NOT_5651( .ZN(g16846), .A(g15903) );
  INV_X1 NOT_5652( .ZN(II22820), .A(g14402) );
  INV_X1 NOT_5653( .ZN(g16848), .A(II22820) );
  INV_X1 NOT_5654( .ZN(II22823), .A(g13613) );
  INV_X1 NOT_5655( .ZN(g16849), .A(II22823) );
  INV_X1 NOT_5656( .ZN(II22828), .A(g14514) );
  INV_X1 NOT_5657( .ZN(g16852), .A(II22828) );
  INV_X1 NOT_5658( .ZN(II22836), .A(g13571) );
  INV_X1 NOT_5659( .ZN(g16858), .A(II22836) );
  INV_X1 NOT_5660( .ZN(II22842), .A(g13580) );
  INV_X1 NOT_5661( .ZN(g16862), .A(II22842) );
  INV_X1 NOT_5662( .ZN(II22845), .A(g13579) );
  INV_X1 NOT_5663( .ZN(g16863), .A(II22845) );
  INV_X1 NOT_5664( .ZN(g16867), .A(g13589) );
  INV_X1 NOT_5665( .ZN(II22852), .A(g13600) );
  INV_X1 NOT_5666( .ZN(g16877), .A(II22852) );
  INV_X1 NOT_5667( .ZN(II22855), .A(g13588) );
  INV_X1 NOT_5668( .ZN(g16878), .A(II22855) );
  INV_X1 NOT_5669( .ZN(II22860), .A(g14885) );
  INV_X1 NOT_5670( .ZN(g16881), .A(II22860) );
  INV_X1 NOT_5671( .ZN(g16884), .A(g13589) );
  INV_X1 NOT_5672( .ZN(g16895), .A(g13589) );
  INV_X1 NOT_5673( .ZN(II22866), .A(g13612) );
  INV_X1 NOT_5674( .ZN(g16905), .A(II22866) );
  INV_X1 NOT_5675( .ZN(II22869), .A(g13608) );
  INV_X1 NOT_5676( .ZN(g16906), .A(II22869) );
  INV_X1 NOT_5677( .ZN(II22875), .A(g14966) );
  INV_X1 NOT_5678( .ZN(g16910), .A(II22875) );
  INV_X1 NOT_5679( .ZN(g16913), .A(g13589) );
  INV_X1 NOT_5680( .ZN(g16924), .A(g13589) );
  INV_X1 NOT_5681( .ZN(II22881), .A(g13622) );
  INV_X1 NOT_5682( .ZN(g16934), .A(II22881) );
  INV_X1 NOT_5683( .ZN(II22893), .A(g15055) );
  INV_X1 NOT_5684( .ZN(g16940), .A(II22893) );
  INV_X1 NOT_5685( .ZN(g16943), .A(g13589) );
  INV_X1 NOT_5686( .ZN(g16954), .A(g13589) );
  INV_X1 NOT_5687( .ZN(II22912), .A(g15151) );
  INV_X1 NOT_5688( .ZN(g16971), .A(II22912) );
  INV_X1 NOT_5689( .ZN(g16974), .A(g13589) );
  INV_X1 NOT_5690( .ZN(g17029), .A(g14685) );
  INV_X1 NOT_5691( .ZN(g17057), .A(g13519) );
  INV_X1 NOT_5692( .ZN(g17063), .A(g14719) );
  INV_X1 NOT_5693( .ZN(g17092), .A(g13530) );
  INV_X1 NOT_5694( .ZN(g17098), .A(g14747) );
  INV_X1 NOT_5695( .ZN(g17130), .A(g13541) );
  INV_X1 NOT_5696( .ZN(g17136), .A(g14768) );
  INV_X1 NOT_5697( .ZN(g17157), .A(g13552) );
  INV_X1 NOT_5698( .ZN(II23253), .A(g13741) );
  INV_X1 NOT_5699( .ZN(g17189), .A(II23253) );
  INV_X1 NOT_5700( .ZN(II23274), .A(g13741) );
  INV_X1 NOT_5701( .ZN(g17200), .A(II23274) );
  INV_X1 NOT_5702( .ZN(g17203), .A(g13568) );
  INV_X1 NOT_5703( .ZN(II23287), .A(g13741) );
  INV_X1 NOT_5704( .ZN(g17207), .A(II23287) );
  INV_X1 NOT_5705( .ZN(g17208), .A(g13576) );
  INV_X1 NOT_5706( .ZN(II23292), .A(g13741) );
  INV_X1 NOT_5707( .ZN(g17212), .A(II23292) );
  INV_X1 NOT_5708( .ZN(g17214), .A(g13585) );
  INV_X1 NOT_5709( .ZN(g17217), .A(g13605) );
  INV_X1 NOT_5710( .ZN(II23309), .A(g16132) );
  INV_X1 NOT_5711( .ZN(g17227), .A(II23309) );
  INV_X1 NOT_5712( .ZN(II23314), .A(g15720) );
  INV_X1 NOT_5713( .ZN(g17230), .A(II23314) );
  INV_X1 NOT_5714( .ZN(II23317), .A(g16181) );
  INV_X1 NOT_5715( .ZN(g17233), .A(II23317) );
  INV_X1 NOT_5716( .ZN(II23323), .A(g15664) );
  INV_X1 NOT_5717( .ZN(g17237), .A(II23323) );
  INV_X1 NOT_5718( .ZN(II23326), .A(g15758) );
  INV_X4 NOT_5719( .ZN(g17240), .A(II23326) );
  INV_X1 NOT_5720( .ZN(II23329), .A(g15760) );
  INV_X1 NOT_5721( .ZN(g17243), .A(II23329) );
  INV_X1 NOT_5722( .ZN(II23335), .A(g16412) );
  INV_X1 NOT_5723( .ZN(g17249), .A(II23335) );
  INV_X1 NOT_5724( .ZN(II23338), .A(g15721) );
  INV_X1 NOT_5725( .ZN(g17252), .A(II23338) );
  INV_X1 NOT_5726( .ZN(II23341), .A(g15784) );
  INV_X1 NOT_5727( .ZN(g17255), .A(II23341) );
  INV_X1 NOT_5728( .ZN(g17258), .A(g16053) );
  INV_X1 NOT_5729( .ZN(II23345), .A(g15723) );
  INV_X1 NOT_5730( .ZN(g17259), .A(II23345) );
  INV_X1 NOT_5731( .ZN(II23348), .A(g15786) );
  INV_X1 NOT_5732( .ZN(g17262), .A(II23348) );
  INV_X1 NOT_5733( .ZN(II23351), .A(g15788) );
  INV_X1 NOT_5734( .ZN(g17265), .A(II23351) );
  INV_X1 NOT_5735( .ZN(II23358), .A(g16442) );
  INV_X1 NOT_5736( .ZN(g17272), .A(II23358) );
  INV_X1 NOT_5737( .ZN(II23361), .A(g15759) );
  INV_X1 NOT_5738( .ZN(g17275), .A(II23361) );
  INV_X1 NOT_5739( .ZN(II23364), .A(g15805) );
  INV_X1 NOT_5740( .ZN(g17278), .A(II23364) );
  INV_X1 NOT_5741( .ZN(g17281), .A(g16081) );
  INV_X1 NOT_5742( .ZN(II23368), .A(g16446) );
  INV_X1 NOT_5743( .ZN(g17282), .A(II23368) );
  INV_X1 NOT_5744( .ZN(II23371), .A(g15761) );
  INV_X1 NOT_5745( .ZN(g17285), .A(II23371) );
  INV_X1 NOT_5746( .ZN(II23374), .A(g15807) );
  INV_X1 NOT_5747( .ZN(g17288), .A(II23374) );
  INV_X1 NOT_5748( .ZN(II23377), .A(g15763) );
  INV_X1 NOT_5749( .ZN(g17291), .A(II23377) );
  INV_X1 NOT_5750( .ZN(II23380), .A(g15809) );
  INV_X1 NOT_5751( .ZN(g17294), .A(II23380) );
  INV_X1 NOT_5752( .ZN(II23383), .A(g15811) );
  INV_X1 NOT_5753( .ZN(g17297), .A(II23383) );
  INV_X1 NOT_5754( .ZN(II23386), .A(g13469) );
  INV_X1 NOT_5755( .ZN(g17300), .A(II23386) );
  INV_X1 NOT_5756( .ZN(II23392), .A(g13476) );
  INV_X1 NOT_5757( .ZN(g17304), .A(II23392) );
  INV_X1 NOT_5758( .ZN(II23395), .A(g15785) );
  INV_X1 NOT_5759( .ZN(g17307), .A(II23395) );
  INV_X1 NOT_5760( .ZN(II23398), .A(g15820) );
  INV_X1 NOT_5761( .ZN(g17310), .A(II23398) );
  INV_X1 NOT_5762( .ZN(g17313), .A(g16109) );
  INV_X1 NOT_5763( .ZN(g17314), .A(g16110) );
  INV_X1 NOT_5764( .ZN(II23403), .A(g13478) );
  INV_X1 NOT_5765( .ZN(g17315), .A(II23403) );
  INV_X1 NOT_5766( .ZN(II23406), .A(g15787) );
  INV_X1 NOT_5767( .ZN(g17318), .A(II23406) );
  INV_X2 NOT_5768( .ZN(II23409), .A(g15822) );
  INV_X2 NOT_5769( .ZN(g17321), .A(II23409) );
  INV_X1 NOT_5770( .ZN(II23412), .A(g13482) );
  INV_X1 NOT_5771( .ZN(g17324), .A(II23412) );
  INV_X1 NOT_5772( .ZN(II23415), .A(g15789) );
  INV_X1 NOT_5773( .ZN(g17327), .A(II23415) );
  INV_X1 NOT_5774( .ZN(II23418), .A(g15824) );
  INV_X1 NOT_5775( .ZN(g17330), .A(II23418) );
  INV_X1 NOT_5776( .ZN(II23421), .A(g15791) );
  INV_X1 NOT_5777( .ZN(g17333), .A(II23421) );
  INV_X1 NOT_5778( .ZN(II23424), .A(g15826) );
  INV_X1 NOT_5779( .ZN(g17336), .A(II23424) );
  INV_X1 NOT_5780( .ZN(II23430), .A(g13494) );
  INV_X1 NOT_5781( .ZN(g17342), .A(II23430) );
  INV_X1 NOT_5782( .ZN(II23433), .A(g15806) );
  INV_X1 NOT_5783( .ZN(g17345), .A(II23433) );
  INV_X1 NOT_5784( .ZN(II23436), .A(g15832) );
  INV_X1 NOT_5785( .ZN(g17348), .A(II23436) );
  INV_X1 NOT_5786( .ZN(g17351), .A(g16152) );
  INV_X1 NOT_5787( .ZN(II23442), .A(g13495) );
  INV_X1 NOT_5788( .ZN(g17354), .A(II23442) );
  INV_X1 NOT_5789( .ZN(II23445), .A(g15808) );
  INV_X1 NOT_5790( .ZN(g17357), .A(II23445) );
  INV_X1 NOT_5791( .ZN(II23448), .A(g15834) );
  INV_X1 NOT_5792( .ZN(g17360), .A(II23448) );
  INV_X1 NOT_5793( .ZN(II23451), .A(g13497) );
  INV_X1 NOT_5794( .ZN(g17363), .A(II23451) );
  INV_X1 NOT_5795( .ZN(II23454), .A(g15810) );
  INV_X1 NOT_5796( .ZN(g17366), .A(II23454) );
  INV_X1 NOT_5797( .ZN(II23457), .A(g15836) );
  INV_X1 NOT_5798( .ZN(g17369), .A(II23457) );
  INV_X1 NOT_5799( .ZN(II23460), .A(g13501) );
  INV_X1 NOT_5800( .ZN(g17372), .A(II23460) );
  INV_X1 NOT_5801( .ZN(II23463), .A(g15812) );
  INV_X1 NOT_5802( .ZN(g17375), .A(II23463) );
  INV_X1 NOT_5803( .ZN(II23466), .A(g15838) );
  INV_X1 NOT_5804( .ZN(g17378), .A(II23466) );
  INV_X1 NOT_5805( .ZN(II23472), .A(g13510) );
  INV_X1 NOT_5806( .ZN(g17384), .A(II23472) );
  INV_X1 NOT_5807( .ZN(II23475), .A(g15821) );
  INV_X1 NOT_5808( .ZN(g17387), .A(II23475) );
  INV_X1 NOT_5809( .ZN(II23478), .A(g15844) );
  INV_X1 NOT_5810( .ZN(g17390), .A(II23478) );
  INV_X1 NOT_5811( .ZN(g17394), .A(g16197) );
  INV_X1 NOT_5812( .ZN(II23487), .A(g13511) );
  INV_X1 NOT_5813( .ZN(g17399), .A(II23487) );
  INV_X1 NOT_5814( .ZN(II23490), .A(g15823) );
  INV_X1 NOT_5815( .ZN(g17402), .A(II23490) );
  INV_X1 NOT_5816( .ZN(II23493), .A(g15846) );
  INV_X1 NOT_5817( .ZN(g17405), .A(II23493) );
  INV_X1 NOT_5818( .ZN(II23498), .A(g13512) );
  INV_X1 NOT_5819( .ZN(g17410), .A(II23498) );
  INV_X1 NOT_5820( .ZN(II23501), .A(g15825) );
  INV_X1 NOT_5821( .ZN(g17413), .A(II23501) );
  INV_X1 NOT_5822( .ZN(II23504), .A(g15848) );
  INV_X1 NOT_5823( .ZN(g17416), .A(II23504) );
  INV_X1 NOT_5824( .ZN(II23507), .A(g13514) );
  INV_X1 NOT_5825( .ZN(g17419), .A(II23507) );
  INV_X1 NOT_5826( .ZN(II23510), .A(g15827) );
  INV_X1 NOT_5827( .ZN(g17422), .A(II23510) );
  INV_X1 NOT_5828( .ZN(II23513), .A(g15850) );
  INV_X1 NOT_5829( .ZN(g17425), .A(II23513) );
  INV_X1 NOT_5830( .ZN(II23518), .A(g15856) );
  INV_X1 NOT_5831( .ZN(g17430), .A(II23518) );
  INV_X1 NOT_5832( .ZN(II23521), .A(g13518) );
  INV_X1 NOT_5833( .ZN(g17433), .A(II23521) );
  INV_X1 NOT_5834( .ZN(II23524), .A(g15833) );
  INV_X1 NOT_5835( .ZN(g17436), .A(II23524) );
  INV_X1 NOT_5836( .ZN(II23527), .A(g15858) );
  INV_X1 NOT_5837( .ZN(g17439), .A(II23527) );
  INV_X1 NOT_5838( .ZN(II23530), .A(g14885) );
  INV_X1 NOT_5839( .ZN(g17442), .A(II23530) );
  INV_X1 NOT_5840( .ZN(g17445), .A(g16250) );
  INV_X1 NOT_5841( .ZN(II23539), .A(g13524) );
  INV_X1 NOT_5842( .ZN(g17451), .A(II23539) );
  INV_X1 NOT_5843( .ZN(II23542), .A(g15835) );
  INV_X1 NOT_5844( .ZN(g17454), .A(II23542) );
  INV_X1 NOT_5845( .ZN(II23545), .A(g15867) );
  INV_X1 NOT_5846( .ZN(g17457), .A(II23545) );
  INV_X1 NOT_5847( .ZN(II23553), .A(g13525) );
  INV_X1 NOT_5848( .ZN(g17465), .A(II23553) );
  INV_X1 NOT_5849( .ZN(II23556), .A(g15837) );
  INV_X1 NOT_5850( .ZN(g17468), .A(II23556) );
  INV_X1 NOT_5851( .ZN(II23559), .A(g15869) );
  INV_X1 NOT_5852( .ZN(g17471), .A(II23559) );
  INV_X1 NOT_5853( .ZN(II23564), .A(g13526) );
  INV_X1 NOT_5854( .ZN(g17476), .A(II23564) );
  INV_X1 NOT_5855( .ZN(II23567), .A(g15839) );
  INV_X1 NOT_5856( .ZN(g17479), .A(II23567) );
  INV_X1 NOT_5857( .ZN(II23570), .A(g15871) );
  INV_X1 NOT_5858( .ZN(g17482), .A(II23570) );
  INV_X1 NOT_5859( .ZN(II23575), .A(g15843) );
  INV_X1 NOT_5860( .ZN(g17487), .A(II23575) );
  INV_X1 NOT_5861( .ZN(II23578), .A(g15879) );
  INV_X1 NOT_5862( .ZN(g17490), .A(II23578) );
  INV_X1 NOT_5863( .ZN(II23581), .A(g13528) );
  INV_X1 NOT_5864( .ZN(g17493), .A(II23581) );
  INV_X1 NOT_5865( .ZN(II23584), .A(g15845) );
  INV_X1 NOT_5866( .ZN(g17496), .A(II23584) );
  INV_X1 NOT_5867( .ZN(g17499), .A(g16292) );
  INV_X1 NOT_5868( .ZN(II23588), .A(g14885) );
  INV_X1 NOT_5869( .ZN(g17500), .A(II23588) );
  INV_X1 NOT_5870( .ZN(II23591), .A(g14885) );
  INV_X1 NOT_5871( .ZN(g17503), .A(II23591) );
  INV_X1 NOT_5872( .ZN(II23599), .A(g15887) );
  INV_X1 NOT_5873( .ZN(g17511), .A(II23599) );
  INV_X1 NOT_5874( .ZN(II23602), .A(g13529) );
  INV_X1 NOT_5875( .ZN(g17514), .A(II23602) );
  INV_X1 NOT_5876( .ZN(II23605), .A(g15847) );
  INV_X1 NOT_5877( .ZN(g17517), .A(II23605) );
  INV_X1 NOT_5878( .ZN(II23608), .A(g15889) );
  INV_X1 NOT_5879( .ZN(g17520), .A(II23608) );
  INV_X1 NOT_5880( .ZN(II23611), .A(g14966) );
  INV_X1 NOT_5881( .ZN(g17523), .A(II23611) );
  INV_X1 NOT_5882( .ZN(II23619), .A(g13535) );
  INV_X1 NOT_5883( .ZN(g17531), .A(II23619) );
  INV_X1 NOT_5884( .ZN(II23622), .A(g15849) );
  INV_X1 NOT_5885( .ZN(g17534), .A(II23622) );
  INV_X1 NOT_5886( .ZN(II23625), .A(g15898) );
  INV_X1 NOT_5887( .ZN(g17537), .A(II23625) );
  INV_X1 NOT_5888( .ZN(II23633), .A(g13536) );
  INV_X1 NOT_5889( .ZN(g17545), .A(II23633) );
  INV_X2 NOT_5890( .ZN(II23636), .A(g15851) );
  INV_X2 NOT_5891( .ZN(g17548), .A(II23636) );
  INV_X1 NOT_5892( .ZN(II23639), .A(g15900) );
  INV_X1 NOT_5893( .ZN(g17551), .A(II23639) );
  INV_X1 NOT_5894( .ZN(II23645), .A(g13537) );
  INV_X1 NOT_5895( .ZN(g17557), .A(II23645) );
  INV_X1 NOT_5896( .ZN(II23648), .A(g15857) );
  INV_X1 NOT_5897( .ZN(g17560), .A(II23648) );
  INV_X1 NOT_5898( .ZN(II23651), .A(g13538) );
  INV_X1 NOT_5899( .ZN(g17563), .A(II23651) );
  INV_X1 NOT_5900( .ZN(g17566), .A(g16346) );
  INV_X1 NOT_5901( .ZN(II23655), .A(g14831) );
  INV_X1 NOT_5902( .ZN(g17567), .A(II23655) );
  INV_X1 NOT_5903( .ZN(II23658), .A(g14885) );
  INV_X1 NOT_5904( .ZN(g17570), .A(II23658) );
  INV_X1 NOT_5905( .ZN(II23661), .A(g16085) );
  INV_X1 NOT_5906( .ZN(g17573), .A(II23661) );
  INV_X1 NOT_5907( .ZN(II23667), .A(g15866) );
  INV_X1 NOT_5908( .ZN(g17579), .A(II23667) );
  INV_X1 NOT_5909( .ZN(II23670), .A(g15912) );
  INV_X1 NOT_5910( .ZN(g17582), .A(II23670) );
  INV_X1 NOT_5911( .ZN(II23673), .A(g13539) );
  INV_X1 NOT_5912( .ZN(g17585), .A(II23673) );
  INV_X1 NOT_5913( .ZN(II23676), .A(g15868) );
  INV_X1 NOT_5914( .ZN(g17588), .A(II23676) );
  INV_X1 NOT_5915( .ZN(II23679), .A(g14966) );
  INV_X1 NOT_5916( .ZN(g17591), .A(II23679) );
  INV_X1 NOT_5917( .ZN(II23682), .A(g14966) );
  INV_X1 NOT_5918( .ZN(g17594), .A(II23682) );
  INV_X1 NOT_5919( .ZN(II23689), .A(g15920) );
  INV_X1 NOT_5920( .ZN(g17601), .A(II23689) );
  INV_X1 NOT_5921( .ZN(II23692), .A(g13540) );
  INV_X1 NOT_5922( .ZN(g17604), .A(II23692) );
  INV_X1 NOT_5923( .ZN(II23695), .A(g15870) );
  INV_X1 NOT_5924( .ZN(g17607), .A(II23695) );
  INV_X1 NOT_5925( .ZN(II23698), .A(g15922) );
  INV_X1 NOT_5926( .ZN(g17610), .A(II23698) );
  INV_X1 NOT_5927( .ZN(II23701), .A(g15055) );
  INV_X1 NOT_5928( .ZN(g17613), .A(II23701) );
  INV_X1 NOT_5929( .ZN(II23709), .A(g13546) );
  INV_X1 NOT_5930( .ZN(g17621), .A(II23709) );
  INV_X1 NOT_5931( .ZN(II23712), .A(g15872) );
  INV_X1 NOT_5932( .ZN(g17624), .A(II23712) );
  INV_X1 NOT_5933( .ZN(II23715), .A(g15931) );
  INV_X1 NOT_5934( .ZN(g17627), .A(II23715) );
  INV_X1 NOT_5935( .ZN(II23725), .A(g13547) );
  INV_X1 NOT_5936( .ZN(g17637), .A(II23725) );
  INV_X1 NOT_5937( .ZN(g17640), .A(g13873) );
  INV_X1 NOT_5938( .ZN(II23729), .A(g14337) );
  INV_X1 NOT_5939( .ZN(g17645), .A(II23729) );
  INV_X1 NOT_5940( .ZN(g17648), .A(g16384) );
  INV_X1 NOT_5941( .ZN(II23733), .A(g14831) );
  INV_X1 NOT_5942( .ZN(g17649), .A(II23733) );
  INV_X1 NOT_5943( .ZN(II23739), .A(g13548) );
  INV_X1 NOT_5944( .ZN(g17655), .A(II23739) );
  INV_X1 NOT_5945( .ZN(II23742), .A(g15888) );
  INV_X1 NOT_5946( .ZN(g17658), .A(II23742) );
  INV_X1 NOT_5947( .ZN(II23745), .A(g13549) );
  INV_X2 NOT_5948( .ZN(g17661), .A(II23745) );
  INV_X2 NOT_5949( .ZN(II23748), .A(g14904) );
  INV_X1 NOT_5950( .ZN(g17664), .A(II23748) );
  INV_X1 NOT_5951( .ZN(II23751), .A(g14966) );
  INV_X1 NOT_5952( .ZN(g17667), .A(II23751) );
  INV_X1 NOT_5953( .ZN(II23754), .A(g16123) );
  INV_X1 NOT_5954( .ZN(g17670), .A(II23754) );
  INV_X1 NOT_5955( .ZN(II23760), .A(g15897) );
  INV_X1 NOT_5956( .ZN(g17676), .A(II23760) );
  INV_X1 NOT_5957( .ZN(II23763), .A(g15941) );
  INV_X1 NOT_5958( .ZN(g17679), .A(II23763) );
  INV_X1 NOT_5959( .ZN(II23766), .A(g13550) );
  INV_X1 NOT_5960( .ZN(g17682), .A(II23766) );
  INV_X1 NOT_5961( .ZN(II23769), .A(g15899) );
  INV_X1 NOT_5962( .ZN(g17685), .A(II23769) );
  INV_X1 NOT_5963( .ZN(II23772), .A(g15055) );
  INV_X1 NOT_5964( .ZN(g17688), .A(II23772) );
  INV_X1 NOT_5965( .ZN(II23775), .A(g15055) );
  INV_X1 NOT_5966( .ZN(g17691), .A(II23775) );
  INV_X1 NOT_5967( .ZN(II23782), .A(g15949) );
  INV_X1 NOT_5968( .ZN(g17698), .A(II23782) );
  INV_X1 NOT_5969( .ZN(II23785), .A(g13551) );
  INV_X1 NOT_5970( .ZN(g17701), .A(II23785) );
  INV_X1 NOT_5971( .ZN(II23788), .A(g15901) );
  INV_X1 NOT_5972( .ZN(g17704), .A(II23788) );
  INV_X1 NOT_5973( .ZN(II23791), .A(g15951) );
  INV_X1 NOT_5974( .ZN(g17707), .A(II23791) );
  INV_X1 NOT_5975( .ZN(II23794), .A(g15151) );
  INV_X1 NOT_5976( .ZN(g17710), .A(II23794) );
  INV_X1 NOT_5977( .ZN(g17720), .A(g15853) );
  INV_X1 NOT_5978( .ZN(g17724), .A(g13886) );
  INV_X1 NOT_5979( .ZN(II23817), .A(g13557) );
  INV_X1 NOT_5980( .ZN(g17738), .A(II23817) );
  INV_X1 NOT_5981( .ZN(g17741), .A(g13895) );
  INV_X1 NOT_5982( .ZN(II23821), .A(g14337) );
  INV_X1 NOT_5983( .ZN(g17746), .A(II23821) );
  INV_X1 NOT_5984( .ZN(II23824), .A(g14904) );
  INV_X1 NOT_5985( .ZN(g17749), .A(II23824) );
  INV_X1 NOT_5986( .ZN(II23830), .A(g13558) );
  INV_X1 NOT_5987( .ZN(g17755), .A(II23830) );
  INV_X1 NOT_5988( .ZN(II23833), .A(g15921) );
  INV_X1 NOT_5989( .ZN(g17758), .A(II23833) );
  INV_X1 NOT_5990( .ZN(II23836), .A(g13559) );
  INV_X1 NOT_5991( .ZN(g17761), .A(II23836) );
  INV_X1 NOT_5992( .ZN(II23839), .A(g14985) );
  INV_X1 NOT_5993( .ZN(g17764), .A(II23839) );
  INV_X1 NOT_5994( .ZN(II23842), .A(g15055) );
  INV_X1 NOT_5995( .ZN(g17767), .A(II23842) );
  INV_X1 NOT_5996( .ZN(II23845), .A(g16174) );
  INV_X1 NOT_5997( .ZN(g17770), .A(II23845) );
  INV_X1 NOT_5998( .ZN(II23851), .A(g15930) );
  INV_X1 NOT_5999( .ZN(g17776), .A(II23851) );
  INV_X1 NOT_6000( .ZN(II23854), .A(g15970) );
  INV_X1 NOT_6001( .ZN(g17779), .A(II23854) );
  INV_X1 NOT_6002( .ZN(II23857), .A(g13560) );
  INV_X1 NOT_6003( .ZN(g17782), .A(II23857) );
  INV_X1 NOT_6004( .ZN(II23860), .A(g15932) );
  INV_X1 NOT_6005( .ZN(g17785), .A(II23860) );
  INV_X1 NOT_6006( .ZN(II23863), .A(g15151) );
  INV_X1 NOT_6007( .ZN(g17788), .A(II23863) );
  INV_X1 NOT_6008( .ZN(II23866), .A(g15151) );
  INV_X1 NOT_6009( .ZN(g17791), .A(II23866) );
  INV_X1 NOT_6010( .ZN(II23874), .A(g15797) );
  INV_X1 NOT_6011( .ZN(g17799), .A(II23874) );
  INV_X1 NOT_6012( .ZN(g17802), .A(g13907) );
  INV_X1 NOT_6013( .ZN(II23888), .A(g14685) );
  INV_X1 NOT_6014( .ZN(g17815), .A(II23888) );
  INV_X1 NOT_6015( .ZN(g17825), .A(g13927) );
  INV_X1 NOT_6016( .ZN(II23904), .A(g13561) );
  INV_X1 NOT_6017( .ZN(g17839), .A(II23904) );
  INV_X1 NOT_6018( .ZN(g17842), .A(g13936) );
  INV_X1 NOT_6019( .ZN(II23908), .A(g14337) );
  INV_X1 NOT_6020( .ZN(g17847), .A(II23908) );
  INV_X1 NOT_6021( .ZN(II23911), .A(g14985) );
  INV_X1 NOT_6022( .ZN(g17850), .A(II23911) );
  INV_X1 NOT_6023( .ZN(II23917), .A(g13562) );
  INV_X1 NOT_6024( .ZN(g17856), .A(II23917) );
  INV_X1 NOT_6025( .ZN(II23920), .A(g15950) );
  INV_X1 NOT_6026( .ZN(g17859), .A(II23920) );
  INV_X1 NOT_6027( .ZN(II23923), .A(g13563) );
  INV_X1 NOT_6028( .ZN(g17862), .A(II23923) );
  INV_X1 NOT_6029( .ZN(II23926), .A(g15074) );
  INV_X1 NOT_6030( .ZN(g17865), .A(II23926) );
  INV_X1 NOT_6031( .ZN(II23929), .A(g15151) );
  INV_X1 NOT_6032( .ZN(g17868), .A(II23929) );
  INV_X1 NOT_6033( .ZN(II23932), .A(g16233) );
  INV_X1 NOT_6034( .ZN(g17871), .A(II23932) );
  INV_X1 NOT_6035( .ZN(g17878), .A(g15830) );
  INV_X1 NOT_6036( .ZN(g17882), .A(g13946) );
  INV_X1 NOT_6037( .ZN(g17892), .A(g13954) );
  INV_X1 NOT_6038( .ZN(g17893), .A(g14165) );
  INV_X1 NOT_6039( .ZN(II23954), .A(g16154) );
  INV_X1 NOT_6040( .ZN(g17903), .A(II23954) );
  INV_X1 NOT_6041( .ZN(g17914), .A(g13963) );
  INV_X1 NOT_6042( .ZN(II23976), .A(g14719) );
  INV_X1 NOT_6043( .ZN(g17927), .A(II23976) );
  INV_X1 NOT_6044( .ZN(g17937), .A(g13983) );
  INV_X1 NOT_6045( .ZN(II23992), .A(g13564) );
  INV_X1 NOT_6046( .ZN(g17951), .A(II23992) );
  INV_X1 NOT_6047( .ZN(g17954), .A(g13992) );
  INV_X1 NOT_6048( .ZN(II23996), .A(g14337) );
  INV_X1 NOT_6049( .ZN(g17959), .A(II23996) );
  INV_X1 NOT_6050( .ZN(II23999), .A(g15074) );
  INV_X1 NOT_6051( .ZN(g17962), .A(II23999) );
  INV_X1 NOT_6052( .ZN(g17969), .A(g15841) );
  INV_X1 NOT_6053( .ZN(g17974), .A(g14001) );
  INV_X1 NOT_6054( .ZN(g17984), .A(g14008) );
  INV_X1 NOT_6055( .ZN(g17988), .A(g14685) );
  INV_X2 NOT_6056( .ZN(g17991), .A(g14450) );
  INV_X2 NOT_6057( .ZN(g17993), .A(g14016) );
  INV_X1 NOT_6058( .ZN(g18003), .A(g14024) );
  INV_X1 NOT_6059( .ZN(g18004), .A(g14280) );
  INV_X1 NOT_6060( .ZN(II24049), .A(g16213) );
  INV_X1 NOT_6061( .ZN(g18014), .A(II24049) );
  INV_X1 NOT_6062( .ZN(g18025), .A(g14033) );
  INV_X1 NOT_6063( .ZN(II24071), .A(g14747) );
  INV_X1 NOT_6064( .ZN(g18038), .A(II24071) );
  INV_X1 NOT_6065( .ZN(g18048), .A(g14053) );
  INV_X1 NOT_6066( .ZN(g18063), .A(g15660) );
  INV_X1 NOT_6067( .ZN(g18070), .A(g15854) );
  INV_X1 NOT_6068( .ZN(g18074), .A(g14062) );
  INV_X1 NOT_6069( .ZN(g18084), .A(g14068) );
  INV_X1 NOT_6070( .ZN(g18089), .A(g14355) );
  INV_X1 NOT_6071( .ZN(g18091), .A(g14092) );
  INV_X1 NOT_6072( .ZN(g18101), .A(g14099) );
  INV_X1 NOT_6073( .ZN(g18105), .A(g14719) );
  INV_X1 NOT_6074( .ZN(g18108), .A(g14537) );
  INV_X1 NOT_6075( .ZN(g18110), .A(g14107) );
  INV_X1 NOT_6076( .ZN(g18120), .A(g14115) );
  INV_X1 NOT_6077( .ZN(g18121), .A(g14402) );
  INV_X1 NOT_6078( .ZN(II24144), .A(g16278) );
  INV_X1 NOT_6079( .ZN(g18131), .A(II24144) );
  INV_X1 NOT_6080( .ZN(g18142), .A(g14124) );
  INV_X1 NOT_6081( .ZN(II24166), .A(g14768) );
  INV_X1 NOT_6082( .ZN(g18155), .A(II24166) );
  INV_X1 NOT_6083( .ZN(II24171), .A(g16439) );
  INV_X1 NOT_6084( .ZN(g18166), .A(II24171) );
  INV_X1 NOT_6085( .ZN(g18170), .A(g15877) );
  INV_X1 NOT_6086( .ZN(g18174), .A(g14148) );
  INV_X1 NOT_6087( .ZN(g18179), .A(g14153) );
  INV_X1 NOT_6088( .ZN(g18188), .A(g14252) );
  INV_X1 NOT_6089( .ZN(g18190), .A(g14177) );
  INV_X1 NOT_6090( .ZN(g18200), .A(g14183) );
  INV_X1 NOT_6091( .ZN(g18205), .A(g14467) );
  INV_X1 NOT_6092( .ZN(g18207), .A(g14207) );
  INV_X1 NOT_6093( .ZN(g18217), .A(g14214) );
  INV_X1 NOT_6094( .ZN(g18221), .A(g14747) );
  INV_X1 NOT_6095( .ZN(g18224), .A(g14592) );
  INV_X1 NOT_6096( .ZN(g18226), .A(g14222) );
  INV_X1 NOT_6097( .ZN(g18236), .A(g14230) );
  INV_X1 NOT_6098( .ZN(g18237), .A(g14514) );
  INV_X1 NOT_6099( .ZN(II24247), .A(g16337) );
  INV_X1 NOT_6100( .ZN(g18247), .A(II24247) );
  INV_X1 NOT_6101( .ZN(II24258), .A(g16463) );
  INV_X1 NOT_6102( .ZN(g18258), .A(II24258) );
  INV_X1 NOT_6103( .ZN(g18261), .A(g15719) );
  INV_X1 NOT_6104( .ZN(g18265), .A(g14238) );
  INV_X1 NOT_6105( .ZN(g18275), .A(g14171) );
  INV_X1 NOT_6106( .ZN(II24285), .A(g15992) );
  INV_X1 NOT_6107( .ZN(g18278), .A(II24285) );
  INV_X1 NOT_6108( .ZN(g18281), .A(g14263) );
  INV_X1 NOT_6109( .ZN(g18286), .A(g14268) );
  INV_X1 NOT_6110( .ZN(g18295), .A(g14374) );
  INV_X1 NOT_6111( .ZN(g18297), .A(g14292) );
  INV_X1 NOT_6112( .ZN(g18307), .A(g14298) );
  INV_X1 NOT_6113( .ZN(g18312), .A(g14554) );
  INV_X1 NOT_6114( .ZN(g18314), .A(g14322) );
  INV_X1 NOT_6115( .ZN(g18324), .A(g14329) );
  INV_X1 NOT_6116( .ZN(g18328), .A(g14768) );
  INV_X1 NOT_6117( .ZN(g18331), .A(g14626) );
  INV_X1 NOT_6118( .ZN(II24346), .A(g15873) );
  INV_X1 NOT_6119( .ZN(g18334), .A(II24346) );
  INV_X1 NOT_6120( .ZN(g18337), .A(g15757) );
  INV_X1 NOT_6121( .ZN(g18341), .A(g14342) );
  INV_X1 NOT_6122( .ZN(g18351), .A(g13741) );
  INV_X1 NOT_6123( .ZN(g18353), .A(g13918) );
  INV_X1 NOT_6124( .ZN(II24368), .A(g15990) );
  INV_X1 NOT_6125( .ZN(g18355), .A(II24368) );
  INV_X1 NOT_6126( .ZN(g18358), .A(g14360) );
  INV_X1 NOT_6127( .ZN(g18368), .A(g14286) );
  INV_X1 NOT_6128( .ZN(II24394), .A(g15995) );
  INV_X1 NOT_6129( .ZN(g18371), .A(II24394) );
  INV_X1 NOT_6130( .ZN(g18374), .A(g14385) );
  INV_X1 NOT_6131( .ZN(g18379), .A(g14390) );
  INV_X1 NOT_6132( .ZN(g18388), .A(g14486) );
  INV_X1 NOT_6133( .ZN(g18390), .A(g14414) );
  INV_X1 NOT_6134( .ZN(g18400), .A(g14420) );
  INV_X1 NOT_6135( .ZN(g18405), .A(g14609) );
  INV_X1 NOT_6136( .ZN(g18407), .A(g15959) );
  INV_X1 NOT_6137( .ZN(g18414), .A(g15718) );
  INV_X1 NOT_6138( .ZN(g18415), .A(g15783) );
  INV_X1 NOT_6139( .ZN(g18429), .A(g14831) );
  INV_X1 NOT_6140( .ZN(II24459), .A(g13599) );
  INV_X1 NOT_6141( .ZN(g18432), .A(II24459) );
  INV_X1 NOT_6142( .ZN(g18435), .A(g14359) );
  INV_X1 NOT_6143( .ZN(g18436), .A(g14454) );
  INV_X1 NOT_6144( .ZN(g18446), .A(g13741) );
  INV_X1 NOT_6145( .ZN(g18448), .A(g13974) );
  INV_X1 NOT_6146( .ZN(II24481), .A(g15993) );
  INV_X1 NOT_6147( .ZN(g18450), .A(II24481) );
  INV_X1 NOT_6148( .ZN(g18453), .A(g14472) );
  INV_X1 NOT_6149( .ZN(g18463), .A(g14408) );
  INV_X1 NOT_6150( .ZN(II24507), .A(g15999) );
  INV_X1 NOT_6151( .ZN(g18466), .A(II24507) );
  INV_X1 NOT_6152( .ZN(g18469), .A(g14497) );
  INV_X1 NOT_6153( .ZN(g18474), .A(g14502) );
  INV_X1 NOT_6154( .ZN(g18483), .A(g14573) );
  INV_X1 NOT_6155( .ZN(g18485), .A(g15756) );
  INV_X1 NOT_6156( .ZN(g18486), .A(g15804) );
  INV_X1 NOT_6157( .ZN(g18490), .A(g13565) );
  INV_X1 NOT_6158( .ZN(g18502), .A(g14904) );
  INV_X1 NOT_6159( .ZN(II24560), .A(g13611) );
  INV_X1 NOT_6160( .ZN(g18505), .A(II24560) );
  INV_X2 NOT_6161( .ZN(g18508), .A(g14471) );
  INV_X2 NOT_6162( .ZN(g18509), .A(g14541) );
  INV_X1 NOT_6163( .ZN(g18519), .A(g13741) );
  INV_X1 NOT_6164( .ZN(g18521), .A(g14044) );
  INV_X1 NOT_6165( .ZN(II24582), .A(g15996) );
  INV_X1 NOT_6166( .ZN(g18523), .A(II24582) );
  INV_X1 NOT_6167( .ZN(g18526), .A(g14559) );
  INV_X1 NOT_6168( .ZN(g18536), .A(g14520) );
  INV_X1 NOT_6169( .ZN(II24608), .A(g16006) );
  INV_X1 NOT_6170( .ZN(g18539), .A(II24608) );
  INV_X1 NOT_6171( .ZN(g18543), .A(g15819) );
  INV_X1 NOT_6172( .ZN(g18552), .A(g16154) );
  INV_X1 NOT_6173( .ZN(g18554), .A(g13573) );
  INV_X1 NOT_6174( .ZN(g18566), .A(g14985) );
  INV_X1 NOT_6175( .ZN(II24662), .A(g13621) );
  INV_X1 NOT_6176( .ZN(g18569), .A(II24662) );
  INV_X1 NOT_6177( .ZN(g18572), .A(g14558) );
  INV_X1 NOT_6178( .ZN(g18573), .A(g14596) );
  INV_X1 NOT_6179( .ZN(g18583), .A(g13741) );
  INV_X1 NOT_6180( .ZN(g18585), .A(g14135) );
  INV_X1 NOT_6181( .ZN(II24684), .A(g16000) );
  INV_X1 NOT_6182( .ZN(g18587), .A(II24684) );
  INV_X1 NOT_6183( .ZN(g18593), .A(g15831) );
  INV_X1 NOT_6184( .ZN(g18602), .A(g16213) );
  INV_X1 NOT_6185( .ZN(g18604), .A(g13582) );
  INV_X1 NOT_6186( .ZN(g18616), .A(g15074) );
  INV_X1 NOT_6187( .ZN(II24732), .A(g13633) );
  INV_X1 NOT_6188( .ZN(g18619), .A(II24732) );
  INV_X1 NOT_6189( .ZN(g18622), .A(g14613) );
  INV_X1 NOT_6190( .ZN(g18634), .A(g16278) );
  INV_X1 NOT_6191( .ZN(g18636), .A(g13602) );
  INV_X1 NOT_6192( .ZN(g18643), .A(g16337) );
  INV_X1 NOT_6193( .ZN(g18646), .A(g16341) );
  INV_X1 NOT_6194( .ZN(g18656), .A(g14776) );
  INV_X1 NOT_6195( .ZN(g18670), .A(g14797) );
  INV_X1 NOT_6196( .ZN(g18679), .A(g14811) );
  INV_X1 NOT_6197( .ZN(g18691), .A(g14885) );
  INV_X1 NOT_6198( .ZN(g18692), .A(g14837) );
  INV_X1 NOT_6199( .ZN(g18699), .A(g14849) );
  INV_X1 NOT_6200( .ZN(g18708), .A(g14863) );
  INV_X1 NOT_6201( .ZN(g18720), .A(g14895) );
  INV_X1 NOT_6202( .ZN(g18725), .A(g13865) );
  INV_X1 NOT_6203( .ZN(g18727), .A(g14966) );
  INV_X1 NOT_6204( .ZN(g18728), .A(g14910) );
  INV_X1 NOT_6205( .ZN(g18735), .A(g14922) );
  INV_X1 NOT_6206( .ZN(g18744), .A(g14936) );
  INV_X1 NOT_6207( .ZN(g18756), .A(g14960) );
  INV_X1 NOT_6208( .ZN(g18757), .A(g14963) );
  INV_X1 NOT_6209( .ZN(g18758), .A(g14976) );
  INV_X1 NOT_6210( .ZN(g18764), .A(g15055) );
  INV_X1 NOT_6211( .ZN(g18765), .A(g14991) );
  INV_X1 NOT_6212( .ZN(g18772), .A(g15003) );
  INV_X1 NOT_6213( .ZN(g18783), .A(g15034) );
  INV_X1 NOT_6214( .ZN(g18784), .A(g15037) );
  INV_X1 NOT_6215( .ZN(g18785), .A(g15040) );
  INV_X1 NOT_6216( .ZN(g18786), .A(g15043) );
  INV_X1 NOT_6217( .ZN(g18787), .A(g15049) );
  INV_X1 NOT_6218( .ZN(g18788), .A(g15052) );
  INV_X1 NOT_6219( .ZN(g18789), .A(g15065) );
  INV_X1 NOT_6220( .ZN(g18795), .A(g15151) );
  INV_X1 NOT_6221( .ZN(g18796), .A(g15080) );
  INV_X1 NOT_6222( .ZN(g18805), .A(g15106) );
  INV_X1 NOT_6223( .ZN(g18806), .A(g15109) );
  INV_X1 NOT_6224( .ZN(g18807), .A(g15112) );
  INV_X1 NOT_6225( .ZN(g18808), .A(g15115) );
  INV_X1 NOT_6226( .ZN(g18809), .A(g15130) );
  INV_X1 NOT_6227( .ZN(g18810), .A(g15133) );
  INV_X1 NOT_6228( .ZN(g18811), .A(g15136) );
  INV_X1 NOT_6229( .ZN(g18812), .A(g15139) );
  INV_X1 NOT_6230( .ZN(g18813), .A(g15145) );
  INV_X1 NOT_6231( .ZN(g18814), .A(g15148) );
  INV_X1 NOT_6232( .ZN(g18815), .A(g15161) );
  INV_X1 NOT_6233( .ZN(g18822), .A(g15179) );
  INV_X1 NOT_6234( .ZN(g18823), .A(g15182) );
  INV_X1 NOT_6235( .ZN(g18824), .A(g15185) );
  INV_X1 NOT_6236( .ZN(g18825), .A(g15198) );
  INV_X1 NOT_6237( .ZN(g18826), .A(g15201) );
  INV_X1 NOT_6238( .ZN(g18827), .A(g15204) );
  INV_X1 NOT_6239( .ZN(g18828), .A(g15207) );
  INV_X1 NOT_6240( .ZN(g18829), .A(g15222) );
  INV_X1 NOT_6241( .ZN(g18830), .A(g15225) );
  INV_X1 NOT_6242( .ZN(g18831), .A(g15228) );
  INV_X1 NOT_6243( .ZN(g18832), .A(g15231) );
  INV_X1 NOT_6244( .ZN(g18833), .A(g15237) );
  INV_X1 NOT_6245( .ZN(g18834), .A(g15240) );
  INV_X1 NOT_6246( .ZN(g18838), .A(g15248) );
  INV_X1 NOT_6247( .ZN(g18839), .A(g15251) );
  INV_X1 NOT_6248( .ZN(g18840), .A(g15254) );
  INV_X1 NOT_6249( .ZN(g18841), .A(g15265) );
  INV_X1 NOT_6250( .ZN(g18842), .A(g15268) );
  INV_X1 NOT_6251( .ZN(g18843), .A(g15271) );
  INV_X1 NOT_6252( .ZN(g18844), .A(g15284) );
  INV_X1 NOT_6253( .ZN(g18845), .A(g15287) );
  INV_X1 NOT_6254( .ZN(g18846), .A(g15290) );
  INV_X1 NOT_6255( .ZN(g18847), .A(g15293) );
  INV_X1 NOT_6256( .ZN(g18848), .A(g15308) );
  INV_X1 NOT_6257( .ZN(g18849), .A(g15311) );
  INV_X1 NOT_6258( .ZN(g18850), .A(g15314) );
  INV_X1 NOT_6259( .ZN(g18851), .A(g15317) );
  INV_X1 NOT_6260( .ZN(g18853), .A(g15326) );
  INV_X1 NOT_6261( .ZN(g18854), .A(g15329) );
  INV_X1 NOT_6262( .ZN(g18855), .A(g15332) );
  INV_X1 NOT_6263( .ZN(g18856), .A(g15340) );
  INV_X1 NOT_6264( .ZN(g18857), .A(g15343) );
  INV_X1 NOT_6265( .ZN(g18858), .A(g15346) );
  INV_X1 NOT_6266( .ZN(g18859), .A(g15357) );
  INV_X1 NOT_6267( .ZN(g18860), .A(g15360) );
  INV_X1 NOT_6268( .ZN(g18861), .A(g15363) );
  INV_X1 NOT_6269( .ZN(g18862), .A(g15376) );
  INV_X1 NOT_6270( .ZN(g18863), .A(g15379) );
  INV_X1 NOT_6271( .ZN(g18864), .A(g15382) );
  INV_X1 NOT_6272( .ZN(g18865), .A(g15385) );
  INV_X1 NOT_6273( .ZN(II24894), .A(g14797) );
  INV_X1 NOT_6274( .ZN(g18869), .A(II24894) );
  INV_X1 NOT_6275( .ZN(g18870), .A(g15393) );
  INV_X1 NOT_6276( .ZN(g18871), .A(g15396) );
  INV_X1 NOT_6277( .ZN(g18872), .A(g15399) );
  INV_X1 NOT_6278( .ZN(g18873), .A(g15404) );
  INV_X1 NOT_6279( .ZN(g18874), .A(g15412) );
  INV_X1 NOT_6280( .ZN(g18875), .A(g15415) );
  INV_X1 NOT_6281( .ZN(g18876), .A(g15418) );
  INV_X1 NOT_6282( .ZN(g18877), .A(g15426) );
  INV_X1 NOT_6283( .ZN(g18878), .A(g15429) );
  INV_X1 NOT_6284( .ZN(g18879), .A(g15432) );
  INV_X1 NOT_6285( .ZN(g18880), .A(g15443) );
  INV_X1 NOT_6286( .ZN(g18881), .A(g15446) );
  INV_X1 NOT_6287( .ZN(g18882), .A(g15449) );
  INV_X1 NOT_6288( .ZN(g18884), .A(g13469) );
  INV_X1 NOT_6289( .ZN(II24913), .A(g15800) );
  INV_X1 NOT_6290( .ZN(g18886), .A(II24913) );
  INV_X1 NOT_6291( .ZN(II24916), .A(g14776) );
  INV_X1 NOT_6292( .ZN(g18890), .A(II24916) );
  INV_X1 NOT_6293( .ZN(g18891), .A(g15461) );
  INV_X1 NOT_6294( .ZN(g18892), .A(g15464) );
  INV_X1 NOT_6295( .ZN(g18893), .A(g15467) );
  INV_X1 NOT_6296( .ZN(g18894), .A(g15471) );
  INV_X1 NOT_6297( .ZN(II24923), .A(g14849) );
  INV_X1 NOT_6298( .ZN(g18895), .A(II24923) );
  INV_X1 NOT_6299( .ZN(g18896), .A(g15477) );
  INV_X1 NOT_6300( .ZN(g18897), .A(g15480) );
  INV_X1 NOT_6301( .ZN(g18898), .A(g15483) );
  INV_X1 NOT_6302( .ZN(g18899), .A(g15488) );
  INV_X1 NOT_6303( .ZN(g18900), .A(g15496) );
  INV_X1 NOT_6304( .ZN(g18901), .A(g15499) );
  INV_X1 NOT_6305( .ZN(g18902), .A(g15502) );
  INV_X1 NOT_6306( .ZN(g18903), .A(g15510) );
  INV_X1 NOT_6307( .ZN(g18904), .A(g15513) );
  INV_X1 NOT_6308( .ZN(g18905), .A(g15516) );
  INV_X1 NOT_6309( .ZN(g18908), .A(g15521) );
  INV_X1 NOT_6310( .ZN(g18909), .A(g15528) );
  INV_X1 NOT_6311( .ZN(g18910), .A(g15531) );
  INV_X1 NOT_6312( .ZN(g18911), .A(g15534) );
  INV_X1 NOT_6313( .ZN(g18912), .A(g15537) );
  INV_X1 NOT_6314( .ZN(II24943), .A(g14811) );
  INV_X1 NOT_6315( .ZN(g18913), .A(II24943) );
  INV_X1 NOT_6316( .ZN(g18914), .A(g15547) );
  INV_X1 NOT_6317( .ZN(g18915), .A(g15550) );
  INV_X1 NOT_6318( .ZN(g18916), .A(g15553) );
  INV_X1 NOT_6319( .ZN(g18917), .A(g15557) );
  INV_X1 NOT_6320( .ZN(II24950), .A(g14922) );
  INV_X1 NOT_6321( .ZN(g18918), .A(II24950) );
  INV_X1 NOT_6322( .ZN(g18919), .A(g15563) );
  INV_X1 NOT_6323( .ZN(g18920), .A(g15566) );
  INV_X1 NOT_6324( .ZN(g18921), .A(g15569) );
  INV_X1 NOT_6325( .ZN(g18922), .A(g15574) );
  INV_X1 NOT_6326( .ZN(g18923), .A(g15582) );
  INV_X1 NOT_6327( .ZN(g18924), .A(g15585) );
  INV_X1 NOT_6328( .ZN(g18925), .A(g15588) );
  INV_X1 NOT_6329( .ZN(g18926), .A(g15596) );
  INV_X1 NOT_6330( .ZN(g18927), .A(g15599) );
  INV_X1 NOT_6331( .ZN(g18928), .A(g15606) );
  INV_X1 NOT_6332( .ZN(g18929), .A(g15609) );
  INV_X1 NOT_6333( .ZN(g18930), .A(g15612) );
  INV_X1 NOT_6334( .ZN(g18931), .A(g15615) );
  INV_X1 NOT_6335( .ZN(II24966), .A(g14863) );
  INV_X1 NOT_6336( .ZN(g18932), .A(II24966) );
  INV_X4 NOT_6337( .ZN(g18933), .A(g15625) );
  INV_X4 NOT_6338( .ZN(g18934), .A(g15628) );
  INV_X1 NOT_6339( .ZN(g18935), .A(g15631) );
  INV_X1 NOT_6340( .ZN(g18936), .A(g15635) );
  INV_X1 NOT_6341( .ZN(II24973), .A(g15003) );
  INV_X1 NOT_6342( .ZN(g18937), .A(II24973) );
  INV_X1 NOT_6343( .ZN(g18938), .A(g15641) );
  INV_X1 NOT_6344( .ZN(g18939), .A(g15644) );
  INV_X1 NOT_6345( .ZN(g18940), .A(g15647) );
  INV_X1 NOT_6346( .ZN(g18941), .A(g15652) );
  INV_X1 NOT_6347( .ZN(g18943), .A(g15655) );
  INV_X1 NOT_6348( .ZN(II24982), .A(g14347) );
  INV_X1 NOT_6349( .ZN(g18944), .A(II24982) );
  INV_X1 NOT_6350( .ZN(g18945), .A(g15667) );
  INV_X1 NOT_6351( .ZN(g18946), .A(g15672) );
  INV_X1 NOT_6352( .ZN(g18947), .A(g15675) );
  INV_X1 NOT_6353( .ZN(g18948), .A(g15682) );
  INV_X1 NOT_6354( .ZN(g18949), .A(g15685) );
  INV_X1 NOT_6355( .ZN(g18950), .A(g15688) );
  INV_X1 NOT_6356( .ZN(g18951), .A(g15691) );
  INV_X1 NOT_6357( .ZN(II24992), .A(g14936) );
  INV_X1 NOT_6358( .ZN(g18952), .A(II24992) );
  INV_X1 NOT_6359( .ZN(g18953), .A(g15701) );
  INV_X1 NOT_6360( .ZN(g18954), .A(g15704) );
  INV_X1 NOT_6361( .ZN(g18955), .A(g15707) );
  INV_X1 NOT_6362( .ZN(g18956), .A(g15711) );
  INV_X1 NOT_6363( .ZN(g18958), .A(g15714) );
  INV_X1 NOT_6364( .ZN(II25001), .A(g14244) );
  INV_X1 NOT_6365( .ZN(g18959), .A(II25001) );
  INV_X1 NOT_6366( .ZN(II25004), .A(g14459) );
  INV_X1 NOT_6367( .ZN(g18960), .A(II25004) );
  INV_X1 NOT_6368( .ZN(g18961), .A(g15726) );
  INV_X1 NOT_6369( .ZN(g18962), .A(g15731) );
  INV_X1 NOT_6370( .ZN(g18963), .A(g15734) );
  INV_X1 NOT_6371( .ZN(g18964), .A(g15741) );
  INV_X1 NOT_6372( .ZN(g18965), .A(g15744) );
  INV_X1 NOT_6373( .ZN(g18966), .A(g15747) );
  INV_X1 NOT_6374( .ZN(g18967), .A(g15750) );
  INV_X1 NOT_6375( .ZN(II25015), .A(g14158) );
  INV_X1 NOT_6376( .ZN(g18969), .A(II25015) );
  INV_X1 NOT_6377( .ZN(II25018), .A(g14366) );
  INV_X1 NOT_6378( .ZN(g18970), .A(II25018) );
  INV_X1 NOT_6379( .ZN(II25021), .A(g14546) );
  INV_X1 NOT_6380( .ZN(g18971), .A(II25021) );
  INV_X1 NOT_6381( .ZN(g18972), .A(g15766) );
  INV_X1 NOT_6382( .ZN(g18973), .A(g15771) );
  INV_X1 NOT_6383( .ZN(g18974), .A(g15774) );
  INV_X1 NOT_6384( .ZN(g18976), .A(g15777) );
  INV_X1 NOT_6385( .ZN(II25037), .A(g14071) );
  INV_X1 NOT_6386( .ZN(g18981), .A(II25037) );
  INV_X1 NOT_6387( .ZN(II25041), .A(g14895) );
  INV_X1 NOT_6388( .ZN(g18983), .A(II25041) );
  INV_X1 NOT_6389( .ZN(II25044), .A(g14273) );
  INV_X1 NOT_6390( .ZN(g18984), .A(II25044) );
  INV_X1 NOT_6391( .ZN(II25047), .A(g14478) );
  INV_X1 NOT_6392( .ZN(g18985), .A(II25047) );
  INV_X1 NOT_6393( .ZN(II25050), .A(g14601) );
  INV_X1 NOT_6394( .ZN(g18986), .A(II25050) );
  INV_X1 NOT_6395( .ZN(g18987), .A(g15794) );
  INV_X1 NOT_6396( .ZN(II25054), .A(g14837) );
  INV_X1 NOT_6397( .ZN(g18988), .A(II25054) );
  INV_X1 NOT_6398( .ZN(II25057), .A(g14186) );
  INV_X1 NOT_6399( .ZN(g18989), .A(II25057) );
  INV_X1 NOT_6400( .ZN(II25061), .A(g14976) );
  INV_X1 NOT_6401( .ZN(g18991), .A(II25061) );
  INV_X1 NOT_6402( .ZN(II25064), .A(g14395) );
  INV_X1 NOT_6403( .ZN(g18992), .A(II25064) );
  INV_X1 NOT_6404( .ZN(II25067), .A(g14565) );
  INV_X1 NOT_6405( .ZN(g18993), .A(II25067) );
  INV_X1 NOT_6406( .ZN(II25071), .A(g14910) );
  INV_X1 NOT_6407( .ZN(g18995), .A(II25071) );
  INV_X1 NOT_6408( .ZN(II25074), .A(g14301) );
  INV_X1 NOT_6409( .ZN(g18996), .A(II25074) );
  INV_X1 NOT_6410( .ZN(II25078), .A(g15065) );
  INV_X1 NOT_6411( .ZN(g18998), .A(II25078) );
  INV_X1 NOT_6412( .ZN(II25081), .A(g14507) );
  INV_X1 NOT_6413( .ZN(g18999), .A(II25081) );
  INV_X1 NOT_6414( .ZN(II25084), .A(g14885) );
  INV_X1 NOT_6415( .ZN(g19000), .A(II25084) );
  INV_X1 NOT_6416( .ZN(g19001), .A(g14071) );
  INV_X1 NOT_6417( .ZN(II25089), .A(g14991) );
  INV_X4 NOT_6418( .ZN(g19008), .A(II25089) );
  INV_X4 NOT_6419( .ZN(II25092), .A(g14423) );
  INV_X1 NOT_6420( .ZN(g19009), .A(II25092) );
  INV_X1 NOT_6421( .ZN(II25096), .A(g15161) );
  INV_X1 NOT_6422( .ZN(g19011), .A(II25096) );
  INV_X1 NOT_6423( .ZN(II25099), .A(g19000) );
  INV_X1 NOT_6424( .ZN(g19012), .A(II25099) );
  INV_X1 NOT_6425( .ZN(II25102), .A(g18944) );
  INV_X1 NOT_6426( .ZN(g19013), .A(II25102) );
  INV_X1 NOT_6427( .ZN(II25105), .A(g18959) );
  INV_X1 NOT_6428( .ZN(g19014), .A(II25105) );
  INV_X1 NOT_6429( .ZN(II25108), .A(g18969) );
  INV_X1 NOT_6430( .ZN(g19015), .A(II25108) );
  INV_X1 NOT_6431( .ZN(II25111), .A(g18981) );
  INV_X1 NOT_6432( .ZN(g19016), .A(II25111) );
  INV_X1 NOT_6433( .ZN(II25114), .A(g18983) );
  INV_X1 NOT_6434( .ZN(g19017), .A(II25114) );
  INV_X1 NOT_6435( .ZN(II25117), .A(g18988) );
  INV_X1 NOT_6436( .ZN(g19018), .A(II25117) );
  INV_X1 NOT_6437( .ZN(II25120), .A(g18869) );
  INV_X1 NOT_6438( .ZN(g19019), .A(II25120) );
  INV_X1 NOT_6439( .ZN(II25123), .A(g18890) );
  INV_X1 NOT_6440( .ZN(g19020), .A(II25123) );
  INV_X1 NOT_6441( .ZN(II25126), .A(g16858) );
  INV_X1 NOT_6442( .ZN(g19021), .A(II25126) );
  INV_X1 NOT_6443( .ZN(II25129), .A(g16813) );
  INV_X1 NOT_6444( .ZN(g19022), .A(II25129) );
  INV_X1 NOT_6445( .ZN(II25132), .A(g16862) );
  INV_X1 NOT_6446( .ZN(g19023), .A(II25132) );
  INV_X1 NOT_6447( .ZN(II25135), .A(g16506) );
  INV_X1 NOT_6448( .ZN(g19024), .A(II25135) );
  INV_X1 NOT_6449( .ZN(II25138), .A(g18960) );
  INV_X1 NOT_6450( .ZN(g19025), .A(II25138) );
  INV_X1 NOT_6451( .ZN(II25141), .A(g18970) );
  INV_X1 NOT_6452( .ZN(g19026), .A(II25141) );
  INV_X1 NOT_6453( .ZN(II25144), .A(g18984) );
  INV_X1 NOT_6454( .ZN(g19027), .A(II25144) );
  INV_X1 NOT_6455( .ZN(II25147), .A(g18989) );
  INV_X1 NOT_6456( .ZN(g19028), .A(II25147) );
  INV_X1 NOT_6457( .ZN(II25150), .A(g18991) );
  INV_X1 NOT_6458( .ZN(g19029), .A(II25150) );
  INV_X1 NOT_6459( .ZN(II25153), .A(g18995) );
  INV_X1 NOT_6460( .ZN(g19030), .A(II25153) );
  INV_X1 NOT_6461( .ZN(II25156), .A(g18895) );
  INV_X1 NOT_6462( .ZN(g19031), .A(II25156) );
  INV_X1 NOT_6463( .ZN(II25159), .A(g18913) );
  INV_X1 NOT_6464( .ZN(g19032), .A(II25159) );
  INV_X1 NOT_6465( .ZN(II25162), .A(g16863) );
  INV_X1 NOT_6466( .ZN(g19033), .A(II25162) );
  INV_X1 NOT_6467( .ZN(II25165), .A(g16831) );
  INV_X1 NOT_6468( .ZN(g19034), .A(II25165) );
  INV_X1 NOT_6469( .ZN(II25168), .A(g16877) );
  INV_X1 NOT_6470( .ZN(g19035), .A(II25168) );
  INV_X1 NOT_6471( .ZN(II25171), .A(g16528) );
  INV_X1 NOT_6472( .ZN(g19036), .A(II25171) );
  INV_X1 NOT_6473( .ZN(II25174), .A(g18971) );
  INV_X1 NOT_6474( .ZN(g19037), .A(II25174) );
  INV_X1 NOT_6475( .ZN(II25177), .A(g18985) );
  INV_X1 NOT_6476( .ZN(g19038), .A(II25177) );
  INV_X1 NOT_6477( .ZN(II25180), .A(g18992) );
  INV_X1 NOT_6478( .ZN(g19039), .A(II25180) );
  INV_X1 NOT_6479( .ZN(II25183), .A(g18996) );
  INV_X1 NOT_6480( .ZN(g19040), .A(II25183) );
  INV_X1 NOT_6481( .ZN(II25186), .A(g18998) );
  INV_X1 NOT_6482( .ZN(g19041), .A(II25186) );
  INV_X1 NOT_6483( .ZN(II25189), .A(g19008) );
  INV_X1 NOT_6484( .ZN(g19042), .A(II25189) );
  INV_X1 NOT_6485( .ZN(II25192), .A(g18918) );
  INV_X1 NOT_6486( .ZN(g19043), .A(II25192) );
  INV_X1 NOT_6487( .ZN(II25195), .A(g18932) );
  INV_X1 NOT_6488( .ZN(g19044), .A(II25195) );
  INV_X1 NOT_6489( .ZN(II25198), .A(g16878) );
  INV_X1 NOT_6490( .ZN(g19045), .A(II25198) );
  INV_X1 NOT_6491( .ZN(II25201), .A(g16843) );
  INV_X1 NOT_6492( .ZN(g19046), .A(II25201) );
  INV_X1 NOT_6493( .ZN(II25204), .A(g16905) );
  INV_X1 NOT_6494( .ZN(g19047), .A(II25204) );
  INV_X1 NOT_6495( .ZN(II25207), .A(g16559) );
  INV_X1 NOT_6496( .ZN(g19048), .A(II25207) );
  INV_X1 NOT_6497( .ZN(II25210), .A(g18986) );
  INV_X2 NOT_6498( .ZN(g19049), .A(II25210) );
  INV_X2 NOT_6499( .ZN(II25213), .A(g18993) );
  INV_X1 NOT_6500( .ZN(g19050), .A(II25213) );
  INV_X1 NOT_6501( .ZN(II25216), .A(g18999) );
  INV_X1 NOT_6502( .ZN(g19051), .A(II25216) );
  INV_X1 NOT_6503( .ZN(II25219), .A(g19009) );
  INV_X1 NOT_6504( .ZN(g19052), .A(II25219) );
  INV_X1 NOT_6505( .ZN(II25222), .A(g19011) );
  INV_X1 NOT_6506( .ZN(g19053), .A(II25222) );
  INV_X1 NOT_6507( .ZN(II25225), .A(g16514) );
  INV_X1 NOT_6508( .ZN(g19054), .A(II25225) );
  INV_X1 NOT_6509( .ZN(II25228), .A(g18937) );
  INV_X1 NOT_6510( .ZN(g19055), .A(II25228) );
  INV_X1 NOT_6511( .ZN(II25231), .A(g18952) );
  INV_X1 NOT_6512( .ZN(g19056), .A(II25231) );
  INV_X1 NOT_6513( .ZN(II25234), .A(g16906) );
  INV_X1 NOT_6514( .ZN(g19057), .A(II25234) );
  INV_X1 NOT_6515( .ZN(II25237), .A(g16849) );
  INV_X1 NOT_6516( .ZN(g19058), .A(II25237) );
  INV_X1 NOT_6517( .ZN(II25240), .A(g16934) );
  INV_X1 NOT_6518( .ZN(g19059), .A(II25240) );
  INV_X1 NOT_6519( .ZN(II25243), .A(g17227) );
  INV_X1 NOT_6520( .ZN(g19060), .A(II25243) );
  INV_X1 NOT_6521( .ZN(II25246), .A(g17233) );
  INV_X1 NOT_6522( .ZN(g19061), .A(II25246) );
  INV_X1 NOT_6523( .ZN(II25249), .A(g17300) );
  INV_X1 NOT_6524( .ZN(g19062), .A(II25249) );
  INV_X1 NOT_6525( .ZN(II25253), .A(g17124) );
  INV_X1 NOT_6526( .ZN(g19064), .A(II25253) );
  INV_X1 NOT_6527( .ZN(g19070), .A(g18583) );
  INV_X1 NOT_6528( .ZN(II25258), .A(g16974) );
  INV_X1 NOT_6529( .ZN(g19075), .A(II25258) );
  INV_X1 NOT_6530( .ZN(g19078), .A(g18619) );
  INV_X1 NOT_6531( .ZN(II25264), .A(g17151) );
  INV_X1 NOT_6532( .ZN(g19081), .A(II25264) );
  INV_X1 NOT_6533( .ZN(II25272), .A(g17051) );
  INV_X1 NOT_6534( .ZN(g19091), .A(II25272) );
  INV_X1 NOT_6535( .ZN(g19096), .A(g18980) );
  INV_X1 NOT_6536( .ZN(II25283), .A(g17086) );
  INV_X1 NOT_6537( .ZN(g19098), .A(II25283) );
  INV_X1 NOT_6538( .ZN(II25294), .A(g17124) );
  INV_X1 NOT_6539( .ZN(g19105), .A(II25294) );
  INV_X1 NOT_6540( .ZN(II25303), .A(g17151) );
  INV_X1 NOT_6541( .ZN(g19110), .A(II25303) );
  INV_X1 NOT_6542( .ZN(II25308), .A(g16867) );
  INV_X1 NOT_6543( .ZN(g19113), .A(II25308) );
  INV_X1 NOT_6544( .ZN(II25315), .A(g16895) );
  INV_X1 NOT_6545( .ZN(g19118), .A(II25315) );
  INV_X1 NOT_6546( .ZN(II25320), .A(g16924) );
  INV_X1 NOT_6547( .ZN(g19125), .A(II25320) );
  INV_X1 NOT_6548( .ZN(II25325), .A(g16954) );
  INV_X1 NOT_6549( .ZN(g19132), .A(II25325) );
  INV_X1 NOT_6550( .ZN(II25334), .A(g17645) );
  INV_X1 NOT_6551( .ZN(g19145), .A(II25334) );
  INV_X1 NOT_6552( .ZN(II25338), .A(g17746) );
  INV_X1 NOT_6553( .ZN(g19147), .A(II25338) );
  INV_X1 NOT_6554( .ZN(II25344), .A(g17847) );
  INV_X1 NOT_6555( .ZN(g19151), .A(II25344) );
  INV_X1 NOT_6556( .ZN(II25351), .A(g17959) );
  INV_X1 NOT_6557( .ZN(g19156), .A(II25351) );
  INV_X1 NOT_6558( .ZN(II25355), .A(g18669) );
  INV_X1 NOT_6559( .ZN(g19158), .A(II25355) );
  INV_X1 NOT_6560( .ZN(II25358), .A(g18678) );
  INV_X1 NOT_6561( .ZN(g19159), .A(II25358) );
  INV_X1 NOT_6562( .ZN(II25365), .A(g18707) );
  INV_X1 NOT_6563( .ZN(g19164), .A(II25365) );
  INV_X1 NOT_6564( .ZN(II25371), .A(g18719) );
  INV_X1 NOT_6565( .ZN(g19168), .A(II25371) );
  INV_X1 NOT_6566( .ZN(II25374), .A(g18726) );
  INV_X1 NOT_6567( .ZN(g19169), .A(II25374) );
  INV_X1 NOT_6568( .ZN(II25377), .A(g18743) );
  INV_X1 NOT_6569( .ZN(g19170), .A(II25377) );
  INV_X2 NOT_6570( .ZN(II25383), .A(g18755) );
  INV_X2 NOT_6571( .ZN(g19174), .A(II25383) );
  INV_X1 NOT_6572( .ZN(II25386), .A(g18763) );
  INV_X1 NOT_6573( .ZN(g19175), .A(II25386) );
  INV_X1 NOT_6574( .ZN(II25389), .A(g18780) );
  INV_X1 NOT_6575( .ZN(g19176), .A(II25389) );
  INV_X1 NOT_6576( .ZN(II25395), .A(g18782) );
  INV_X1 NOT_6577( .ZN(g19180), .A(II25395) );
  INV_X1 NOT_6578( .ZN(II25399), .A(g18794) );
  INV_X1 NOT_6579( .ZN(g19182), .A(II25399) );
  INV_X1 NOT_6580( .ZN(II25402), .A(g18821) );
  INV_X1 NOT_6581( .ZN(g19183), .A(II25402) );
  INV_X1 NOT_6582( .ZN(II25406), .A(g18804) );
  INV_X1 NOT_6583( .ZN(g19185), .A(II25406) );
  INV_X1 NOT_6584( .ZN(II25412), .A(g18820) );
  INV_X1 NOT_6585( .ZN(g19189), .A(II25412) );
  INV_X1 NOT_6586( .ZN(II25415), .A(g18835) );
  INV_X1 NOT_6587( .ZN(g19190), .A(II25415) );
  INV_X1 NOT_6588( .ZN(II25423), .A(g18852) );
  INV_X1 NOT_6589( .ZN(g19196), .A(II25423) );
  INV_X1 NOT_6590( .ZN(II25426), .A(g18836) );
  INV_X1 NOT_6591( .ZN(g19197), .A(II25426) );
  INV_X1 NOT_6592( .ZN(II25429), .A(g18975) );
  INV_X1 NOT_6593( .ZN(g19198), .A(II25429) );
  INV_X1 NOT_6594( .ZN(II25432), .A(g18837) );
  INV_X1 NOT_6595( .ZN(g19199), .A(II25432) );
  INV_X1 NOT_6596( .ZN(II25442), .A(g18866) );
  INV_X1 NOT_6597( .ZN(g19207), .A(II25442) );
  INV_X1 NOT_6598( .ZN(II25445), .A(g18968) );
  INV_X1 NOT_6599( .ZN(g19208), .A(II25445) );
  INV_X1 NOT_6600( .ZN(II25456), .A(g18883) );
  INV_X1 NOT_6601( .ZN(g19217), .A(II25456) );
  INV_X1 NOT_6602( .ZN(II25459), .A(g18867) );
  INV_X1 NOT_6603( .ZN(g19218), .A(II25459) );
  INV_X1 NOT_6604( .ZN(II25463), .A(g18868) );
  INV_X1 NOT_6605( .ZN(g19220), .A(II25463) );
  INV_X1 NOT_6606( .ZN(II25474), .A(g18885) );
  INV_X1 NOT_6607( .ZN(g19229), .A(II25474) );
  INV_X1 NOT_6608( .ZN(II25486), .A(g18754) );
  INV_X1 NOT_6609( .ZN(g19237), .A(II25486) );
  INV_X1 NOT_6610( .ZN(II25489), .A(g18906) );
  INV_X1 NOT_6611( .ZN(g19238), .A(II25489) );
  INV_X1 NOT_6612( .ZN(II25492), .A(g18907) );
  INV_X1 NOT_6613( .ZN(g19239), .A(II25492) );
  INV_X1 NOT_6614( .ZN(II25506), .A(g18781) );
  INV_X1 NOT_6615( .ZN(g19247), .A(II25506) );
  INV_X1 NOT_6616( .ZN(II25510), .A(g18542) );
  INV_X1 NOT_6617( .ZN(g19249), .A(II25510) );
  INV_X1 NOT_6618( .ZN(g19251), .A(g16540) );
  INV_X1 NOT_6619( .ZN(II25525), .A(g18803) );
  INV_X1 NOT_6620( .ZN(g19258), .A(II25525) );
  INV_X1 NOT_6621( .ZN(II25528), .A(g18942) );
  INV_X1 NOT_6622( .ZN(g19259), .A(II25528) );
  INV_X1 NOT_6623( .ZN(g19265), .A(g16572) );
  INV_X1 NOT_6624( .ZN(II25557), .A(g18957) );
  INV_X1 NOT_6625( .ZN(g19270), .A(II25557) );
  INV_X1 NOT_6626( .ZN(II25567), .A(g17186) );
  INV_X1 NOT_6627( .ZN(g19272), .A(II25567) );
  INV_X1 NOT_6628( .ZN(g19280), .A(g16596) );
  INV_X1 NOT_6629( .ZN(g19287), .A(g16608) );
  INV_X1 NOT_6630( .ZN(II25612), .A(g17197) );
  INV_X1 NOT_6631( .ZN(g19291), .A(II25612) );
  INV_X1 NOT_6632( .ZN(g19299), .A(g16616) );
  INV_X1 NOT_6633( .ZN(g19301), .A(g16622) );
  INV_X1 NOT_6634( .ZN(g19302), .A(g17025) );
  INV_X2 NOT_6635( .ZN(g19305), .A(g16626) );
  INV_X2 NOT_6636( .ZN(II25660), .A(g17204) );
  INV_X1 NOT_6637( .ZN(g19309), .A(II25660) );
  INV_X1 NOT_6638( .ZN(g19319), .A(g16633) );
  INV_X1 NOT_6639( .ZN(g19322), .A(g16636) );
  INV_X1 NOT_6640( .ZN(g19323), .A(g17059) );
  INV_X1 NOT_6641( .ZN(g19326), .A(g16640) );
  INV_X1 NOT_6642( .ZN(II25717), .A(g17209) );
  INV_X1 NOT_6643( .ZN(g19330), .A(II25717) );
  INV_X1 NOT_6644( .ZN(II25728), .A(g17118) );
  INV_X1 NOT_6645( .ZN(g19335), .A(II25728) );
  INV_X1 NOT_6646( .ZN(g19346), .A(g16644) );
  INV_X1 NOT_6647( .ZN(g19349), .A(g16647) );
  INV_X1 NOT_6648( .ZN(g19350), .A(g17094) );
  INV_X1 NOT_6649( .ZN(g19353), .A(g16651) );
  INV_X1 NOT_6650( .ZN(II25768), .A(g17139) );
  INV_X1 NOT_6651( .ZN(g19358), .A(II25768) );
  INV_X1 NOT_6652( .ZN(II25778), .A(g17145) );
  INV_X1 NOT_6653( .ZN(g19369), .A(II25778) );
  INV_X1 NOT_6654( .ZN(g19380), .A(g16656) );
  INV_X1 NOT_6655( .ZN(g19383), .A(g16659) );
  INV_X1 NOT_6656( .ZN(g19384), .A(g17132) );
  INV_X1 NOT_6657( .ZN(g19387), .A(g16567) );
  INV_X1 NOT_6658( .ZN(g19388), .A(g17139) );
  INV_X1 NOT_6659( .ZN(II25816), .A(g17162) );
  INV_X1 NOT_6660( .ZN(g19390), .A(II25816) );
  INV_X1 NOT_6661( .ZN(II25826), .A(g17168) );
  INV_X1 NOT_6662( .ZN(g19401), .A(II25826) );
  INV_X1 NOT_6663( .ZN(g19412), .A(g16673) );
  INV_X1 NOT_6664( .ZN(g19415), .A(g16676) );
  INV_X1 NOT_6665( .ZN(g19417), .A(g16591) );
  INV_X1 NOT_6666( .ZN(g19418), .A(g17162) );
  INV_X1 NOT_6667( .ZN(II25862), .A(g17177) );
  INV_X1 NOT_6668( .ZN(g19420), .A(II25862) );
  INV_X1 NOT_6669( .ZN(II25872), .A(g17183) );
  INV_X1 NOT_6670( .ZN(g19431), .A(II25872) );
  INV_X1 NOT_6671( .ZN(g19441), .A(g17213) );
  INV_X1 NOT_6672( .ZN(g19444), .A(g17985) );
  INV_X1 NOT_6673( .ZN(g19448), .A(g16694) );
  INV_X1 NOT_6674( .ZN(g19452), .A(g16702) );
  INV_X1 NOT_6675( .ZN(g19454), .A(g16611) );
  INV_X1 NOT_6676( .ZN(g19455), .A(g17177) );
  INV_X1 NOT_6677( .ZN(II25904), .A(g17194) );
  INV_X1 NOT_6678( .ZN(g19457), .A(II25904) );
  INV_X1 NOT_6679( .ZN(g19467), .A(g16719) );
  INV_X1 NOT_6680( .ZN(g19468), .A(g17216) );
  INV_X1 NOT_6681( .ZN(g19471), .A(g18102) );
  INV_X1 NOT_6682( .ZN(g19475), .A(g16725) );
  INV_X1 NOT_6683( .ZN(g19479), .A(g16733) );
  INV_X1 NOT_6684( .ZN(g19481), .A(g16629) );
  INV_X1 NOT_6685( .ZN(g19482), .A(g17194) );
  INV_X1 NOT_6686( .ZN(g19483), .A(g16758) );
  INV_X1 NOT_6687( .ZN(g19484), .A(g16867) );
  INV_X1 NOT_6688( .ZN(g19490), .A(g16761) );
  INV_X1 NOT_6689( .ZN(g19491), .A(g17219) );
  INV_X1 NOT_6690( .ZN(g19494), .A(g18218) );
  INV_X1 NOT_6691( .ZN(g19498), .A(g16767) );
  INV_X1 NOT_6692( .ZN(g19502), .A(g16775) );
  INV_X1 NOT_6693( .ZN(g19504), .A(g16785) );
  INV_X1 NOT_6694( .ZN(g19505), .A(g16895) );
  INV_X1 NOT_6695( .ZN(g19511), .A(g16788) );
  INV_X1 NOT_6696( .ZN(g19512), .A(g17221) );
  INV_X1 NOT_6697( .ZN(g19515), .A(g18325) );
  INV_X1 NOT_6698( .ZN(g19519), .A(g16794) );
  INV_X1 NOT_6699( .ZN(g19523), .A(g16814) );
  INV_X1 NOT_6700( .ZN(g19524), .A(g16924) );
  INV_X1 NOT_6701( .ZN(g19530), .A(g16817) );
  INV_X1 NOT_6702( .ZN(g19533), .A(g16832) );
  INV_X1 NOT_6703( .ZN(g19534), .A(g16954) );
  INV_X1 NOT_6704( .ZN(II25966), .A(g16654) );
  INV_X1 NOT_6705( .ZN(g19543), .A(II25966) );
  INV_X1 NOT_6706( .ZN(II25971), .A(g16671) );
  INV_X1 NOT_6707( .ZN(g19546), .A(II25971) );
  INV_X1 NOT_6708( .ZN(II25977), .A(g16692) );
  INV_X1 NOT_6709( .ZN(g19550), .A(II25977) );
  INV_X1 NOT_6710( .ZN(II25985), .A(g16718) );
  INV_X1 NOT_6711( .ZN(g19556), .A(II25985) );
  INV_X1 NOT_6712( .ZN(II25994), .A(g16860) );
  INV_X1 NOT_6713( .ZN(g19563), .A(II25994) );
  INV_X1 NOT_6714( .ZN(II26006), .A(g16866) );
  INV_X1 NOT_6715( .ZN(g19573), .A(II26006) );
  INV_X1 NOT_6716( .ZN(g19577), .A(g16881) );
  INV_X1 NOT_6717( .ZN(g19578), .A(g16884) );
  INV_X1 NOT_6718( .ZN(II26025), .A(g16803) );
  INV_X1 NOT_6719( .ZN(g19595), .A(II26025) );
  INV_X1 NOT_6720( .ZN(II26028), .A(g16566) );
  INV_X1 NOT_6721( .ZN(g19596), .A(II26028) );
  INV_X1 NOT_6722( .ZN(g19607), .A(g16910) );
  INV_X1 NOT_6723( .ZN(g19608), .A(g16913) );
  INV_X1 NOT_6724( .ZN(II26051), .A(g16824) );
  INV_X1 NOT_6725( .ZN(g19622), .A(II26051) );
  INV_X1 NOT_6726( .ZN(g19640), .A(g16940) );
  INV_X1 NOT_6727( .ZN(g19641), .A(g16943) );
  INV_X1 NOT_6728( .ZN(II26078), .A(g16835) );
  INV_X1 NOT_6729( .ZN(g19652), .A(II26078) );
  INV_X1 NOT_6730( .ZN(II26085), .A(g18085) );
  INV_X1 NOT_6731( .ZN(g19657), .A(II26085) );
  INV_X1 NOT_6732( .ZN(g19680), .A(g16971) );
  INV_X1 NOT_6733( .ZN(g19681), .A(g16974) );
  INV_X1 NOT_6734( .ZN(II26112), .A(g16844) );
  INV_X1 NOT_6735( .ZN(g19689), .A(II26112) );
  INV_X1 NOT_6736( .ZN(II26115), .A(g16845) );
  INV_X1 NOT_6737( .ZN(g19690), .A(II26115) );
  INV_X1 NOT_6738( .ZN(II26123), .A(g17503) );
  INV_X1 NOT_6739( .ZN(g19696), .A(II26123) );
  INV_X1 NOT_6740( .ZN(II26134), .A(g18201) );
  INV_X2 NOT_6741( .ZN(g19705), .A(II26134) );
  INV_X2 NOT_6742( .ZN(II26154), .A(g16851) );
  INV_X1 NOT_6743( .ZN(g19725), .A(II26154) );
  INV_X1 NOT_6744( .ZN(II26171), .A(g17594) );
  INV_X1 NOT_6745( .ZN(g19740), .A(II26171) );
  INV_X1 NOT_6746( .ZN(II26182), .A(g18308) );
  INV_X1 NOT_6747( .ZN(g19749), .A(II26182) );
  INV_X1 NOT_6748( .ZN(II26195), .A(g16853) );
  INV_X1 NOT_6749( .ZN(g19762), .A(II26195) );
  INV_X1 NOT_6750( .ZN(II26198), .A(g16854) );
  INV_X1 NOT_6751( .ZN(g19763), .A(II26198) );
  INV_X1 NOT_6752( .ZN(II26220), .A(g17691) );
  INV_X1 NOT_6753( .ZN(g19783), .A(II26220) );
  INV_X1 NOT_6754( .ZN(II26231), .A(g18401) );
  INV_X1 NOT_6755( .ZN(g19792), .A(II26231) );
  INV_X1 NOT_6756( .ZN(II26237), .A(g16857) );
  INV_X1 NOT_6757( .ZN(g19798), .A(II26237) );
  INV_X1 NOT_6758( .ZN(II26266), .A(g17791) );
  INV_X1 NOT_6759( .ZN(g19825), .A(II26266) );
  INV_X1 NOT_6760( .ZN(g19830), .A(g18886) );
  INV_X1 NOT_6761( .ZN(II26276), .A(g16861) );
  INV_X1 NOT_6762( .ZN(g19838), .A(II26276) );
  INV_X1 NOT_6763( .ZN(II26334), .A(g18977) );
  INV_X1 NOT_6764( .ZN(g19890), .A(II26334) );
  INV_X1 NOT_6765( .ZN(II26337), .A(g16880) );
  INV_X1 NOT_6766( .ZN(g19893), .A(II26337) );
  INV_X1 NOT_6767( .ZN(II26340), .A(g17025) );
  INV_X1 NOT_6768( .ZN(g19894), .A(II26340) );
  INV_X1 NOT_6769( .ZN(II26365), .A(g18626) );
  INV_X1 NOT_6770( .ZN(g19915), .A(II26365) );
  INV_X1 NOT_6771( .ZN(g19918), .A(g18646) );
  INV_X1 NOT_6772( .ZN(II26369), .A(g17059) );
  INV_X1 NOT_6773( .ZN(g19919), .A(II26369) );
  INV_X1 NOT_6774( .ZN(g19933), .A(g18548) );
  INV_X1 NOT_6775( .ZN(II26388), .A(g17094) );
  INV_X1 NOT_6776( .ZN(g19934), .A(II26388) );
  INV_X1 NOT_6777( .ZN(II26401), .A(g17012) );
  INV_X1 NOT_6778( .ZN(g19945), .A(II26401) );
  INV_X1 NOT_6779( .ZN(g19948), .A(g17896) );
  INV_X1 NOT_6780( .ZN(g19950), .A(g18598) );
  INV_X1 NOT_6781( .ZN(II26407), .A(g17132) );
  INV_X1 NOT_6782( .ZN(g19951), .A(II26407) );
  INV_X1 NOT_6783( .ZN(II26413), .A(g16643) );
  INV_X1 NOT_6784( .ZN(g19957), .A(II26413) );
  INV_X1 NOT_6785( .ZN(II26420), .A(g17042) );
  INV_X1 NOT_6786( .ZN(g19972), .A(II26420) );
  INV_X1 NOT_6787( .ZN(g19975), .A(g18007) );
  INV_X1 NOT_6788( .ZN(g19977), .A(g18630) );
  INV_X1 NOT_6789( .ZN(II26426), .A(g16536) );
  INV_X1 NOT_6790( .ZN(g19978), .A(II26426) );
  INV_X1 NOT_6791( .ZN(II26437), .A(g16655) );
  INV_X1 NOT_6792( .ZN(g19987), .A(II26437) );
  INV_X1 NOT_6793( .ZN(II26444), .A(g17076) );
  INV_X1 NOT_6794( .ZN(g20002), .A(II26444) );
  INV_X1 NOT_6795( .ZN(g20005), .A(g18124) );
  INV_X1 NOT_6796( .ZN(g20007), .A(g18639) );
  INV_X1 NOT_6797( .ZN(II26458), .A(g17985) );
  INV_X1 NOT_6798( .ZN(g20016), .A(II26458) );
  INV_X1 NOT_6799( .ZN(II26469), .A(g16672) );
  INV_X1 NOT_6800( .ZN(g20025), .A(II26469) );
  INV_X1 NOT_6801( .ZN(II26476), .A(g17111) );
  INV_X1 NOT_6802( .ZN(g20040), .A(II26476) );
  INV_X1 NOT_6803( .ZN(g20043), .A(g18240) );
  INV_X1 NOT_6804( .ZN(II26481), .A(g18590) );
  INV_X1 NOT_6805( .ZN(g20045), .A(II26481) );
  INV_X1 NOT_6806( .ZN(II26494), .A(g18102) );
  INV_X1 NOT_6807( .ZN(g20058), .A(II26494) );
  INV_X1 NOT_6808( .ZN(II26505), .A(g16693) );
  INV_X1 NOT_6809( .ZN(g20067), .A(II26505) );
  INV_X1 NOT_6810( .ZN(II26512), .A(g16802) );
  INV_X1 NOT_6811( .ZN(g20082), .A(II26512) );
  INV_X1 NOT_6812( .ZN(g20083), .A(g17968) );
  INV_X1 NOT_6813( .ZN(II26535), .A(g18218) );
  INV_X1 NOT_6814( .ZN(g20099), .A(II26535) );
  INV_X1 NOT_6815( .ZN(II26545), .A(g16823) );
  INV_X1 NOT_6816( .ZN(g20105), .A(II26545) );
  INV_X1 NOT_6817( .ZN(II26574), .A(g18325) );
  INV_X1 NOT_6818( .ZN(g20124), .A(II26574) );
  INV_X1 NOT_6819( .ZN(g20127), .A(g18623) );
  INV_X1 NOT_6820( .ZN(g20140), .A(g16830) );
  INV_X1 NOT_6821( .ZN(g20163), .A(g17973) );
  INV_X1 NOT_6822( .ZN(II26612), .A(g17645) );
  INV_X1 NOT_6823( .ZN(g20164), .A(II26612) );
  INV_X1 NOT_6824( .ZN(g20178), .A(g16842) );
  INV_X1 NOT_6825( .ZN(g20193), .A(g18691) );
  INV_X1 NOT_6826( .ZN(II26642), .A(g17746) );
  INV_X1 NOT_6827( .ZN(g20198), .A(II26642) );
  INV_X1 NOT_6828( .ZN(g20212), .A(g16848) );
  INV_X1 NOT_6829( .ZN(g20223), .A(g18727) );
  INV_X1 NOT_6830( .ZN(II26664), .A(g17847) );
  INV_X1 NOT_6831( .ZN(g20228), .A(II26664) );
  INV_X1 NOT_6832( .ZN(g20242), .A(g16852) );
  INV_X1 NOT_6833( .ZN(g20250), .A(g18764) );
  INV_X1 NOT_6834( .ZN(II26679), .A(g17959) );
  INV_X1 NOT_6835( .ZN(g20255), .A(II26679) );
  INV_X1 NOT_6836( .ZN(g20269), .A(g17230) );
  INV_X1 NOT_6837( .ZN(g20273), .A(g18795) );
  INV_X1 NOT_6838( .ZN(g20278), .A(g17237) );
  INV_X1 NOT_6839( .ZN(g20279), .A(g17240) );
  INV_X1 NOT_6840( .ZN(g20281), .A(g17243) );
  INV_X1 NOT_6841( .ZN(g20286), .A(g17249) );
  INV_X1 NOT_6842( .ZN(g20287), .A(g17252) );
  INV_X1 NOT_6843( .ZN(g20288), .A(g17255) );
  INV_X1 NOT_6844( .ZN(g20289), .A(g17259) );
  INV_X1 NOT_6845( .ZN(g20290), .A(g17262) );
  INV_X1 NOT_6846( .ZN(g20292), .A(g17265) );
  INV_X1 NOT_6847( .ZN(II26714), .A(g17720) );
  INV_X1 NOT_6848( .ZN(g20295), .A(II26714) );
  INV_X1 NOT_6849( .ZN(g20296), .A(g17272) );
  INV_X1 NOT_6850( .ZN(g20297), .A(g17275) );
  INV_X1 NOT_6851( .ZN(g20298), .A(g17278) );
  INV_X1 NOT_6852( .ZN(g20302), .A(g17282) );
  INV_X1 NOT_6853( .ZN(g20303), .A(g17285) );
  INV_X1 NOT_6854( .ZN(g20304), .A(g17288) );
  INV_X1 NOT_6855( .ZN(g20305), .A(g17291) );
  INV_X1 NOT_6856( .ZN(g20306), .A(g17294) );
  INV_X1 NOT_6857( .ZN(g20308), .A(g17297) );
  INV_X1 NOT_6858( .ZN(g20311), .A(g17304) );
  INV_X1 NOT_6859( .ZN(g20312), .A(g17307) );
  INV_X1 NOT_6860( .ZN(g20313), .A(g17310) );
  INV_X1 NOT_6861( .ZN(g20315), .A(g17315) );
  INV_X1 NOT_6862( .ZN(g20316), .A(g17318) );
  INV_X1 NOT_6863( .ZN(g20317), .A(g17321) );
  INV_X1 NOT_6864( .ZN(g20321), .A(g17324) );
  INV_X1 NOT_6865( .ZN(g20322), .A(g17327) );
  INV_X1 NOT_6866( .ZN(g20323), .A(g17330) );
  INV_X1 NOT_6867( .ZN(g20324), .A(g17333) );
  INV_X1 NOT_6868( .ZN(g20325), .A(g17336) );
  INV_X1 NOT_6869( .ZN(g20327), .A(g17342) );
  INV_X1 NOT_6870( .ZN(g20328), .A(g17345) );
  INV_X1 NOT_6871( .ZN(g20329), .A(g17348) );
  INV_X1 NOT_6872( .ZN(g20330), .A(g17354) );
  INV_X1 NOT_6873( .ZN(g20331), .A(g17357) );
  INV_X1 NOT_6874( .ZN(g20332), .A(g17360) );
  INV_X1 NOT_6875( .ZN(g20334), .A(g17363) );
  INV_X1 NOT_6876( .ZN(g20335), .A(g17366) );
  INV_X1 NOT_6877( .ZN(g20336), .A(g17369) );
  INV_X1 NOT_6878( .ZN(g20340), .A(g17372) );
  INV_X1 NOT_6879( .ZN(g20341), .A(g17375) );
  INV_X1 NOT_6880( .ZN(g20342), .A(g17378) );
  INV_X1 NOT_6881( .ZN(g20344), .A(g17384) );
  INV_X1 NOT_6882( .ZN(g20345), .A(g17387) );
  INV_X1 NOT_6883( .ZN(g20346), .A(g17390) );
  INV_X1 NOT_6884( .ZN(g20347), .A(g17399) );
  INV_X1 NOT_6885( .ZN(g20348), .A(g17402) );
  INV_X1 NOT_6886( .ZN(g20349), .A(g17405) );
  INV_X1 NOT_6887( .ZN(g20350), .A(g17410) );
  INV_X1 NOT_6888( .ZN(g20351), .A(g17413) );
  INV_X1 NOT_6889( .ZN(g20352), .A(g17416) );
  INV_X1 NOT_6890( .ZN(g20354), .A(g17419) );
  INV_X1 NOT_6891( .ZN(g20355), .A(g17422) );
  INV_X1 NOT_6892( .ZN(g20356), .A(g17425) );
  INV_X1 NOT_6893( .ZN(II26777), .A(g17222) );
  INV_X1 NOT_6894( .ZN(g20360), .A(II26777) );
  INV_X1 NOT_6895( .ZN(g20361), .A(g17430) );
  INV_X1 NOT_6896( .ZN(g20362), .A(g17433) );
  INV_X1 NOT_6897( .ZN(g20363), .A(g17436) );
  INV_X1 NOT_6898( .ZN(g20364), .A(g17439) );
  INV_X1 NOT_6899( .ZN(g20365), .A(g17442) );
  INV_X1 NOT_6900( .ZN(g20366), .A(g17451) );
  INV_X1 NOT_6901( .ZN(g20367), .A(g17454) );
  INV_X1 NOT_6902( .ZN(g20368), .A(g17457) );
  INV_X1 NOT_6903( .ZN(g20369), .A(g17465) );
  INV_X1 NOT_6904( .ZN(g20370), .A(g17468) );
  INV_X1 NOT_6905( .ZN(g20371), .A(g17471) );
  INV_X1 NOT_6906( .ZN(g20372), .A(g17476) );
  INV_X1 NOT_6907( .ZN(g20373), .A(g17479) );
  INV_X1 NOT_6908( .ZN(g20374), .A(g17482) );
  INV_X1 NOT_6909( .ZN(II26796), .A(g17224) );
  INV_X1 NOT_6910( .ZN(g20377), .A(II26796) );
  INV_X1 NOT_6911( .ZN(g20378), .A(g17487) );
  INV_X1 NOT_6912( .ZN(g20379), .A(g17490) );
  INV_X1 NOT_6913( .ZN(g20380), .A(g17493) );
  INV_X1 NOT_6914( .ZN(g20381), .A(g17496) );
  INV_X1 NOT_6915( .ZN(g20382), .A(g17500) );
  INV_X1 NOT_6916( .ZN(g20383), .A(g17503) );
  INV_X1 NOT_6917( .ZN(g20384), .A(g17511) );
  INV_X1 NOT_6918( .ZN(g20385), .A(g17514) );
  INV_X1 NOT_6919( .ZN(g20386), .A(g17517) );
  INV_X1 NOT_6920( .ZN(g20387), .A(g17520) );
  INV_X1 NOT_6921( .ZN(g20388), .A(g17523) );
  INV_X1 NOT_6922( .ZN(g20389), .A(g17531) );
  INV_X1 NOT_6923( .ZN(g20390), .A(g17534) );
  INV_X1 NOT_6924( .ZN(g20391), .A(g17537) );
  INV_X1 NOT_6925( .ZN(g20392), .A(g17545) );
  INV_X1 NOT_6926( .ZN(g20393), .A(g17548) );
  INV_X1 NOT_6927( .ZN(g20394), .A(g17551) );
  INV_X1 NOT_6928( .ZN(II26816), .A(g17225) );
  INV_X1 NOT_6929( .ZN(g20395), .A(II26816) );
  INV_X1 NOT_6930( .ZN(II26819), .A(g17226) );
  INV_X1 NOT_6931( .ZN(g20396), .A(II26819) );
  INV_X1 NOT_6932( .ZN(g20397), .A(g17557) );
  INV_X1 NOT_6933( .ZN(g20398), .A(g17560) );
  INV_X1 NOT_6934( .ZN(g20399), .A(g17563) );
  INV_X1 NOT_6935( .ZN(g20400), .A(g17567) );
  INV_X1 NOT_6936( .ZN(g20401), .A(g17570) );
  INV_X2 NOT_6937( .ZN(g20402), .A(g17573) );
  INV_X2 NOT_6938( .ZN(g20403), .A(g17579) );
  INV_X1 NOT_6939( .ZN(g20404), .A(g17582) );
  INV_X1 NOT_6940( .ZN(g20405), .A(g17585) );
  INV_X1 NOT_6941( .ZN(g20406), .A(g17588) );
  INV_X1 NOT_6942( .ZN(g20407), .A(g17591) );
  INV_X1 NOT_6943( .ZN(g20408), .A(g17594) );
  INV_X1 NOT_6944( .ZN(g20409), .A(g17601) );
  INV_X1 NOT_6945( .ZN(g20410), .A(g17604) );
  INV_X1 NOT_6946( .ZN(g20411), .A(g17607) );
  INV_X1 NOT_6947( .ZN(g20412), .A(g17610) );
  INV_X1 NOT_6948( .ZN(g20413), .A(g17613) );
  INV_X1 NOT_6949( .ZN(g20414), .A(g17621) );
  INV_X1 NOT_6950( .ZN(g20415), .A(g17624) );
  INV_X1 NOT_6951( .ZN(g20416), .A(g17627) );
  INV_X1 NOT_6952( .ZN(II26843), .A(g17228) );
  INV_X1 NOT_6953( .ZN(g20418), .A(II26843) );
  INV_X1 NOT_6954( .ZN(II26846), .A(g17229) );
  INV_X1 NOT_6955( .ZN(g20419), .A(II26846) );
  INV_X1 NOT_6956( .ZN(g20420), .A(g17637) );
  INV_X1 NOT_6957( .ZN(g20421), .A(g17649) );
  INV_X1 NOT_6958( .ZN(g20422), .A(g17655) );
  INV_X1 NOT_6959( .ZN(g20423), .A(g17658) );
  INV_X1 NOT_6960( .ZN(g20424), .A(g17661) );
  INV_X1 NOT_6961( .ZN(g20425), .A(g17664) );
  INV_X1 NOT_6962( .ZN(g20426), .A(g17667) );
  INV_X1 NOT_6963( .ZN(g20427), .A(g17670) );
  INV_X1 NOT_6964( .ZN(g20428), .A(g17676) );
  INV_X1 NOT_6965( .ZN(g20429), .A(g17679) );
  INV_X1 NOT_6966( .ZN(g20430), .A(g17682) );
  INV_X1 NOT_6967( .ZN(g20431), .A(g17685) );
  INV_X1 NOT_6968( .ZN(g20432), .A(g17688) );
  INV_X1 NOT_6969( .ZN(g20433), .A(g17691) );
  INV_X1 NOT_6970( .ZN(g20434), .A(g17698) );
  INV_X1 NOT_6971( .ZN(g20435), .A(g17701) );
  INV_X1 NOT_6972( .ZN(g20436), .A(g17704) );
  INV_X1 NOT_6973( .ZN(g20437), .A(g17707) );
  INV_X1 NOT_6974( .ZN(g20438), .A(g17710) );
  INV_X1 NOT_6975( .ZN(II26868), .A(g17234) );
  INV_X1 NOT_6976( .ZN(g20439), .A(II26868) );
  INV_X1 NOT_6977( .ZN(II26871), .A(g17235) );
  INV_X1 NOT_6978( .ZN(g20440), .A(II26871) );
  INV_X1 NOT_6979( .ZN(II26874), .A(g17236) );
  INV_X1 NOT_6980( .ZN(g20441), .A(II26874) );
  INV_X1 NOT_6981( .ZN(g20442), .A(g17738) );
  INV_X1 NOT_6982( .ZN(g20443), .A(g17749) );
  INV_X1 NOT_6983( .ZN(g20444), .A(g17755) );
  INV_X1 NOT_6984( .ZN(g20445), .A(g17758) );
  INV_X1 NOT_6985( .ZN(g20446), .A(g17761) );
  INV_X1 NOT_6986( .ZN(g20447), .A(g17764) );
  INV_X1 NOT_6987( .ZN(g20448), .A(g17767) );
  INV_X1 NOT_6988( .ZN(g20449), .A(g17770) );
  INV_X1 NOT_6989( .ZN(g20450), .A(g17776) );
  INV_X1 NOT_6990( .ZN(g20451), .A(g17779) );
  INV_X1 NOT_6991( .ZN(g20452), .A(g17782) );
  INV_X1 NOT_6992( .ZN(g20453), .A(g17785) );
  INV_X1 NOT_6993( .ZN(g20454), .A(g17788) );
  INV_X1 NOT_6994( .ZN(g20455), .A(g17791) );
  INV_X1 NOT_6995( .ZN(g20456), .A(g17799) );
  INV_X1 NOT_6996( .ZN(II26892), .A(g17246) );
  INV_X1 NOT_6997( .ZN(g20457), .A(II26892) );
  INV_X1 NOT_6998( .ZN(II26895), .A(g17247) );
  INV_X1 NOT_6999( .ZN(g20458), .A(II26895) );
  INV_X1 NOT_7000( .ZN(II26898), .A(g17248) );
  INV_X1 NOT_7001( .ZN(g20459), .A(II26898) );
  INV_X1 NOT_7002( .ZN(g20461), .A(g17839) );
  INV_X1 NOT_7003( .ZN(g20462), .A(g17850) );
  INV_X1 NOT_7004( .ZN(g20463), .A(g17856) );
  INV_X1 NOT_7005( .ZN(g20464), .A(g17859) );
  INV_X1 NOT_7006( .ZN(g20465), .A(g17862) );
  INV_X1 NOT_7007( .ZN(g20466), .A(g17865) );
  INV_X1 NOT_7008( .ZN(g20467), .A(g17868) );
  INV_X1 NOT_7009( .ZN(g20468), .A(g17871) );
  INV_X1 NOT_7010( .ZN(II26910), .A(g17269) );
  INV_X1 NOT_7011( .ZN(g20469), .A(II26910) );
  INV_X1 NOT_7012( .ZN(II26913), .A(g17270) );
  INV_X1 NOT_7013( .ZN(g20470), .A(II26913) );
  INV_X1 NOT_7014( .ZN(II26916), .A(g17271) );
  INV_X1 NOT_7015( .ZN(g20471), .A(II26916) );
  INV_X1 NOT_7016( .ZN(g20476), .A(g17951) );
  INV_X1 NOT_7017( .ZN(g20477), .A(g17962) );
  INV_X1 NOT_7018( .ZN(II26923), .A(g17302) );
  INV_X1 NOT_7019( .ZN(g20478), .A(II26923) );
  INV_X1 NOT_7020( .ZN(II26926), .A(g17303) );
  INV_X1 NOT_7021( .ZN(g20479), .A(II26926) );
  INV_X1 NOT_7022( .ZN(II26931), .A(g17340) );
  INV_X1 NOT_7023( .ZN(g20484), .A(II26931) );
  INV_X1 NOT_7024( .ZN(II26934), .A(g17341) );
  INV_X1 NOT_7025( .ZN(g20485), .A(II26934) );
  INV_X1 NOT_7026( .ZN(g20490), .A(g18166) );
  INV_X1 NOT_7027( .ZN(II26940), .A(g17383) );
  INV_X1 NOT_7028( .ZN(g20491), .A(II26940) );
  INV_X1 NOT_7029( .ZN(g20496), .A(g18258) );
  INV_X1 NOT_7030( .ZN(II26947), .A(g17429) );
  INV_X1 NOT_7031( .ZN(g20498), .A(II26947) );
  INV_X1 NOT_7032( .ZN(g20500), .A(g18278) );
  INV_X1 NOT_7033( .ZN(g20501), .A(g18334) );
  INV_X1 NOT_7034( .ZN(g20504), .A(g18355) );
  INV_X1 NOT_7035( .ZN(g20505), .A(g18371) );
  INV_X1 NOT_7036( .ZN(g20507), .A(g18351) );
  INV_X1 NOT_7037( .ZN(II26960), .A(g16884) );
  INV_X1 NOT_7038( .ZN(g20513), .A(II26960) );
  INV_X1 NOT_7039( .ZN(g20516), .A(g18432) );
  INV_X1 NOT_7040( .ZN(g20517), .A(g18450) );
  INV_X1 NOT_7041( .ZN(g20518), .A(g18466) );
  INV_X1 NOT_7042( .ZN(II26966), .A(g17051) );
  INV_X1 NOT_7043( .ZN(g20519), .A(II26966) );
  INV_X1 NOT_7044( .ZN(g20526), .A(g18446) );
  INV_X1 NOT_7045( .ZN(II26972), .A(g16913) );
  INV_X1 NOT_7046( .ZN(g20531), .A(II26972) );
  INV_X1 NOT_7047( .ZN(g20534), .A(g18505) );
  INV_X1 NOT_7048( .ZN(g20535), .A(g18523) );
  INV_X1 NOT_7049( .ZN(g20536), .A(g18539) );
  INV_X1 NOT_7050( .ZN(II26980), .A(g17086) );
  INV_X1 NOT_7051( .ZN(g20539), .A(II26980) );
  INV_X1 NOT_7052( .ZN(g20545), .A(g18519) );
  INV_X1 NOT_7053( .ZN(II26985), .A(g16943) );
  INV_X1 NOT_7054( .ZN(g20550), .A(II26985) );
  INV_X1 NOT_7055( .ZN(g20553), .A(g18569) );
  INV_X1 NOT_7056( .ZN(g20554), .A(g18587) );
  INV_X1 NOT_7057( .ZN(II26990), .A(g19145) );
  INV_X1 NOT_7058( .ZN(g20555), .A(II26990) );
  INV_X1 NOT_7059( .ZN(II26993), .A(g19159) );
  INV_X1 NOT_7060( .ZN(g20556), .A(II26993) );
  INV_X1 NOT_7061( .ZN(II26996), .A(g19169) );
  INV_X1 NOT_7062( .ZN(g20557), .A(II26996) );
  INV_X1 NOT_7063( .ZN(II26999), .A(g19543) );
  INV_X1 NOT_7064( .ZN(g20558), .A(II26999) );
  INV_X1 NOT_7065( .ZN(II27002), .A(g19147) );
  INV_X1 NOT_7066( .ZN(g20559), .A(II27002) );
  INV_X1 NOT_7067( .ZN(II27005), .A(g19164) );
  INV_X1 NOT_7068( .ZN(g20560), .A(II27005) );
  INV_X1 NOT_7069( .ZN(II27008), .A(g19175) );
  INV_X1 NOT_7070( .ZN(g20561), .A(II27008) );
  INV_X1 NOT_7071( .ZN(II27011), .A(g19546) );
  INV_X1 NOT_7072( .ZN(g20562), .A(II27011) );
  INV_X1 NOT_7073( .ZN(II27014), .A(g19151) );
  INV_X1 NOT_7074( .ZN(g20563), .A(II27014) );
  INV_X1 NOT_7075( .ZN(II27017), .A(g19170) );
  INV_X1 NOT_7076( .ZN(g20564), .A(II27017) );
  INV_X1 NOT_7077( .ZN(II27020), .A(g19182) );
  INV_X1 NOT_7078( .ZN(g20565), .A(II27020) );
  INV_X1 NOT_7079( .ZN(II27023), .A(g19550) );
  INV_X1 NOT_7080( .ZN(g20566), .A(II27023) );
  INV_X1 NOT_7081( .ZN(II27026), .A(g19156) );
  INV_X1 NOT_7082( .ZN(g20567), .A(II27026) );
  INV_X1 NOT_7083( .ZN(II27029), .A(g19176) );
  INV_X1 NOT_7084( .ZN(g20568), .A(II27029) );
  INV_X1 NOT_7085( .ZN(II27032), .A(g19189) );
  INV_X1 NOT_7086( .ZN(g20569), .A(II27032) );
  INV_X1 NOT_7087( .ZN(II27035), .A(g19556) );
  INV_X1 NOT_7088( .ZN(g20570), .A(II27035) );
  INV_X1 NOT_7089( .ZN(II27038), .A(g20082) );
  INV_X1 NOT_7090( .ZN(g20571), .A(II27038) );
  INV_X1 NOT_7091( .ZN(II27041), .A(g19237) );
  INV_X1 NOT_7092( .ZN(g20572), .A(II27041) );
  INV_X1 NOT_7093( .ZN(II27044), .A(g19247) );
  INV_X1 NOT_7094( .ZN(g20573), .A(II27044) );
  INV_X1 NOT_7095( .ZN(II27047), .A(g19258) );
  INV_X1 NOT_7096( .ZN(g20574), .A(II27047) );
  INV_X1 NOT_7097( .ZN(II27050), .A(g19183) );
  INV_X1 NOT_7098( .ZN(g20575), .A(II27050) );
  INV_X1 NOT_7099( .ZN(II27053), .A(g19190) );
  INV_X1 NOT_7100( .ZN(g20576), .A(II27053) );
  INV_X1 NOT_7101( .ZN(II27056), .A(g19196) );
  INV_X1 NOT_7102( .ZN(g20577), .A(II27056) );
  INV_X1 NOT_7103( .ZN(II27059), .A(g19207) );
  INV_X1 NOT_7104( .ZN(g20578), .A(II27059) );
  INV_X1 NOT_7105( .ZN(II27062), .A(g19217) );
  INV_X1 NOT_7106( .ZN(g20579), .A(II27062) );
  INV_X1 NOT_7107( .ZN(II27065), .A(g19270) );
  INV_X1 NOT_7108( .ZN(g20580), .A(II27065) );
  INV_X1 NOT_7109( .ZN(II27068), .A(g19197) );
  INV_X1 NOT_7110( .ZN(g20581), .A(II27068) );
  INV_X1 NOT_7111( .ZN(II27071), .A(g19218) );
  INV_X1 NOT_7112( .ZN(g20582), .A(II27071) );
  INV_X1 NOT_7113( .ZN(II27074), .A(g19238) );
  INV_X1 NOT_7114( .ZN(g20583), .A(II27074) );
  INV_X1 NOT_7115( .ZN(II27077), .A(g19259) );
  INV_X1 NOT_7116( .ZN(g20584), .A(II27077) );
  INV_X1 NOT_7117( .ZN(II27080), .A(g19198) );
  INV_X1 NOT_7118( .ZN(g20585), .A(II27080) );
  INV_X1 NOT_7119( .ZN(II27083), .A(g19208) );
  INV_X1 NOT_7120( .ZN(g20586), .A(II27083) );
  INV_X1 NOT_7121( .ZN(II27086), .A(g19229) );
  INV_X4 NOT_7122( .ZN(g20587), .A(II27086) );
  INV_X4 NOT_7123( .ZN(II27089), .A(g20105) );
  INV_X4 NOT_7124( .ZN(g20588), .A(II27089) );
  INV_X1 NOT_7125( .ZN(II27092), .A(g19174) );
  INV_X1 NOT_7126( .ZN(g20589), .A(II27092) );
  INV_X1 NOT_7127( .ZN(II27095), .A(g19185) );
  INV_X1 NOT_7128( .ZN(g20590), .A(II27095) );
  INV_X1 NOT_7129( .ZN(II27098), .A(g19199) );
  INV_X1 NOT_7130( .ZN(g20591), .A(II27098) );
  INV_X1 NOT_7131( .ZN(II27101), .A(g19220) );
  INV_X1 NOT_7132( .ZN(g20592), .A(II27101) );
  INV_X1 NOT_7133( .ZN(II27104), .A(g19239) );
  INV_X1 NOT_7134( .ZN(g20593), .A(II27104) );
  INV_X1 NOT_7135( .ZN(II27107), .A(g19249) );
  INV_X1 NOT_7136( .ZN(g20594), .A(II27107) );
  INV_X1 NOT_7137( .ZN(II27110), .A(g19622) );
  INV_X1 NOT_7138( .ZN(g20595), .A(II27110) );
  INV_X1 NOT_7139( .ZN(II27113), .A(g19689) );
  INV_X1 NOT_7140( .ZN(g20596), .A(II27113) );
  INV_X1 NOT_7141( .ZN(II27116), .A(g19762) );
  INV_X1 NOT_7142( .ZN(g20597), .A(II27116) );
  INV_X1 NOT_7143( .ZN(II27119), .A(g19563) );
  INV_X1 NOT_7144( .ZN(g20598), .A(II27119) );
  INV_X1 NOT_7145( .ZN(II27122), .A(g19595) );
  INV_X1 NOT_7146( .ZN(g20599), .A(II27122) );
  INV_X1 NOT_7147( .ZN(II27125), .A(g19652) );
  INV_X1 NOT_7148( .ZN(g20600), .A(II27125) );
  INV_X1 NOT_7149( .ZN(II27128), .A(g19725) );
  INV_X1 NOT_7150( .ZN(g20601), .A(II27128) );
  INV_X1 NOT_7151( .ZN(II27131), .A(g19798) );
  INV_X1 NOT_7152( .ZN(g20602), .A(II27131) );
  INV_X1 NOT_7153( .ZN(II27134), .A(g19573) );
  INV_X1 NOT_7154( .ZN(g20603), .A(II27134) );
  INV_X1 NOT_7155( .ZN(II27137), .A(g19596) );
  INV_X1 NOT_7156( .ZN(g20604), .A(II27137) );
  INV_X1 NOT_7157( .ZN(II27140), .A(g19690) );
  INV_X1 NOT_7158( .ZN(g20605), .A(II27140) );
  INV_X1 NOT_7159( .ZN(II27143), .A(g19763) );
  INV_X1 NOT_7160( .ZN(g20606), .A(II27143) );
  INV_X1 NOT_7161( .ZN(II27146), .A(g19838) );
  INV_X1 NOT_7162( .ZN(g20607), .A(II27146) );
  INV_X1 NOT_7163( .ZN(II27149), .A(g19893) );
  INV_X1 NOT_7164( .ZN(g20608), .A(II27149) );
  INV_X1 NOT_7165( .ZN(II27152), .A(g20360) );
  INV_X1 NOT_7166( .ZN(g20609), .A(II27152) );
  INV_X1 NOT_7167( .ZN(II27155), .A(g20395) );
  INV_X1 NOT_7168( .ZN(g20610), .A(II27155) );
  INV_X1 NOT_7169( .ZN(II27158), .A(g20439) );
  INV_X1 NOT_7170( .ZN(g20611), .A(II27158) );
  INV_X1 NOT_7171( .ZN(II27161), .A(g20377) );
  INV_X1 NOT_7172( .ZN(g20612), .A(II27161) );
  INV_X1 NOT_7173( .ZN(II27164), .A(g20418) );
  INV_X1 NOT_7174( .ZN(g20613), .A(II27164) );
  INV_X1 NOT_7175( .ZN(II27167), .A(g20457) );
  INV_X1 NOT_7176( .ZN(g20614), .A(II27167) );
  INV_X1 NOT_7177( .ZN(II27170), .A(g20396) );
  INV_X1 NOT_7178( .ZN(g20615), .A(II27170) );
  INV_X1 NOT_7179( .ZN(II27173), .A(g20440) );
  INV_X1 NOT_7180( .ZN(g20616), .A(II27173) );
  INV_X1 NOT_7181( .ZN(II27176), .A(g20469) );
  INV_X1 NOT_7182( .ZN(g20617), .A(II27176) );
  INV_X1 NOT_7183( .ZN(II27179), .A(g20419) );
  INV_X1 NOT_7184( .ZN(g20618), .A(II27179) );
  INV_X1 NOT_7185( .ZN(II27182), .A(g20458) );
  INV_X1 NOT_7186( .ZN(g20619), .A(II27182) );
  INV_X1 NOT_7187( .ZN(II27185), .A(g20478) );
  INV_X1 NOT_7188( .ZN(g20620), .A(II27185) );
  INV_X1 NOT_7189( .ZN(II27188), .A(g20441) );
  INV_X1 NOT_7190( .ZN(g20621), .A(II27188) );
  INV_X1 NOT_7191( .ZN(II27191), .A(g20470) );
  INV_X1 NOT_7192( .ZN(g20622), .A(II27191) );
  INV_X1 NOT_7193( .ZN(II27194), .A(g20484) );
  INV_X1 NOT_7194( .ZN(g20623), .A(II27194) );
  INV_X1 NOT_7195( .ZN(II27197), .A(g20459) );
  INV_X1 NOT_7196( .ZN(g20624), .A(II27197) );
  INV_X1 NOT_7197( .ZN(II27200), .A(g20479) );
  INV_X1 NOT_7198( .ZN(g20625), .A(II27200) );
  INV_X1 NOT_7199( .ZN(II27203), .A(g20491) );
  INV_X1 NOT_7200( .ZN(g20626), .A(II27203) );
  INV_X1 NOT_7201( .ZN(II27206), .A(g20471) );
  INV_X1 NOT_7202( .ZN(g20627), .A(II27206) );
  INV_X1 NOT_7203( .ZN(II27209), .A(g20485) );
  INV_X1 NOT_7204( .ZN(g20628), .A(II27209) );
  INV_X1 NOT_7205( .ZN(II27212), .A(g20498) );
  INV_X1 NOT_7206( .ZN(g20629), .A(II27212) );
  INV_X1 NOT_7207( .ZN(II27215), .A(g19158) );
  INV_X1 NOT_7208( .ZN(g20630), .A(II27215) );
  INV_X1 NOT_7209( .ZN(II27218), .A(g19168) );
  INV_X1 NOT_7210( .ZN(g20631), .A(II27218) );
  INV_X1 NOT_7211( .ZN(II27221), .A(g19180) );
  INV_X1 NOT_7212( .ZN(g20632), .A(II27221) );
  INV_X1 NOT_7213( .ZN(II27225), .A(g19358) );
  INV_X1 NOT_7214( .ZN(g20634), .A(II27225) );
  INV_X1 NOT_7215( .ZN(II27228), .A(g19390) );
  INV_X1 NOT_7216( .ZN(g20637), .A(II27228) );
  INV_X1 NOT_7217( .ZN(II27232), .A(g19401) );
  INV_X1 NOT_7218( .ZN(g20641), .A(II27232) );
  INV_X1 NOT_7219( .ZN(II27235), .A(g19420) );
  INV_X1 NOT_7220( .ZN(g20644), .A(II27235) );
  INV_X1 NOT_7221( .ZN(II27240), .A(g19335) );
  INV_X1 NOT_7222( .ZN(g20649), .A(II27240) );
  INV_X1 NOT_7223( .ZN(II27243), .A(g19335) );
  INV_X1 NOT_7224( .ZN(g20652), .A(II27243) );
  INV_X1 NOT_7225( .ZN(II27246), .A(g19335) );
  INV_X1 NOT_7226( .ZN(g20655), .A(II27246) );
  INV_X1 NOT_7227( .ZN(II27250), .A(g19390) );
  INV_X1 NOT_7228( .ZN(g20659), .A(II27250) );
  INV_X1 NOT_7229( .ZN(II27253), .A(g19420) );
  INV_X1 NOT_7230( .ZN(g20662), .A(II27253) );
  INV_X1 NOT_7231( .ZN(II27257), .A(g19431) );
  INV_X1 NOT_7232( .ZN(g20666), .A(II27257) );
  INV_X1 NOT_7233( .ZN(II27260), .A(g19457) );
  INV_X1 NOT_7234( .ZN(g20669), .A(II27260) );
  INV_X1 NOT_7235( .ZN(II27264), .A(g19358) );
  INV_X1 NOT_7236( .ZN(g20673), .A(II27264) );
  INV_X1 NOT_7237( .ZN(II27267), .A(g19358) );
  INV_X1 NOT_7238( .ZN(g20676), .A(II27267) );
  INV_X1 NOT_7239( .ZN(II27270), .A(g19335) );
  INV_X1 NOT_7240( .ZN(g20679), .A(II27270) );
  INV_X1 NOT_7241( .ZN(II27275), .A(g19369) );
  INV_X1 NOT_7242( .ZN(g20684), .A(II27275) );
  INV_X1 NOT_7243( .ZN(II27278), .A(g19369) );
  INV_X1 NOT_7244( .ZN(g20687), .A(II27278) );
  INV_X1 NOT_7245( .ZN(II27281), .A(g19369) );
  INV_X1 NOT_7246( .ZN(g20690), .A(II27281) );
  INV_X1 NOT_7247( .ZN(II27285), .A(g19420) );
  INV_X1 NOT_7248( .ZN(g20694), .A(II27285) );
  INV_X1 NOT_7249( .ZN(II27288), .A(g19457) );
  INV_X1 NOT_7250( .ZN(g20697), .A(II27288) );
  INV_X1 NOT_7251( .ZN(II27293), .A(g19335) );
  INV_X1 NOT_7252( .ZN(g20704), .A(II27293) );
  INV_X1 NOT_7253( .ZN(II27297), .A(g19390) );
  INV_X1 NOT_7254( .ZN(g20708), .A(II27297) );
  INV_X1 NOT_7255( .ZN(II27300), .A(g19390) );
  INV_X1 NOT_7256( .ZN(g20711), .A(II27300) );
  INV_X1 NOT_7257( .ZN(II27303), .A(g19369) );
  INV_X1 NOT_7258( .ZN(g20714), .A(II27303) );
  INV_X1 NOT_7259( .ZN(II27308), .A(g19401) );
  INV_X1 NOT_7260( .ZN(g20719), .A(II27308) );
  INV_X1 NOT_7261( .ZN(II27311), .A(g19401) );
  INV_X1 NOT_7262( .ZN(g20722), .A(II27311) );
  INV_X1 NOT_7263( .ZN(II27314), .A(g19401) );
  INV_X1 NOT_7264( .ZN(g20725), .A(II27314) );
  INV_X1 NOT_7265( .ZN(II27318), .A(g19457) );
  INV_X1 NOT_7266( .ZN(g20729), .A(II27318) );
  INV_X1 NOT_7267( .ZN(II27321), .A(g19335) );
  INV_X1 NOT_7268( .ZN(g20732), .A(II27321) );
  INV_X1 NOT_7269( .ZN(II27324), .A(g19358) );
  INV_X1 NOT_7270( .ZN(g20735), .A(II27324) );
  INV_X1 NOT_7271( .ZN(II27328), .A(g19369) );
  INV_X1 NOT_7272( .ZN(g20739), .A(II27328) );
  INV_X1 NOT_7273( .ZN(II27332), .A(g19420) );
  INV_X1 NOT_7274( .ZN(g20743), .A(II27332) );
  INV_X1 NOT_7275( .ZN(II27335), .A(g19420) );
  INV_X1 NOT_7276( .ZN(g20746), .A(II27335) );
  INV_X1 NOT_7277( .ZN(II27338), .A(g19401) );
  INV_X1 NOT_7278( .ZN(g20749), .A(II27338) );
  INV_X1 NOT_7279( .ZN(II27343), .A(g19431) );
  INV_X1 NOT_7280( .ZN(g20754), .A(II27343) );
  INV_X1 NOT_7281( .ZN(II27346), .A(g19431) );
  INV_X1 NOT_7282( .ZN(g20757), .A(II27346) );
  INV_X1 NOT_7283( .ZN(II27349), .A(g19431) );
  INV_X1 NOT_7284( .ZN(g20760), .A(II27349) );
  INV_X1 NOT_7285( .ZN(II27352), .A(g19358) );
  INV_X1 NOT_7286( .ZN(g20763), .A(II27352) );
  INV_X1 NOT_7287( .ZN(II27355), .A(g19335) );
  INV_X1 NOT_7288( .ZN(g20766), .A(II27355) );
  INV_X1 NOT_7289( .ZN(II27358), .A(g19369) );
  INV_X1 NOT_7290( .ZN(g20769), .A(II27358) );
  INV_X1 NOT_7291( .ZN(II27361), .A(g19390) );
  INV_X1 NOT_7292( .ZN(g20772), .A(II27361) );
  INV_X1 NOT_7293( .ZN(II27365), .A(g19401) );
  INV_X4 NOT_7294( .ZN(g20776), .A(II27365) );
  INV_X4 NOT_7295( .ZN(II27369), .A(g19457) );
  INV_X4 NOT_7296( .ZN(g20780), .A(II27369) );
  INV_X1 NOT_7297( .ZN(II27372), .A(g19457) );
  INV_X1 NOT_7298( .ZN(g20783), .A(II27372) );
  INV_X1 NOT_7299( .ZN(II27375), .A(g19431) );
  INV_X1 NOT_7300( .ZN(g20786), .A(II27375) );
  INV_X1 NOT_7301( .ZN(II27379), .A(g19358) );
  INV_X1 NOT_7302( .ZN(g20790), .A(II27379) );
  INV_X1 NOT_7303( .ZN(II27382), .A(g19390) );
  INV_X1 NOT_7304( .ZN(g20793), .A(II27382) );
  INV_X1 NOT_7305( .ZN(II27385), .A(g19369) );
  INV_X1 NOT_7306( .ZN(g20796), .A(II27385) );
  INV_X1 NOT_7307( .ZN(II27388), .A(g19401) );
  INV_X1 NOT_7308( .ZN(g20799), .A(II27388) );
  INV_X1 NOT_7309( .ZN(II27391), .A(g19420) );
  INV_X1 NOT_7310( .ZN(g20802), .A(II27391) );
  INV_X1 NOT_7311( .ZN(II27395), .A(g19431) );
  INV_X1 NOT_7312( .ZN(g20806), .A(II27395) );
  INV_X1 NOT_7313( .ZN(II27399), .A(g19390) );
  INV_X1 NOT_7314( .ZN(g20810), .A(II27399) );
  INV_X1 NOT_7315( .ZN(II27402), .A(g19420) );
  INV_X1 NOT_7316( .ZN(g20813), .A(II27402) );
  INV_X1 NOT_7317( .ZN(II27405), .A(g19401) );
  INV_X1 NOT_7318( .ZN(g20816), .A(II27405) );
  INV_X1 NOT_7319( .ZN(II27408), .A(g19431) );
  INV_X1 NOT_7320( .ZN(g20819), .A(II27408) );
  INV_X1 NOT_7321( .ZN(II27411), .A(g19457) );
  INV_X1 NOT_7322( .ZN(g20822), .A(II27411) );
  INV_X1 NOT_7323( .ZN(II27416), .A(g19420) );
  INV_X1 NOT_7324( .ZN(g20827), .A(II27416) );
  INV_X1 NOT_7325( .ZN(II27419), .A(g19457) );
  INV_X1 NOT_7326( .ZN(g20830), .A(II27419) );
  INV_X1 NOT_7327( .ZN(II27422), .A(g19431) );
  INV_X1 NOT_7328( .ZN(g20833), .A(II27422) );
  INV_X1 NOT_7329( .ZN(II27426), .A(g19457) );
  INV_X1 NOT_7330( .ZN(g20837), .A(II27426) );
  INV_X1 NOT_7331( .ZN(g20842), .A(g19441) );
  INV_X1 NOT_7332( .ZN(g20850), .A(g19468) );
  INV_X1 NOT_7333( .ZN(g20858), .A(g19491) );
  INV_X1 NOT_7334( .ZN(g20866), .A(g19512) );
  INV_X1 NOT_7335( .ZN(g20885), .A(g19865) );
  INV_X1 NOT_7336( .ZN(g20904), .A(g19896) );
  INV_X1 NOT_7337( .ZN(g20928), .A(g19921) );
  INV_X1 NOT_7338( .ZN(II27488), .A(g20310) );
  INV_X1 NOT_7339( .ZN(g20942), .A(II27488) );
  INV_X1 NOT_7340( .ZN(II27491), .A(g20314) );
  INV_X1 NOT_7341( .ZN(g20943), .A(II27491) );
  INV_X1 NOT_7342( .ZN(g20956), .A(g19936) );
  INV_X1 NOT_7343( .ZN(II27516), .A(g20333) );
  INV_X1 NOT_7344( .ZN(g20971), .A(II27516) );
  INV_X1 NOT_7345( .ZN(II27531), .A(g20343) );
  INV_X1 NOT_7346( .ZN(g20984), .A(II27531) );
  INV_X1 NOT_7347( .ZN(II27534), .A(g20083) );
  INV_X1 NOT_7348( .ZN(g20985), .A(II27534) );
  INV_X1 NOT_7349( .ZN(II27537), .A(g19957) );
  INV_X1 NOT_7350( .ZN(g20986), .A(II27537) );
  INV_X1 NOT_7351( .ZN(II27549), .A(g20353) );
  INV_X1 NOT_7352( .ZN(g20998), .A(II27549) );
  INV_X1 NOT_7353( .ZN(II27565), .A(g19987) );
  INV_X1 NOT_7354( .ZN(g21012), .A(II27565) );
  INV_X1 NOT_7355( .ZN(II27577), .A(g20375) );
  INV_X1 NOT_7356( .ZN(g21024), .A(II27577) );
  INV_X1 NOT_7357( .ZN(II27585), .A(g20376) );
  INV_X1 NOT_7358( .ZN(g21030), .A(II27585) );
  INV_X1 NOT_7359( .ZN(II27593), .A(g20025) );
  INV_X1 NOT_7360( .ZN(g21036), .A(II27593) );
  INV_X1 NOT_7361( .ZN(g21050), .A(g20513) );
  INV_X1 NOT_7362( .ZN(II27614), .A(g20067) );
  INV_X1 NOT_7363( .ZN(g21057), .A(II27614) );
  INV_X1 NOT_7364( .ZN(II27621), .A(g20417) );
  INV_X1 NOT_7365( .ZN(g21064), .A(II27621) );
  INV_X1 NOT_7366( .ZN(g21066), .A(g20519) );
  INV_X1 NOT_7367( .ZN(g21069), .A(g20531) );
  INV_X1 NOT_7368( .ZN(g21076), .A(g20539) );
  INV_X1 NOT_7369( .ZN(g21079), .A(g20550) );
  INV_X1 NOT_7370( .ZN(II27646), .A(g20507) );
  INV_X1 NOT_7371( .ZN(g21087), .A(II27646) );
  INV_X1 NOT_7372( .ZN(g21090), .A(g19064) );
  INV_X1 NOT_7373( .ZN(g21093), .A(g19075) );
  INV_X1 NOT_7374( .ZN(II27658), .A(g20526) );
  INV_X1 NOT_7375( .ZN(g21099), .A(II27658) );
  INV_X1 NOT_7376( .ZN(g21102), .A(g19081) );
  INV_X1 NOT_7377( .ZN(II27667), .A(g20507) );
  INV_X1 NOT_7378( .ZN(g21108), .A(II27667) );
  INV_X1 NOT_7379( .ZN(II27672), .A(g20545) );
  INV_X1 NOT_7380( .ZN(g21113), .A(II27672) );
  INV_X1 NOT_7381( .ZN(II27684), .A(g20526) );
  INV_X1 NOT_7382( .ZN(g21125), .A(II27684) );
  INV_X1 NOT_7383( .ZN(II27689), .A(g19070) );
  INV_X1 NOT_7384( .ZN(g21130), .A(II27689) );
  INV_X1 NOT_7385( .ZN(II27705), .A(g20545) );
  INV_X1 NOT_7386( .ZN(g21144), .A(II27705) );
  INV_X1 NOT_7387( .ZN(II27727), .A(g19070) );
  INV_X1 NOT_7388( .ZN(g21164), .A(II27727) );
  INV_X1 NOT_7389( .ZN(II27749), .A(g19954) );
  INV_X1 NOT_7390( .ZN(g21184), .A(II27749) );
  INV_X1 NOT_7391( .ZN(g21187), .A(g19113) );
  INV_X1 NOT_7392( .ZN(II27766), .A(g19984) );
  INV_X1 NOT_7393( .ZN(g21199), .A(II27766) );
  INV_X1 NOT_7394( .ZN(g21202), .A(g19118) );
  INV_X1 NOT_7395( .ZN(II27779), .A(g20022) );
  INV_X1 NOT_7396( .ZN(g21214), .A(II27779) );
  INV_X1 NOT_7397( .ZN(g21217), .A(g19125) );
  INV_X1 NOT_7398( .ZN(II27785), .A(g20064) );
  INV_X1 NOT_7399( .ZN(g21222), .A(II27785) );
  INV_X1 NOT_7400( .ZN(g21225), .A(g19132) );
  INV_X1 NOT_7401( .ZN(g21241), .A(g19945) );
  INV_X1 NOT_7402( .ZN(g21249), .A(g19972) );
  INV_X1 NOT_7403( .ZN(g21258), .A(g20002) );
  INV_X1 NOT_7404( .ZN(g21266), .A(g20040) );
  INV_X1 NOT_7405( .ZN(II27822), .A(g19865) );
  INV_X1 NOT_7406( .ZN(g21271), .A(II27822) );
  INV_X1 NOT_7407( .ZN(II27827), .A(g19896) );
  INV_X1 NOT_7408( .ZN(g21278), .A(II27827) );
  INV_X1 NOT_7409( .ZN(II27832), .A(g19921) );
  INV_X1 NOT_7410( .ZN(g21285), .A(II27832) );
  INV_X1 NOT_7411( .ZN(II27838), .A(g19936) );
  INV_X1 NOT_7412( .ZN(g21293), .A(II27838) );
  INV_X1 NOT_7413( .ZN(II27868), .A(g19144) );
  INV_X1 NOT_7414( .ZN(g21327), .A(II27868) );
  INV_X1 NOT_7415( .ZN(II27897), .A(g19149) );
  INV_X1 NOT_7416( .ZN(g21358), .A(II27897) );
  INV_X1 NOT_7417( .ZN(II27900), .A(g19096) );
  INV_X1 NOT_7418( .ZN(g21359), .A(II27900) );
  INV_X1 NOT_7419( .ZN(II27917), .A(g19153) );
  INV_X1 NOT_7420( .ZN(g21376), .A(II27917) );
  INV_X1 NOT_7421( .ZN(II27920), .A(g19154) );
  INV_X1 NOT_7422( .ZN(g21377), .A(II27920) );
  INV_X1 NOT_7423( .ZN(II27927), .A(g19957) );
  INV_X1 NOT_7424( .ZN(g21382), .A(II27927) );
  INV_X1 NOT_7425( .ZN(II27942), .A(g19157) );
  INV_X1 NOT_7426( .ZN(g21399), .A(II27942) );
  INV_X1 NOT_7427( .ZN(g21400), .A(g19918) );
  INV_X1 NOT_7428( .ZN(II27949), .A(g19957) );
  INV_X1 NOT_7429( .ZN(g21404), .A(II27949) );
  INV_X1 NOT_7430( .ZN(II27958), .A(g19987) );
  INV_X1 NOT_7431( .ZN(g21415), .A(II27958) );
  INV_X1 NOT_7432( .ZN(II27969), .A(g19162) );
  INV_X1 NOT_7433( .ZN(g21426), .A(II27969) );
  INV_X1 NOT_7434( .ZN(II27972), .A(g19163) );
  INV_X1 NOT_7435( .ZN(g21427), .A(II27972) );
  INV_X1 NOT_7436( .ZN(II27976), .A(g19957) );
  INV_X1 NOT_7437( .ZN(g21429), .A(II27976) );
  INV_X1 NOT_7438( .ZN(II27984), .A(g19987) );
  INV_X1 NOT_7439( .ZN(g21441), .A(II27984) );
  INV_X1 NOT_7440( .ZN(II27992), .A(g20025) );
  INV_X1 NOT_7441( .ZN(g21449), .A(II27992) );
  INV_X1 NOT_7442( .ZN(II28000), .A(g19167) );
  INV_X1 NOT_7443( .ZN(g21457), .A(II28000) );
  INV_X1 NOT_7444( .ZN(II28003), .A(g19957) );
  INV_X1 NOT_7445( .ZN(g21458), .A(II28003) );
  INV_X1 NOT_7446( .ZN(g21461), .A(g19957) );
  INV_X1 NOT_7447( .ZN(II28009), .A(g20473) );
  INV_X1 NOT_7448( .ZN(g21473), .A(II28009) );
  INV_X1 NOT_7449( .ZN(II28013), .A(g19987) );
  INV_X1 NOT_7450( .ZN(g21477), .A(II28013) );
  INV_X1 NOT_7451( .ZN(II28019), .A(g20025) );
  INV_X1 NOT_7452( .ZN(g21483), .A(II28019) );
  INV_X1 NOT_7453( .ZN(II28027), .A(g20067) );
  INV_X1 NOT_7454( .ZN(g21491), .A(II28027) );
  INV_X1 NOT_7455( .ZN(II28031), .A(g19172) );
  INV_X1 NOT_7456( .ZN(g21495), .A(II28031) );
  INV_X1 NOT_7457( .ZN(II28034), .A(g19173) );
  INV_X1 NOT_7458( .ZN(g21496), .A(II28034) );
  INV_X1 NOT_7459( .ZN(II28038), .A(g19957) );
  INV_X1 NOT_7460( .ZN(g21498), .A(II28038) );
  INV_X1 NOT_7461( .ZN(II28043), .A(g19987) );
  INV_X1 NOT_7462( .ZN(g21505), .A(II28043) );
  INV_X1 NOT_7463( .ZN(g21508), .A(g19987) );
  INV_X1 NOT_7464( .ZN(II28047), .A(g20481) );
  INV_X1 NOT_7465( .ZN(g21514), .A(II28047) );
  INV_X1 NOT_7466( .ZN(II28051), .A(g20025) );
  INV_X1 NOT_7467( .ZN(g21518), .A(II28051) );
  INV_X1 NOT_7468( .ZN(II28057), .A(g20067) );
  INV_X1 NOT_7469( .ZN(g21524), .A(II28057) );
  INV_X4 NOT_7470( .ZN(II28061), .A(g19178) );
  INV_X4 NOT_7471( .ZN(g21528), .A(II28061) );
  INV_X4 NOT_7472( .ZN(g21529), .A(g19272) );
  INV_X1 NOT_7473( .ZN(II28065), .A(g19957) );
  INV_X1 NOT_7474( .ZN(g21530), .A(II28065) );
  INV_X1 NOT_7475( .ZN(II28072), .A(g19987) );
  INV_X1 NOT_7476( .ZN(g21537), .A(II28072) );
  INV_X1 NOT_7477( .ZN(II28076), .A(g20025) );
  INV_X1 NOT_7478( .ZN(g21541), .A(II28076) );
  INV_X1 NOT_7479( .ZN(g21544), .A(g20025) );
  INV_X1 NOT_7480( .ZN(II28080), .A(g20487) );
  INV_X1 NOT_7481( .ZN(g21550), .A(II28080) );
  INV_X1 NOT_7482( .ZN(II28084), .A(g20067) );
  INV_X1 NOT_7483( .ZN(g21554), .A(II28084) );
  INV_X1 NOT_7484( .ZN(II28087), .A(g19184) );
  INV_X1 NOT_7485( .ZN(g21557), .A(II28087) );
  INV_X1 NOT_7486( .ZN(II28090), .A(g20008) );
  INV_X1 NOT_7487( .ZN(g21558), .A(II28090) );
  INV_X1 NOT_7488( .ZN(II28093), .A(g19957) );
  INV_X1 NOT_7489( .ZN(g21561), .A(II28093) );
  INV_X1 NOT_7490( .ZN(g21565), .A(g19291) );
  INV_X1 NOT_7491( .ZN(II28100), .A(g19987) );
  INV_X1 NOT_7492( .ZN(g21566), .A(II28100) );
  INV_X1 NOT_7493( .ZN(II28107), .A(g20025) );
  INV_X1 NOT_7494( .ZN(g21573), .A(II28107) );
  INV_X1 NOT_7495( .ZN(II28111), .A(g20067) );
  INV_X1 NOT_7496( .ZN(g21577), .A(II28111) );
  INV_X1 NOT_7497( .ZN(g21580), .A(g20067) );
  INV_X1 NOT_7498( .ZN(II28115), .A(g20493) );
  INV_X1 NOT_7499( .ZN(g21586), .A(II28115) );
  INV_X1 NOT_7500( .ZN(II28119), .A(g19957) );
  INV_X1 NOT_7501( .ZN(g21590), .A(II28119) );
  INV_X1 NOT_7502( .ZN(II28123), .A(g19987) );
  INV_X1 NOT_7503( .ZN(g21594), .A(II28123) );
  INV_X1 NOT_7504( .ZN(g21598), .A(g19309) );
  INV_X1 NOT_7505( .ZN(II28130), .A(g20025) );
  INV_X1 NOT_7506( .ZN(g21599), .A(II28130) );
  INV_X1 NOT_7507( .ZN(II28137), .A(g20067) );
  INV_X1 NOT_7508( .ZN(g21606), .A(II28137) );
  INV_X1 NOT_7509( .ZN(II28143), .A(g19957) );
  INV_X1 NOT_7510( .ZN(g21612), .A(II28143) );
  INV_X1 NOT_7511( .ZN(II28148), .A(g19987) );
  INV_X1 NOT_7512( .ZN(g21619), .A(II28148) );
  INV_X1 NOT_7513( .ZN(II28152), .A(g20025) );
  INV_X1 NOT_7514( .ZN(g21623), .A(II28152) );
  INV_X1 NOT_7515( .ZN(g21627), .A(g19330) );
  INV_X1 NOT_7516( .ZN(II28159), .A(g20067) );
  INV_X1 NOT_7517( .ZN(g21628), .A(II28159) );
  INV_X1 NOT_7518( .ZN(II28169), .A(g19987) );
  INV_X1 NOT_7519( .ZN(g21640), .A(II28169) );
  INV_X1 NOT_7520( .ZN(II28174), .A(g20025) );
  INV_X1 NOT_7521( .ZN(g21647), .A(II28174) );
  INV_X1 NOT_7522( .ZN(II28178), .A(g20067) );
  INV_X1 NOT_7523( .ZN(g21651), .A(II28178) );
  INV_X1 NOT_7524( .ZN(II28184), .A(g19103) );
  INV_X1 NOT_7525( .ZN(g21655), .A(II28184) );
  INV_X1 NOT_7526( .ZN(g21661), .A(g19091) );
  INV_X1 NOT_7527( .ZN(II28201), .A(g20025) );
  INV_X1 NOT_7528( .ZN(g21671), .A(II28201) );
  INV_X1 NOT_7529( .ZN(II28206), .A(g20067) );
  INV_X1 NOT_7530( .ZN(g21678), .A(II28206) );
  INV_X1 NOT_7531( .ZN(II28210), .A(g20537) );
  INV_X1 NOT_7532( .ZN(g21682), .A(II28210) );
  INV_X1 NOT_7533( .ZN(g21690), .A(g19098) );
  INV_X1 NOT_7534( .ZN(II28229), .A(g20067) );
  INV_X1 NOT_7535( .ZN(g21700), .A(II28229) );
  INV_X1 NOT_7536( .ZN(II28235), .A(g20153) );
  INV_X1 NOT_7537( .ZN(g21708), .A(II28235) );
  INV_X1 NOT_7538( .ZN(g21716), .A(g19894) );
  INV_X1 NOT_7539( .ZN(g21726), .A(g19105) );
  INV_X1 NOT_7540( .ZN(g21742), .A(g19919) );
  INV_X1 NOT_7541( .ZN(g21752), .A(g19110) );
  INV_X1 NOT_7542( .ZN(g21766), .A(g19934) );
  INV_X1 NOT_7543( .ZN(g21782), .A(g19951) );
  INV_X1 NOT_7544( .ZN(II28314), .A(g19152) );
  INV_X1 NOT_7545( .ZN(g21795), .A(II28314) );
  INV_X1 NOT_7546( .ZN(II28357), .A(g20497) );
  INV_X1 NOT_7547( .ZN(g21824), .A(II28357) );
  INV_X1 NOT_7548( .ZN(II28360), .A(g20163) );
  INV_X1 NOT_7549( .ZN(g21825), .A(II28360) );
  INV_X1 NOT_7550( .ZN(g21861), .A(g19657) );
  INV_X1 NOT_7551( .ZN(g21867), .A(g19705) );
  INV_X1 NOT_7552( .ZN(g21872), .A(g19749) );
  INV_X1 NOT_7553( .ZN(g21876), .A(g19792) );
  INV_X1 NOT_7554( .ZN(g21883), .A(g19890) );
  INV_X1 NOT_7555( .ZN(g21886), .A(g19915) );
  INV_X1 NOT_7556( .ZN(g21895), .A(g19945) );
  INV_X1 NOT_7557( .ZN(g21902), .A(g19978) );
  INV_X1 NOT_7558( .ZN(g21907), .A(g19972) );
  INV_X1 NOT_7559( .ZN(II28432), .A(g19335) );
  INV_X1 NOT_7560( .ZN(g21914), .A(II28432) );
  INV_X1 NOT_7561( .ZN(II28435), .A(g19358) );
  INV_X1 NOT_7562( .ZN(g21917), .A(II28435) );
  INV_X1 NOT_7563( .ZN(g21921), .A(g20002) );
  INV_X1 NOT_7564( .ZN(g21927), .A(g20045) );
  INV_X1 NOT_7565( .ZN(II28443), .A(g19358) );
  INV_X1 NOT_7566( .ZN(g21928), .A(II28443) );
  INV_X1 NOT_7567( .ZN(II28447), .A(g19369) );
  INV_X1 NOT_7568( .ZN(g21932), .A(II28447) );
  INV_X1 NOT_7569( .ZN(II28450), .A(g19390) );
  INV_X1 NOT_7570( .ZN(g21935), .A(II28450) );
  INV_X1 NOT_7571( .ZN(g21939), .A(g20040) );
  INV_X1 NOT_7572( .ZN(II28455), .A(g20943) );
  INV_X1 NOT_7573( .ZN(g21943), .A(II28455) );
  INV_X1 NOT_7574( .ZN(II28458), .A(g20971) );
  INV_X1 NOT_7575( .ZN(g21944), .A(II28458) );
  INV_X1 NOT_7576( .ZN(II28461), .A(g20998) );
  INV_X1 NOT_7577( .ZN(g21945), .A(II28461) );
  INV_X1 NOT_7578( .ZN(II28464), .A(g21024) );
  INV_X1 NOT_7579( .ZN(g21946), .A(II28464) );
  INV_X1 NOT_7580( .ZN(II28467), .A(g20942) );
  INV_X1 NOT_7581( .ZN(g21947), .A(II28467) );
  INV_X1 NOT_7582( .ZN(II28470), .A(g20984) );
  INV_X1 NOT_7583( .ZN(g21948), .A(II28470) );
  INV_X1 NOT_7584( .ZN(II28473), .A(g21030) );
  INV_X1 NOT_7585( .ZN(g21949), .A(II28473) );
  INV_X1 NOT_7586( .ZN(II28476), .A(g21064) );
  INV_X1 NOT_7587( .ZN(g21950), .A(II28476) );
  INV_X1 NOT_7588( .ZN(II28479), .A(g21795) );
  INV_X1 NOT_7589( .ZN(g21951), .A(II28479) );
  INV_X1 NOT_7590( .ZN(II28482), .A(g21376) );
  INV_X1 NOT_7591( .ZN(g21952), .A(II28482) );
  INV_X1 NOT_7592( .ZN(II28485), .A(g21426) );
  INV_X1 NOT_7593( .ZN(g21953), .A(II28485) );
  INV_X1 NOT_7594( .ZN(II28488), .A(g21495) );
  INV_X1 NOT_7595( .ZN(g21954), .A(II28488) );
  INV_X1 NOT_7596( .ZN(II28491), .A(g21327) );
  INV_X1 NOT_7597( .ZN(g21955), .A(II28491) );
  INV_X1 NOT_7598( .ZN(II28494), .A(g21358) );
  INV_X1 NOT_7599( .ZN(g21956), .A(II28494) );
  INV_X1 NOT_7600( .ZN(II28497), .A(g21399) );
  INV_X1 NOT_7601( .ZN(g21957), .A(II28497) );
  INV_X1 NOT_7602( .ZN(II28500), .A(g21457) );
  INV_X1 NOT_7603( .ZN(g21958), .A(II28500) );
  INV_X1 NOT_7604( .ZN(II28503), .A(g21528) );
  INV_X1 NOT_7605( .ZN(g21959), .A(II28503) );
  INV_X1 NOT_7606( .ZN(II28506), .A(g21377) );
  INV_X1 NOT_7607( .ZN(g21960), .A(II28506) );
  INV_X1 NOT_7608( .ZN(II28509), .A(g21427) );
  INV_X1 NOT_7609( .ZN(g21961), .A(II28509) );
  INV_X1 NOT_7610( .ZN(II28512), .A(g21496) );
  INV_X1 NOT_7611( .ZN(g21962), .A(II28512) );
  INV_X1 NOT_7612( .ZN(II28515), .A(g21557) );
  INV_X1 NOT_7613( .ZN(g21963), .A(II28515) );
  INV_X1 NOT_7614( .ZN(II28518), .A(g20985) );
  INV_X1 NOT_7615( .ZN(g21964), .A(II28518) );
  INV_X1 NOT_7616( .ZN(II28521), .A(g21824) );
  INV_X1 NOT_7617( .ZN(g21965), .A(II28521) );
  INV_X1 NOT_7618( .ZN(II28524), .A(g21359) );
  INV_X1 NOT_7619( .ZN(g21966), .A(II28524) );
  INV_X1 NOT_7620( .ZN(II28527), .A(g21407) );
  INV_X1 NOT_7621( .ZN(g21967), .A(II28527) );
  INV_X1 NOT_7622( .ZN(II28541), .A(g21467) );
  INV_X1 NOT_7623( .ZN(g21982), .A(II28541) );
  INV_X1 NOT_7624( .ZN(II28550), .A(g21432) );
  INV_X1 NOT_7625( .ZN(g21995), .A(II28550) );
  INV_X1 NOT_7626( .ZN(II28557), .A(g21407) );
  INV_X1 NOT_7627( .ZN(g22003), .A(II28557) );
  INV_X1 NOT_7628( .ZN(II28564), .A(g21385) );
  INV_X1 NOT_7629( .ZN(g22014), .A(II28564) );
  INV_X1 NOT_7630( .ZN(II28628), .A(g21842) );
  INV_X1 NOT_7631( .ZN(g22082), .A(II28628) );
  INV_X1 NOT_7632( .ZN(II28649), .A(g21843) );
  INV_X1 NOT_7633( .ZN(g22107), .A(II28649) );
  INV_X1 NOT_7634( .ZN(II28671), .A(g21845) );
  INV_X1 NOT_7635( .ZN(g22133), .A(II28671) );
  INV_X1 NOT_7636( .ZN(II28693), .A(g21847) );
  INV_X1 NOT_7637( .ZN(g22156), .A(II28693) );
  INV_X1 NOT_7638( .ZN(II28712), .A(g21851) );
  INV_X1 NOT_7639( .ZN(g22176), .A(II28712) );
  INV_X1 NOT_7640( .ZN(g22212), .A(g21914) );
  INV_X1 NOT_7641( .ZN(g22213), .A(g21917) );
  INV_X4 NOT_7642( .ZN(g22217), .A(g21928) );
  INV_X4 NOT_7643( .ZN(II28781), .A(g21331) );
  INV_X4 NOT_7644( .ZN(g22219), .A(II28781) );
  INV_X1 NOT_7645( .ZN(g22221), .A(g21932) );
  INV_X1 NOT_7646( .ZN(g22222), .A(g21935) );
  INV_X1 NOT_7647( .ZN(II28789), .A(g21878) );
  INV_X1 NOT_7648( .ZN(g22225), .A(II28789) );
  INV_X1 NOT_7649( .ZN(II28792), .A(g21880) );
  INV_X1 NOT_7650( .ZN(g22226), .A(II28792) );
  INV_X1 NOT_7651( .ZN(g22230), .A(g20634) );
  INV_X1 NOT_7652( .ZN(II28800), .A(g21316) );
  INV_X1 NOT_7653( .ZN(g22232), .A(II28800) );
  INV_X1 NOT_7654( .ZN(g22233), .A(g20637) );
  INV_X1 NOT_7655( .ZN(g22236), .A(g20641) );
  INV_X1 NOT_7656( .ZN(g22237), .A(g20644) );
  INV_X1 NOT_7657( .ZN(g22239), .A(g20649) );
  INV_X1 NOT_7658( .ZN(g22240), .A(g20652) );
  INV_X1 NOT_7659( .ZN(g22241), .A(g20655) );
  INV_X1 NOT_7660( .ZN(II28813), .A(g21502) );
  INV_X1 NOT_7661( .ZN(g22243), .A(II28813) );
  INV_X1 NOT_7662( .ZN(g22246), .A(g20659) );
  INV_X1 NOT_7663( .ZN(g22248), .A(g20662) );
  INV_X1 NOT_7664( .ZN(g22251), .A(g20666) );
  INV_X1 NOT_7665( .ZN(g22252), .A(g20669) );
  INV_X1 NOT_7666( .ZN(II28825), .A(g21882) );
  INV_X1 NOT_7667( .ZN(g22253), .A(II28825) );
  INV_X1 NOT_7668( .ZN(g22256), .A(g20673) );
  INV_X1 NOT_7669( .ZN(g22257), .A(g20676) );
  INV_X1 NOT_7670( .ZN(g22258), .A(g20679) );
  INV_X1 NOT_7671( .ZN(II28833), .A(g21470) );
  INV_X1 NOT_7672( .ZN(g22259), .A(II28833) );
  INV_X1 NOT_7673( .ZN(g22260), .A(g20684) );
  INV_X1 NOT_7674( .ZN(g22261), .A(g20687) );
  INV_X1 NOT_7675( .ZN(g22262), .A(g20690) );
  INV_X1 NOT_7676( .ZN(g22266), .A(g20694) );
  INV_X1 NOT_7677( .ZN(g22268), .A(g20697) );
  INV_X1 NOT_7678( .ZN(g22271), .A(g20704) );
  INV_X1 NOT_7679( .ZN(g22274), .A(g20708) );
  INV_X1 NOT_7680( .ZN(g22275), .A(g20711) );
  INV_X1 NOT_7681( .ZN(g22276), .A(g20714) );
  INV_X1 NOT_7682( .ZN(g22277), .A(g20719) );
  INV_X1 NOT_7683( .ZN(g22278), .A(g20722) );
  INV_X1 NOT_7684( .ZN(g22279), .A(g20725) );
  INV_X1 NOT_7685( .ZN(g22283), .A(g20729) );
  INV_X1 NOT_7686( .ZN(g22286), .A(g20732) );
  INV_X1 NOT_7687( .ZN(g22287), .A(g20735) );
  INV_X1 NOT_7688( .ZN(g22290), .A(g20739) );
  INV_X1 NOT_7689( .ZN(g22293), .A(g20743) );
  INV_X1 NOT_7690( .ZN(g22294), .A(g20746) );
  INV_X1 NOT_7691( .ZN(g22295), .A(g20749) );
  INV_X1 NOT_7692( .ZN(g22296), .A(g20754) );
  INV_X1 NOT_7693( .ZN(g22297), .A(g20757) );
  INV_X1 NOT_7694( .ZN(g22298), .A(g20760) );
  INV_X1 NOT_7695( .ZN(II28876), .A(g21238) );
  INV_X1 NOT_7696( .ZN(g22300), .A(II28876) );
  INV_X1 NOT_7697( .ZN(g22303), .A(g20763) );
  INV_X1 NOT_7698( .ZN(g22304), .A(g20766) );
  INV_X1 NOT_7699( .ZN(g22306), .A(g20769) );
  INV_X1 NOT_7700( .ZN(g22307), .A(g20772) );
  INV_X1 NOT_7701( .ZN(g22310), .A(g20776) );
  INV_X1 NOT_7702( .ZN(g22313), .A(g20780) );
  INV_X1 NOT_7703( .ZN(g22314), .A(g20783) );
  INV_X1 NOT_7704( .ZN(g22315), .A(g20786) );
  INV_X1 NOT_7705( .ZN(g22316), .A(g21149) );
  INV_X1 NOT_7706( .ZN(g22318), .A(g20790) );
  INV_X1 NOT_7707( .ZN(g22319), .A(g21228) );
  INV_X1 NOT_7708( .ZN(II28896), .A(g21246) );
  INV_X1 NOT_7709( .ZN(g22328), .A(II28896) );
  INV_X1 NOT_7710( .ZN(g22331), .A(g20793) );
  INV_X1 NOT_7711( .ZN(g22332), .A(g20796) );
  INV_X1 NOT_7712( .ZN(g22334), .A(g20799) );
  INV_X1 NOT_7713( .ZN(g22335), .A(g20802) );
  INV_X1 NOT_7714( .ZN(g22338), .A(g20806) );
  INV_X1 NOT_7715( .ZN(g22341), .A(g21169) );
  INV_X1 NOT_7716( .ZN(g22343), .A(g20810) );
  INV_X1 NOT_7717( .ZN(g22344), .A(g21233) );
  INV_X1 NOT_7718( .ZN(II28913), .A(g21255) );
  INV_X1 NOT_7719( .ZN(g22353), .A(II28913) );
  INV_X1 NOT_7720( .ZN(g22356), .A(g20813) );
  INV_X1 NOT_7721( .ZN(g22357), .A(g20816) );
  INV_X1 NOT_7722( .ZN(g22359), .A(g20819) );
  INV_X1 NOT_7723( .ZN(g22360), .A(g20822) );
  INV_X1 NOT_7724( .ZN(g22364), .A(g21189) );
  INV_X1 NOT_7725( .ZN(g22366), .A(g20827) );
  INV_X1 NOT_7726( .ZN(g22367), .A(g21242) );
  INV_X1 NOT_7727( .ZN(II28928), .A(g21263) );
  INV_X1 NOT_7728( .ZN(g22376), .A(II28928) );
  INV_X1 NOT_7729( .ZN(g22379), .A(g20830) );
  INV_X1 NOT_7730( .ZN(g22380), .A(g20833) );
  INV_X1 NOT_7731( .ZN(g22384), .A(g21204) );
  INV_X1 NOT_7732( .ZN(g22386), .A(g20837) );
  INV_X1 NOT_7733( .ZN(g22387), .A(g21250) );
  INV_X1 NOT_7734( .ZN(g22401), .A(g21533) );
  INV_X1 NOT_7735( .ZN(g22402), .A(g21569) );
  INV_X1 NOT_7736( .ZN(g22403), .A(g21602) );
  INV_X1 NOT_7737( .ZN(g22404), .A(g21631) );
  INV_X1 NOT_7738( .ZN(II28949), .A(g21685) );
  INV_X1 NOT_7739( .ZN(g22405), .A(II28949) );
  INV_X1 NOT_7740( .ZN(g22408), .A(g20986) );
  INV_X1 NOT_7741( .ZN(II28953), .A(g21659) );
  INV_X1 NOT_7742( .ZN(g22409), .A(II28953) );
  INV_X1 NOT_7743( .ZN(II28956), .A(g21714) );
  INV_X1 NOT_7744( .ZN(g22412), .A(II28956) );
  INV_X1 NOT_7745( .ZN(II28959), .A(g21636) );
  INV_X1 NOT_7746( .ZN(g22415), .A(II28959) );
  INV_X1 NOT_7747( .ZN(II28962), .A(g21721) );
  INV_X1 NOT_7748( .ZN(g22418), .A(II28962) );
  INV_X1 NOT_7749( .ZN(g22421), .A(g21012) );
  INV_X1 NOT_7750( .ZN(II28966), .A(g20633) );
  INV_X1 NOT_7751( .ZN(g22422), .A(II28966) );
  INV_X1 NOT_7752( .ZN(II28969), .A(g21686) );
  INV_X1 NOT_7753( .ZN(g22425), .A(II28969) );
  INV_X1 NOT_7754( .ZN(II28972), .A(g21736) );
  INV_X1 NOT_7755( .ZN(g22428), .A(II28972) );
  INV_X1 NOT_7756( .ZN(II28975), .A(g21688) );
  INV_X1 NOT_7757( .ZN(g22431), .A(II28975) );
  INV_X1 NOT_7758( .ZN(II28978), .A(g21740) );
  INV_X1 NOT_7759( .ZN(g22434), .A(II28978) );
  INV_X1 NOT_7760( .ZN(II28981), .A(g21667) );
  INV_X1 NOT_7761( .ZN(g22437), .A(II28981) );
  INV_X1 NOT_7762( .ZN(II28984), .A(g21747) );
  INV_X1 NOT_7763( .ZN(g22440), .A(II28984) );
  INV_X1 NOT_7764( .ZN(g22443), .A(g21036) );
  INV_X1 NOT_7765( .ZN(II28988), .A(g20874) );
  INV_X1 NOT_7766( .ZN(g22444), .A(II28988) );
  INV_X1 NOT_7767( .ZN(II28991), .A(g20648) );
  INV_X1 NOT_7768( .ZN(g22445), .A(II28991) );
  INV_X1 NOT_7769( .ZN(II28994), .A(g21715) );
  INV_X1 NOT_7770( .ZN(g22448), .A(II28994) );
  INV_X1 NOT_7771( .ZN(II28997), .A(g21759) );
  INV_X1 NOT_7772( .ZN(g22451), .A(II28997) );
  INV_X1 NOT_7773( .ZN(II29001), .A(g20658) );
  INV_X1 NOT_7774( .ZN(g22455), .A(II29001) );
  INV_X1 NOT_7775( .ZN(II29004), .A(g21722) );
  INV_X1 NOT_7776( .ZN(g22458), .A(II29004) );
  INV_X1 NOT_7777( .ZN(II29007), .A(g21760) );
  INV_X1 NOT_7778( .ZN(g22461), .A(II29007) );
  INV_X1 NOT_7779( .ZN(II29010), .A(g21724) );
  INV_X1 NOT_7780( .ZN(g22464), .A(II29010) );
  INV_X1 NOT_7781( .ZN(II29013), .A(g21764) );
  INV_X1 NOT_7782( .ZN(g22467), .A(II29013) );
  INV_X1 NOT_7783( .ZN(II29016), .A(g21696) );
  INV_X1 NOT_7784( .ZN(g22470), .A(II29016) );
  INV_X1 NOT_7785( .ZN(II29019), .A(g21771) );
  INV_X1 NOT_7786( .ZN(g22473), .A(II29019) );
  INV_X1 NOT_7787( .ZN(g22476), .A(g21057) );
  INV_X1 NOT_7788( .ZN(II29023), .A(g20672) );
  INV_X1 NOT_7789( .ZN(g22477), .A(II29023) );
  INV_X1 NOT_7790( .ZN(II29026), .A(g21737) );
  INV_X1 NOT_7791( .ZN(g22480), .A(II29026) );
  INV_X1 NOT_7792( .ZN(II29030), .A(g20683) );
  INV_X1 NOT_7793( .ZN(g22484), .A(II29030) );
  INV_X1 NOT_7794( .ZN(II29033), .A(g21741) );
  INV_X1 NOT_7795( .ZN(g22487), .A(II29033) );
  INV_X1 NOT_7796( .ZN(II29036), .A(g21775) );
  INV_X1 NOT_7797( .ZN(g22490), .A(II29036) );
  INV_X1 NOT_7798( .ZN(II29040), .A(g20693) );
  INV_X1 NOT_7799( .ZN(g22494), .A(II29040) );
  INV_X1 NOT_7800( .ZN(II29043), .A(g21748) );
  INV_X1 NOT_7801( .ZN(g22497), .A(II29043) );
  INV_X1 NOT_7802( .ZN(II29046), .A(g21776) );
  INV_X1 NOT_7803( .ZN(g22500), .A(II29046) );
  INV_X1 NOT_7804( .ZN(II29049), .A(g21750) );
  INV_X1 NOT_7805( .ZN(g22503), .A(II29049) );
  INV_X1 NOT_7806( .ZN(II29052), .A(g21780) );
  INV_X1 NOT_7807( .ZN(g22506), .A(II29052) );
  INV_X1 NOT_7808( .ZN(II29055), .A(g21732) );
  INV_X1 NOT_7809( .ZN(g22509), .A(II29055) );
  INV_X1 NOT_7810( .ZN(II29058), .A(g20703) );
  INV_X1 NOT_7811( .ZN(g22512), .A(II29058) );
  INV_X1 NOT_7812( .ZN(II29064), .A(g20875) );
  INV_X1 NOT_7813( .ZN(g22518), .A(II29064) );
  INV_X1 NOT_7814( .ZN(II29067), .A(g20876) );
  INV_X1 NOT_7815( .ZN(g22519), .A(II29067) );
  INV_X4 NOT_7816( .ZN(II29070), .A(g20707) );
  INV_X4 NOT_7817( .ZN(g22520), .A(II29070) );
  INV_X4 NOT_7818( .ZN(II29073), .A(g21761) );
  INV_X1 NOT_7819( .ZN(g22523), .A(II29073) );
  INV_X1 NOT_7820( .ZN(II29077), .A(g20718) );
  INV_X1 NOT_7821( .ZN(g22527), .A(II29077) );
  INV_X1 NOT_7822( .ZN(II29080), .A(g21765) );
  INV_X1 NOT_7823( .ZN(g22530), .A(II29080) );
  INV_X1 NOT_7824( .ZN(II29083), .A(g21790) );
  INV_X1 NOT_7825( .ZN(g22533), .A(II29083) );
  INV_X1 NOT_7826( .ZN(II29087), .A(g20728) );
  INV_X1 NOT_7827( .ZN(g22537), .A(II29087) );
  INV_X1 NOT_7828( .ZN(II29090), .A(g21772) );
  INV_X1 NOT_7829( .ZN(g22540), .A(II29090) );
  INV_X1 NOT_7830( .ZN(II29093), .A(g21791) );
  INV_X1 NOT_7831( .ZN(g22543), .A(II29093) );
  INV_X1 NOT_7832( .ZN(g22547), .A(g21087) );
  INV_X1 NOT_7833( .ZN(II29098), .A(g20879) );
  INV_X1 NOT_7834( .ZN(g22548), .A(II29098) );
  INV_X1 NOT_7835( .ZN(II29101), .A(g20880) );
  INV_X1 NOT_7836( .ZN(g22549), .A(II29101) );
  INV_X1 NOT_7837( .ZN(II29104), .A(g20881) );
  INV_X1 NOT_7838( .ZN(g22550), .A(II29104) );
  INV_X1 NOT_7839( .ZN(II29107), .A(g21435) );
  INV_X1 NOT_7840( .ZN(g22551), .A(II29107) );
  INV_X1 NOT_7841( .ZN(II29110), .A(g20738) );
  INV_X1 NOT_7842( .ZN(g22552), .A(II29110) );
  INV_X1 NOT_7843( .ZN(II29116), .A(g20882) );
  INV_X1 NOT_7844( .ZN(g22558), .A(II29116) );
  INV_X1 NOT_7845( .ZN(II29119), .A(g20883) );
  INV_X1 NOT_7846( .ZN(g22559), .A(II29119) );
  INV_X1 NOT_7847( .ZN(II29122), .A(g20742) );
  INV_X1 NOT_7848( .ZN(g22560), .A(II29122) );
  INV_X1 NOT_7849( .ZN(II29125), .A(g21777) );
  INV_X1 NOT_7850( .ZN(g22563), .A(II29125) );
  INV_X1 NOT_7851( .ZN(II29129), .A(g20753) );
  INV_X1 NOT_7852( .ZN(g22567), .A(II29129) );
  INV_X1 NOT_7853( .ZN(II29132), .A(g21781) );
  INV_X1 NOT_7854( .ZN(g22570), .A(II29132) );
  INV_X1 NOT_7855( .ZN(II29135), .A(g21804) );
  INV_X1 NOT_7856( .ZN(g22573), .A(II29135) );
  INV_X1 NOT_7857( .ZN(II29142), .A(g20682) );
  INV_X1 NOT_7858( .ZN(g22582), .A(II29142) );
  INV_X1 NOT_7859( .ZN(II29145), .A(g20891) );
  INV_X1 NOT_7860( .ZN(g22583), .A(II29145) );
  INV_X1 NOT_7861( .ZN(II29148), .A(g20892) );
  INV_X1 NOT_7862( .ZN(g22584), .A(II29148) );
  INV_X1 NOT_7863( .ZN(II29151), .A(g20893) );
  INV_X1 NOT_7864( .ZN(g22585), .A(II29151) );
  INV_X1 NOT_7865( .ZN(II29154), .A(g20894) );
  INV_X1 NOT_7866( .ZN(g22586), .A(II29154) );
  INV_X1 NOT_7867( .ZN(g22588), .A(g21099) );
  INV_X1 NOT_7868( .ZN(II29159), .A(g20896) );
  INV_X1 NOT_7869( .ZN(g22589), .A(II29159) );
  INV_X1 NOT_7870( .ZN(II29162), .A(g20897) );
  INV_X1 NOT_7871( .ZN(g22590), .A(II29162) );
  INV_X1 NOT_7872( .ZN(II29165), .A(g20898) );
  INV_X1 NOT_7873( .ZN(g22591), .A(II29165) );
  INV_X1 NOT_7874( .ZN(II29168), .A(g20775) );
  INV_X1 NOT_7875( .ZN(g22592), .A(II29168) );
  INV_X1 NOT_7876( .ZN(II29174), .A(g20899) );
  INV_X1 NOT_7877( .ZN(g22598), .A(II29174) );
  INV_X1 NOT_7878( .ZN(II29177), .A(g20900) );
  INV_X1 NOT_7879( .ZN(g22599), .A(II29177) );
  INV_X1 NOT_7880( .ZN(II29180), .A(g20779) );
  INV_X1 NOT_7881( .ZN(g22600), .A(II29180) );
  INV_X1 NOT_7882( .ZN(II29183), .A(g21792) );
  INV_X1 NOT_7883( .ZN(g22603), .A(II29183) );
  INV_X1 NOT_7884( .ZN(g22609), .A(g21108) );
  INV_X1 NOT_7885( .ZN(II29191), .A(g20901) );
  INV_X1 NOT_7886( .ZN(g22611), .A(II29191) );
  INV_X1 NOT_7887( .ZN(II29194), .A(g20902) );
  INV_X1 NOT_7888( .ZN(g22612), .A(II29194) );
  INV_X1 NOT_7889( .ZN(II29197), .A(g20903) );
  INV_X1 NOT_7890( .ZN(g22613), .A(II29197) );
  INV_X1 NOT_7891( .ZN(II29203), .A(g20717) );
  INV_X1 NOT_7892( .ZN(g22619), .A(II29203) );
  INV_X1 NOT_7893( .ZN(II29206), .A(g20910) );
  INV_X1 NOT_7894( .ZN(g22620), .A(II29206) );
  INV_X1 NOT_7895( .ZN(II29209), .A(g20911) );
  INV_X1 NOT_7896( .ZN(g22621), .A(II29209) );
  INV_X1 NOT_7897( .ZN(II29212), .A(g20912) );
  INV_X1 NOT_7898( .ZN(g22622), .A(II29212) );
  INV_X1 NOT_7899( .ZN(II29215), .A(g20913) );
  INV_X1 NOT_7900( .ZN(g22623), .A(II29215) );
  INV_X1 NOT_7901( .ZN(g22625), .A(g21113) );
  INV_X1 NOT_7902( .ZN(II29220), .A(g20915) );
  INV_X1 NOT_7903( .ZN(g22626), .A(II29220) );
  INV_X1 NOT_7904( .ZN(II29223), .A(g20916) );
  INV_X1 NOT_7905( .ZN(g22627), .A(II29223) );
  INV_X1 NOT_7906( .ZN(II29226), .A(g20917) );
  INV_X1 NOT_7907( .ZN(g22628), .A(II29226) );
  INV_X1 NOT_7908( .ZN(II29229), .A(g20805) );
  INV_X1 NOT_7909( .ZN(g22629), .A(II29229) );
  INV_X1 NOT_7910( .ZN(II29235), .A(g20918) );
  INV_X1 NOT_7911( .ZN(g22635), .A(II29235) );
  INV_X1 NOT_7912( .ZN(II29238), .A(g20919) );
  INV_X1 NOT_7913( .ZN(g22636), .A(II29238) );
  INV_X1 NOT_7914( .ZN(II29243), .A(g20921) );
  INV_X1 NOT_7915( .ZN(g22639), .A(II29243) );
  INV_X1 NOT_7916( .ZN(II29246), .A(g20922) );
  INV_X1 NOT_7917( .ZN(g22640), .A(II29246) );
  INV_X1 NOT_7918( .ZN(II29249), .A(g20923) );
  INV_X1 NOT_7919( .ZN(g22641), .A(II29249) );
  INV_X1 NOT_7920( .ZN(II29252), .A(g20924) );
  INV_X1 NOT_7921( .ZN(g22642), .A(II29252) );
  INV_X1 NOT_7922( .ZN(g22645), .A(g21125) );
  INV_X1 NOT_7923( .ZN(II29259), .A(g20925) );
  INV_X1 NOT_7924( .ZN(g22647), .A(II29259) );
  INV_X1 NOT_7925( .ZN(II29262), .A(g20926) );
  INV_X1 NOT_7926( .ZN(g22648), .A(II29262) );
  INV_X1 NOT_7927( .ZN(II29265), .A(g20927) );
  INV_X1 NOT_7928( .ZN(g22649), .A(II29265) );
  INV_X1 NOT_7929( .ZN(II29271), .A(g20752) );
  INV_X1 NOT_7930( .ZN(g22655), .A(II29271) );
  INV_X1 NOT_7931( .ZN(II29274), .A(g20934) );
  INV_X1 NOT_7932( .ZN(g22656), .A(II29274) );
  INV_X1 NOT_7933( .ZN(II29277), .A(g20935) );
  INV_X1 NOT_7934( .ZN(g22657), .A(II29277) );
  INV_X1 NOT_7935( .ZN(II29280), .A(g20936) );
  INV_X1 NOT_7936( .ZN(g22658), .A(II29280) );
  INV_X1 NOT_7937( .ZN(II29283), .A(g20937) );
  INV_X1 NOT_7938( .ZN(g22659), .A(II29283) );
  INV_X1 NOT_7939( .ZN(g22661), .A(g21130) );
  INV_X1 NOT_7940( .ZN(II29288), .A(g20939) );
  INV_X1 NOT_7941( .ZN(g22662), .A(II29288) );
  INV_X1 NOT_7942( .ZN(II29291), .A(g20940) );
  INV_X1 NOT_7943( .ZN(g22663), .A(II29291) );
  INV_X1 NOT_7944( .ZN(II29294), .A(g20941) );
  INV_X1 NOT_7945( .ZN(g22664), .A(II29294) );
  INV_X1 NOT_7946( .ZN(II29301), .A(g20944) );
  INV_X1 NOT_7947( .ZN(g22669), .A(II29301) );
  INV_X1 NOT_7948( .ZN(II29304), .A(g20945) );
  INV_X1 NOT_7949( .ZN(g22670), .A(II29304) );
  INV_X1 NOT_7950( .ZN(II29307), .A(g20946) );
  INV_X1 NOT_7951( .ZN(g22671), .A(II29307) );
  INV_X1 NOT_7952( .ZN(II29310), .A(g20947) );
  INV_X1 NOT_7953( .ZN(g22672), .A(II29310) );
  INV_X1 NOT_7954( .ZN(II29313), .A(g20948) );
  INV_X1 NOT_7955( .ZN(g22673), .A(II29313) );
  INV_X1 NOT_7956( .ZN(II29317), .A(g20949) );
  INV_X1 NOT_7957( .ZN(g22675), .A(II29317) );
  INV_X1 NOT_7958( .ZN(II29320), .A(g20950) );
  INV_X1 NOT_7959( .ZN(g22676), .A(II29320) );
  INV_X1 NOT_7960( .ZN(II29323), .A(g20951) );
  INV_X1 NOT_7961( .ZN(g22677), .A(II29323) );
  INV_X1 NOT_7962( .ZN(II29326), .A(g20952) );
  INV_X1 NOT_7963( .ZN(g22678), .A(II29326) );
  INV_X1 NOT_7964( .ZN(g22681), .A(g21144) );
  INV_X1 NOT_7965( .ZN(II29333), .A(g20953) );
  INV_X1 NOT_7966( .ZN(g22683), .A(II29333) );
  INV_X1 NOT_7967( .ZN(II29336), .A(g20954) );
  INV_X1 NOT_7968( .ZN(g22684), .A(II29336) );
  INV_X1 NOT_7969( .ZN(II29339), .A(g20955) );
  INV_X1 NOT_7970( .ZN(g22685), .A(II29339) );
  INV_X1 NOT_7971( .ZN(II29345), .A(g20789) );
  INV_X1 NOT_7972( .ZN(g22691), .A(II29345) );
  INV_X1 NOT_7973( .ZN(II29348), .A(g20962) );
  INV_X1 NOT_7974( .ZN(g22692), .A(II29348) );
  INV_X1 NOT_7975( .ZN(II29351), .A(g20963) );
  INV_X1 NOT_7976( .ZN(g22693), .A(II29351) );
  INV_X1 NOT_7977( .ZN(II29354), .A(g20964) );
  INV_X1 NOT_7978( .ZN(g22694), .A(II29354) );
  INV_X1 NOT_7979( .ZN(II29357), .A(g20965) );
  INV_X1 NOT_7980( .ZN(g22695), .A(II29357) );
  INV_X1 NOT_7981( .ZN(II29360), .A(g21796) );
  INV_X1 NOT_7982( .ZN(g22696), .A(II29360) );
  INV_X1 NOT_7983( .ZN(II29366), .A(g20966) );
  INV_X1 NOT_7984( .ZN(g22702), .A(II29366) );
  INV_X4 NOT_7985( .ZN(II29369), .A(g20967) );
  INV_X4 NOT_7986( .ZN(g22703), .A(II29369) );
  INV_X4 NOT_7987( .ZN(II29372), .A(g20968) );
  INV_X1 NOT_7988( .ZN(g22704), .A(II29372) );
  INV_X1 NOT_7989( .ZN(II29375), .A(g20969) );
  INV_X1 NOT_7990( .ZN(g22705), .A(II29375) );
  INV_X1 NOT_7991( .ZN(II29378), .A(g20970) );
  INV_X1 NOT_7992( .ZN(g22706), .A(II29378) );
  INV_X1 NOT_7993( .ZN(II29383), .A(g20972) );
  INV_X1 NOT_7994( .ZN(g22709), .A(II29383) );
  INV_X1 NOT_7995( .ZN(II29386), .A(g20973) );
  INV_X1 NOT_7996( .ZN(g22710), .A(II29386) );
  INV_X1 NOT_7997( .ZN(II29389), .A(g20974) );
  INV_X1 NOT_7998( .ZN(g22711), .A(II29389) );
  INV_X1 NOT_7999( .ZN(II29392), .A(g20975) );
  INV_X1 NOT_8000( .ZN(g22712), .A(II29392) );
  INV_X1 NOT_8001( .ZN(II29395), .A(g20976) );
  INV_X1 NOT_8002( .ZN(g22713), .A(II29395) );
  INV_X1 NOT_8003( .ZN(II29399), .A(g20977) );
  INV_X1 NOT_8004( .ZN(g22715), .A(II29399) );
  INV_X1 NOT_8005( .ZN(II29402), .A(g20978) );
  INV_X1 NOT_8006( .ZN(g22716), .A(II29402) );
  INV_X1 NOT_8007( .ZN(II29405), .A(g20979) );
  INV_X1 NOT_8008( .ZN(g22717), .A(II29405) );
  INV_X1 NOT_8009( .ZN(II29408), .A(g20980) );
  INV_X1 NOT_8010( .ZN(g22718), .A(II29408) );
  INV_X1 NOT_8011( .ZN(g22721), .A(g21164) );
  INV_X1 NOT_8012( .ZN(II29415), .A(g20981) );
  INV_X1 NOT_8013( .ZN(g22723), .A(II29415) );
  INV_X1 NOT_8014( .ZN(II29418), .A(g20982) );
  INV_X1 NOT_8015( .ZN(g22724), .A(II29418) );
  INV_X1 NOT_8016( .ZN(II29421), .A(g20983) );
  INV_X1 NOT_8017( .ZN(g22725), .A(II29421) );
  INV_X1 NOT_8018( .ZN(II29426), .A(g20989) );
  INV_X1 NOT_8019( .ZN(g22728), .A(II29426) );
  INV_X1 NOT_8020( .ZN(II29429), .A(g20990) );
  INV_X1 NOT_8021( .ZN(g22729), .A(II29429) );
  INV_X1 NOT_8022( .ZN(II29432), .A(g20991) );
  INV_X1 NOT_8023( .ZN(g22730), .A(II29432) );
  INV_X1 NOT_8024( .ZN(II29435), .A(g20992) );
  INV_X1 NOT_8025( .ZN(g22731), .A(II29435) );
  INV_X1 NOT_8026( .ZN(II29439), .A(g20993) );
  INV_X1 NOT_8027( .ZN(g22733), .A(II29439) );
  INV_X1 NOT_8028( .ZN(II29442), .A(g20994) );
  INV_X1 NOT_8029( .ZN(g22734), .A(II29442) );
  INV_X1 NOT_8030( .ZN(II29445), .A(g20995) );
  INV_X1 NOT_8031( .ZN(g22735), .A(II29445) );
  INV_X1 NOT_8032( .ZN(II29448), .A(g20996) );
  INV_X1 NOT_8033( .ZN(g22736), .A(II29448) );
  INV_X1 NOT_8034( .ZN(II29451), .A(g20997) );
  INV_X1 NOT_8035( .ZN(g22737), .A(II29451) );
  INV_X1 NOT_8036( .ZN(II29456), .A(g20999) );
  INV_X1 NOT_8037( .ZN(g22740), .A(II29456) );
  INV_X1 NOT_8038( .ZN(II29459), .A(g21000) );
  INV_X1 NOT_8039( .ZN(g22741), .A(II29459) );
  INV_X1 NOT_8040( .ZN(II29462), .A(g21001) );
  INV_X1 NOT_8041( .ZN(g22742), .A(II29462) );
  INV_X1 NOT_8042( .ZN(II29465), .A(g21002) );
  INV_X1 NOT_8043( .ZN(g22743), .A(II29465) );
  INV_X1 NOT_8044( .ZN(II29468), .A(g21003) );
  INV_X1 NOT_8045( .ZN(g22744), .A(II29468) );
  INV_X1 NOT_8046( .ZN(II29472), .A(g21004) );
  INV_X1 NOT_8047( .ZN(g22746), .A(II29472) );
  INV_X1 NOT_8048( .ZN(II29475), .A(g21005) );
  INV_X1 NOT_8049( .ZN(g22747), .A(II29475) );
  INV_X1 NOT_8050( .ZN(II29478), .A(g21006) );
  INV_X1 NOT_8051( .ZN(g22748), .A(II29478) );
  INV_X1 NOT_8052( .ZN(II29481), .A(g21007) );
  INV_X1 NOT_8053( .ZN(g22749), .A(II29481) );
  INV_X1 NOT_8054( .ZN(II29484), .A(g21903) );
  INV_X1 NOT_8055( .ZN(g22750), .A(II29484) );
  INV_X1 NOT_8056( .ZN(g22753), .A(g21184) );
  INV_X1 NOT_8057( .ZN(II29490), .A(g21009) );
  INV_X1 NOT_8058( .ZN(g22756), .A(II29490) );
  INV_X1 NOT_8059( .ZN(II29493), .A(g21010) );
  INV_X1 NOT_8060( .ZN(g22757), .A(II29493) );
  INV_X1 NOT_8061( .ZN(II29496), .A(g21011) );
  INV_X1 NOT_8062( .ZN(g22758), .A(II29496) );
  INV_X1 NOT_8063( .ZN(II29500), .A(g21015) );
  INV_X1 NOT_8064( .ZN(g22760), .A(II29500) );
  INV_X1 NOT_8065( .ZN(II29503), .A(g21016) );
  INV_X1 NOT_8066( .ZN(g22761), .A(II29503) );
  INV_X1 NOT_8067( .ZN(II29506), .A(g21017) );
  INV_X1 NOT_8068( .ZN(g22762), .A(II29506) );
  INV_X1 NOT_8069( .ZN(II29509), .A(g21018) );
  INV_X1 NOT_8070( .ZN(g22763), .A(II29509) );
  INV_X1 NOT_8071( .ZN(II29513), .A(g21019) );
  INV_X1 NOT_8072( .ZN(g22765), .A(II29513) );
  INV_X1 NOT_8073( .ZN(II29516), .A(g21020) );
  INV_X1 NOT_8074( .ZN(g22766), .A(II29516) );
  INV_X1 NOT_8075( .ZN(II29519), .A(g21021) );
  INV_X1 NOT_8076( .ZN(g22767), .A(II29519) );
  INV_X1 NOT_8077( .ZN(II29522), .A(g21022) );
  INV_X1 NOT_8078( .ZN(g22768), .A(II29522) );
  INV_X1 NOT_8079( .ZN(II29525), .A(g21023) );
  INV_X1 NOT_8080( .ZN(g22769), .A(II29525) );
  INV_X1 NOT_8081( .ZN(II29530), .A(g21025) );
  INV_X1 NOT_8082( .ZN(g22772), .A(II29530) );
  INV_X1 NOT_8083( .ZN(II29533), .A(g21026) );
  INV_X1 NOT_8084( .ZN(g22773), .A(II29533) );
  INV_X1 NOT_8085( .ZN(II29536), .A(g21027) );
  INV_X1 NOT_8086( .ZN(g22774), .A(II29536) );
  INV_X1 NOT_8087( .ZN(II29539), .A(g21028) );
  INV_X1 NOT_8088( .ZN(g22775), .A(II29539) );
  INV_X1 NOT_8089( .ZN(II29542), .A(g21029) );
  INV_X1 NOT_8090( .ZN(g22776), .A(II29542) );
  INV_X1 NOT_8091( .ZN(g22777), .A(g21796) );
  INV_X1 NOT_8092( .ZN(II29547), .A(g21031) );
  INV_X1 NOT_8093( .ZN(g22785), .A(II29547) );
  INV_X1 NOT_8094( .ZN(II29550), .A(g21032) );
  INV_X1 NOT_8095( .ZN(g22786), .A(II29550) );
  INV_X1 NOT_8096( .ZN(g22787), .A(g21199) );
  INV_X1 NOT_8097( .ZN(II29556), .A(g21033) );
  INV_X1 NOT_8098( .ZN(g22790), .A(II29556) );
  INV_X1 NOT_8099( .ZN(II29559), .A(g21034) );
  INV_X1 NOT_8100( .ZN(g22791), .A(II29559) );
  INV_X1 NOT_8101( .ZN(II29562), .A(g21035) );
  INV_X1 NOT_8102( .ZN(g22792), .A(II29562) );
  INV_X1 NOT_8103( .ZN(II29566), .A(g21039) );
  INV_X1 NOT_8104( .ZN(g22794), .A(II29566) );
  INV_X1 NOT_8105( .ZN(II29569), .A(g21040) );
  INV_X1 NOT_8106( .ZN(g22795), .A(II29569) );
  INV_X1 NOT_8107( .ZN(II29572), .A(g21041) );
  INV_X1 NOT_8108( .ZN(g22796), .A(II29572) );
  INV_X1 NOT_8109( .ZN(II29575), .A(g21042) );
  INV_X1 NOT_8110( .ZN(g22797), .A(II29575) );
  INV_X1 NOT_8111( .ZN(II29579), .A(g21043) );
  INV_X1 NOT_8112( .ZN(g22799), .A(II29579) );
  INV_X1 NOT_8113( .ZN(II29582), .A(g21044) );
  INV_X1 NOT_8114( .ZN(g22800), .A(II29582) );
  INV_X1 NOT_8115( .ZN(II29585), .A(g21045) );
  INV_X1 NOT_8116( .ZN(g22801), .A(II29585) );
  INV_X1 NOT_8117( .ZN(II29588), .A(g21046) );
  INV_X1 NOT_8118( .ZN(g22802), .A(II29588) );
  INV_X1 NOT_8119( .ZN(II29591), .A(g21047) );
  INV_X1 NOT_8120( .ZN(g22803), .A(II29591) );
  INV_X1 NOT_8121( .ZN(g22805), .A(g21894) );
  INV_X1 NOT_8122( .ZN(g22806), .A(g21615) );
  INV_X1 NOT_8123( .ZN(II29600), .A(g21720) );
  INV_X1 NOT_8124( .ZN(g22812), .A(II29600) );
  INV_X1 NOT_8125( .ZN(II29603), .A(g21051) );
  INV_X1 NOT_8126( .ZN(g22824), .A(II29603) );
  INV_X1 NOT_8127( .ZN(II29606), .A(g21364) );
  INV_X1 NOT_8128( .ZN(g22825), .A(II29606) );
  INV_X1 NOT_8129( .ZN(II29610), .A(g21052) );
  INV_X1 NOT_8130( .ZN(g22827), .A(II29610) );
  INV_X1 NOT_8131( .ZN(II29613), .A(g21053) );
  INV_X1 NOT_8132( .ZN(g22828), .A(II29613) );
  INV_X1 NOT_8133( .ZN(g22829), .A(g21214) );
  INV_X1 NOT_8134( .ZN(II29619), .A(g21054) );
  INV_X1 NOT_8135( .ZN(g22832), .A(II29619) );
  INV_X1 NOT_8136( .ZN(II29622), .A(g21055) );
  INV_X1 NOT_8137( .ZN(g22833), .A(II29622) );
  INV_X1 NOT_8138( .ZN(II29625), .A(g21056) );
  INV_X1 NOT_8139( .ZN(g22834), .A(II29625) );
  INV_X1 NOT_8140( .ZN(II29629), .A(g21060) );
  INV_X1 NOT_8141( .ZN(g22836), .A(II29629) );
  INV_X1 NOT_8142( .ZN(II29632), .A(g21061) );
  INV_X1 NOT_8143( .ZN(g22837), .A(II29632) );
  INV_X1 NOT_8144( .ZN(II29635), .A(g21062) );
  INV_X1 NOT_8145( .ZN(g22838), .A(II29635) );
  INV_X1 NOT_8146( .ZN(II29638), .A(g21063) );
  INV_X1 NOT_8147( .ZN(g22839), .A(II29638) );
  INV_X1 NOT_8148( .ZN(II29641), .A(g20825) );
  INV_X1 NOT_8149( .ZN(g22840), .A(II29641) );
  INV_X1 NOT_8150( .ZN(g22843), .A(g21889) );
  INV_X1 NOT_8151( .ZN(g22847), .A(g21643) );
  INV_X1 NOT_8152( .ZN(II29653), .A(g21746) );
  INV_X1 NOT_8153( .ZN(g22852), .A(II29653) );
  INV_X1 NOT_8154( .ZN(II29656), .A(g21070) );
  INV_X1 NOT_8155( .ZN(g22864), .A(II29656) );
  INV_X1 NOT_8156( .ZN(II29660), .A(g21071) );
  INV_X1 NOT_8157( .ZN(g22866), .A(II29660) );
  INV_X1 NOT_8158( .ZN(II29663), .A(g21072) );
  INV_X1 NOT_8159( .ZN(g22867), .A(II29663) );
  INV_X8 NOT_8160( .ZN(g22868), .A(g21222) );
  INV_X8 NOT_8161( .ZN(II29669), .A(g21073) );
  INV_X1 NOT_8162( .ZN(g22871), .A(II29669) );
  INV_X1 NOT_8163( .ZN(II29672), .A(g21074) );
  INV_X1 NOT_8164( .ZN(g22872), .A(II29672) );
  INV_X1 NOT_8165( .ZN(II29675), .A(g21075) );
  INV_X1 NOT_8166( .ZN(g22873), .A(II29675) );
  INV_X1 NOT_8167( .ZN(g22875), .A(g21884) );
  INV_X1 NOT_8168( .ZN(g22882), .A(g21674) );
  INV_X1 NOT_8169( .ZN(II29687), .A(g21770) );
  INV_X1 NOT_8170( .ZN(g22887), .A(II29687) );
  INV_X1 NOT_8171( .ZN(II29690), .A(g21080) );
  INV_X1 NOT_8172( .ZN(g22899), .A(II29690) );
  INV_X1 NOT_8173( .ZN(II29694), .A(g21081) );
  INV_X1 NOT_8174( .ZN(g22901), .A(II29694) );
  INV_X1 NOT_8175( .ZN(II29697), .A(g21082) );
  INV_X1 NOT_8176( .ZN(g22902), .A(II29697) );
  INV_X1 NOT_8177( .ZN(II29700), .A(g20700) );
  INV_X1 NOT_8178( .ZN(g22903), .A(II29700) );
  INV_X1 NOT_8179( .ZN(g22907), .A(g21711) );
  INV_X1 NOT_8180( .ZN(g22917), .A(g21703) );
  INV_X1 NOT_8181( .ZN(II29712), .A(g21786) );
  INV_X1 NOT_8182( .ZN(g22922), .A(II29712) );
  INV_X1 NOT_8183( .ZN(II29715), .A(g21094) );
  INV_X1 NOT_8184( .ZN(g22934), .A(II29715) );
  INV_X1 NOT_8185( .ZN(II29724), .A(g21851) );
  INV_X1 NOT_8186( .ZN(g22945), .A(II29724) );
  INV_X1 NOT_8187( .ZN(II29727), .A(g20877) );
  INV_X1 NOT_8188( .ZN(g22948), .A(II29727) );
  INV_X1 NOT_8189( .ZN(g22949), .A(g21665) );
  INV_X1 NOT_8190( .ZN(g22954), .A(g21739) );
  INV_X1 NOT_8191( .ZN(g22958), .A(g21694) );
  INV_X1 NOT_8192( .ZN(g22962), .A(g21763) );
  INV_X1 NOT_8193( .ZN(g22966), .A(g21730) );
  INV_X1 NOT_8194( .ZN(II29736), .A(g20884) );
  INV_X1 NOT_8195( .ZN(g22970), .A(II29736) );
  INV_X1 NOT_8196( .ZN(g22971), .A(g21779) );
  INV_X1 NOT_8197( .ZN(g22975), .A(g21756) );
  INV_X1 NOT_8198( .ZN(II29741), .A(g21346) );
  INV_X1 NOT_8199( .ZN(g22979), .A(II29741) );
  INV_X1 NOT_8200( .ZN(g22980), .A(g21794) );
  INV_X1 NOT_8201( .ZN(g22986), .A(g21382) );
  INV_X1 NOT_8202( .ZN(g22988), .A(g21404) );
  INV_X1 NOT_8203( .ZN(g22989), .A(g21415) );
  INV_X1 NOT_8204( .ZN(g22991), .A(g21429) );
  INV_X1 NOT_8205( .ZN(g22995), .A(g21441) );
  INV_X1 NOT_8206( .ZN(g22996), .A(g21449) );
  INV_X1 NOT_8207( .ZN(g22998), .A(g21458) );
  INV_X1 NOT_8208( .ZN(g23001), .A(g21473) );
  INV_X1 NOT_8209( .ZN(g23002), .A(g21477) );
  INV_X1 NOT_8210( .ZN(g23006), .A(g21483) );
  INV_X1 NOT_8211( .ZN(g23007), .A(g21491) );
  INV_X1 NOT_8212( .ZN(g23008), .A(g21498) );
  INV_X1 NOT_8213( .ZN(g23012), .A(g21505) );
  INV_X1 NOT_8214( .ZN(g23015), .A(g21514) );
  INV_X1 NOT_8215( .ZN(g23016), .A(g21518) );
  INV_X1 NOT_8216( .ZN(g23020), .A(g21524) );
  INV_X1 NOT_8217( .ZN(g23021), .A(g21530) );
  INV_X1 NOT_8218( .ZN(g23024), .A(g21537) );
  INV_X1 NOT_8219( .ZN(g23028), .A(g21541) );
  INV_X1 NOT_8220( .ZN(g23031), .A(g21550) );
  INV_X1 NOT_8221( .ZN(g23032), .A(g21554) );
  INV_X1 NOT_8222( .ZN(g23036), .A(g21558) );
  INV_X1 NOT_8223( .ZN(g23037), .A(g21561) );
  INV_X1 NOT_8224( .ZN(g23038), .A(g21566) );
  INV_X1 NOT_8225( .ZN(g23041), .A(g21573) );
  INV_X1 NOT_8226( .ZN(g23045), .A(g21577) );
  INV_X1 NOT_8227( .ZN(g23048), .A(g21586) );
  INV_X1 NOT_8228( .ZN(g23049), .A(g21590) );
  INV_X1 NOT_8229( .ZN(II29797), .A(g21432) );
  INV_X1 NOT_8230( .ZN(g23050), .A(II29797) );
  INV_X1 NOT_8231( .ZN(II29802), .A(g21435) );
  INV_X1 NOT_8232( .ZN(g23055), .A(II29802) );
  INV_X1 NOT_8233( .ZN(g23056), .A(g21594) );
  INV_X1 NOT_8234( .ZN(g23057), .A(g21599) );
  INV_X1 NOT_8235( .ZN(g23060), .A(g21606) );
  INV_X1 NOT_8236( .ZN(g23064), .A(g21612) );
  INV_X1 NOT_8237( .ZN(II29812), .A(g21467) );
  INV_X1 NOT_8238( .ZN(g23065), .A(II29812) );
  INV_X1 NOT_8239( .ZN(II29817), .A(g21470) );
  INV_X1 NOT_8240( .ZN(g23068), .A(II29817) );
  INV_X1 NOT_8241( .ZN(g23069), .A(g21619) );
  INV_X1 NOT_8242( .ZN(g23074), .A(g21623) );
  INV_X1 NOT_8243( .ZN(g23075), .A(g21628) );
  INV_X1 NOT_8244( .ZN(II29827), .A(g21502) );
  INV_X1 NOT_8245( .ZN(g23078), .A(II29827) );
  INV_X1 NOT_8246( .ZN(g23079), .A(g21640) );
  INV_X1 NOT_8247( .ZN(g23082), .A(g21647) );
  INV_X1 NOT_8248( .ZN(g23087), .A(g21651) );
  INV_X1 NOT_8249( .ZN(g23088), .A(g21655) );
  INV_X1 NOT_8250( .ZN(II29841), .A(g21316) );
  INV_X1 NOT_8251( .ZN(g23094), .A(II29841) );
  INV_X1 NOT_8252( .ZN(g23095), .A(g21671) );
  INV_X1 NOT_8253( .ZN(g23098), .A(g21678) );
  INV_X1 NOT_8254( .ZN(g23103), .A(g21682) );
  INV_X1 NOT_8255( .ZN(II29852), .A(g21331) );
  INV_X1 NOT_8256( .ZN(g23105), .A(II29852) );
  INV_X1 NOT_8257( .ZN(g23112), .A(g21700) );
  INV_X1 NOT_8258( .ZN(g23115), .A(g21708) );
  INV_X1 NOT_8259( .ZN(II29863), .A(g21346) );
  INV_X1 NOT_8260( .ZN(g23116), .A(II29863) );
  INV_X1 NOT_8261( .ZN(II29872), .A(g21364) );
  INV_X1 NOT_8262( .ZN(g23125), .A(II29872) );
  INV_X1 NOT_8263( .ZN(II29881), .A(g21385) );
  INV_X1 NOT_8264( .ZN(g23134), .A(II29881) );
  INV_X1 NOT_8265( .ZN(g23140), .A(g21825) );
  INV_X1 NOT_8266( .ZN(g23141), .A(g21825) );
  INV_X1 NOT_8267( .ZN(g23142), .A(g21825) );
  INV_X1 NOT_8268( .ZN(g23143), .A(g21825) );
  INV_X1 NOT_8269( .ZN(g23144), .A(g21825) );
  INV_X1 NOT_8270( .ZN(g23145), .A(g21825) );
  INV_X1 NOT_8271( .ZN(g23146), .A(g21825) );
  INV_X1 NOT_8272( .ZN(g23147), .A(g21825) );
  INV_X1 NOT_8273( .ZN(II29897), .A(g23116) );
  INV_X1 NOT_8274( .ZN(g23148), .A(II29897) );
  INV_X1 NOT_8275( .ZN(II29900), .A(g23125) );
  INV_X1 NOT_8276( .ZN(g23149), .A(II29900) );
  INV_X1 NOT_8277( .ZN(II29903), .A(g23134) );
  INV_X1 NOT_8278( .ZN(g23150), .A(II29903) );
  INV_X1 NOT_8279( .ZN(II29906), .A(g21967) );
  INV_X1 NOT_8280( .ZN(g23151), .A(II29906) );
  INV_X1 NOT_8281( .ZN(II29909), .A(g23050) );
  INV_X1 NOT_8282( .ZN(g23152), .A(II29909) );
  INV_X1 NOT_8283( .ZN(II29912), .A(g23065) );
  INV_X1 NOT_8284( .ZN(g23153), .A(II29912) );
  INV_X1 NOT_8285( .ZN(II29915), .A(g23055) );
  INV_X1 NOT_8286( .ZN(g23154), .A(II29915) );
  INV_X1 NOT_8287( .ZN(II29918), .A(g23068) );
  INV_X1 NOT_8288( .ZN(g23155), .A(II29918) );
  INV_X1 NOT_8289( .ZN(II29921), .A(g23078) );
  INV_X1 NOT_8290( .ZN(g23156), .A(II29921) );
  INV_X1 NOT_8291( .ZN(II29924), .A(g23094) );
  INV_X1 NOT_8292( .ZN(g23157), .A(II29924) );
  INV_X1 NOT_8293( .ZN(II29927), .A(g23105) );
  INV_X1 NOT_8294( .ZN(g23158), .A(II29927) );
  INV_X1 NOT_8295( .ZN(II29930), .A(g22176) );
  INV_X1 NOT_8296( .ZN(g23159), .A(II29930) );
  INV_X1 NOT_8297( .ZN(II29933), .A(g22082) );
  INV_X1 NOT_8298( .ZN(g23160), .A(II29933) );
  INV_X1 NOT_8299( .ZN(II29936), .A(g22582) );
  INV_X1 NOT_8300( .ZN(g23161), .A(II29936) );
  INV_X1 NOT_8301( .ZN(II29939), .A(g22518) );
  INV_X1 NOT_8302( .ZN(g23162), .A(II29939) );
  INV_X1 NOT_8303( .ZN(II29942), .A(g22548) );
  INV_X1 NOT_8304( .ZN(g23163), .A(II29942) );
  INV_X1 NOT_8305( .ZN(II29945), .A(g22583) );
  INV_X1 NOT_8306( .ZN(g23164), .A(II29945) );
  INV_X1 NOT_8307( .ZN(II29948), .A(g22549) );
  INV_X1 NOT_8308( .ZN(g23165), .A(II29948) );
  INV_X1 NOT_8309( .ZN(II29951), .A(g22584) );
  INV_X1 NOT_8310( .ZN(g23166), .A(II29951) );
  INV_X1 NOT_8311( .ZN(II29954), .A(g22611) );
  INV_X1 NOT_8312( .ZN(g23167), .A(II29954) );
  INV_X1 NOT_8313( .ZN(II29957), .A(g22585) );
  INV_X1 NOT_8314( .ZN(g23168), .A(II29957) );
  INV_X1 NOT_8315( .ZN(II29960), .A(g22612) );
  INV_X1 NOT_8316( .ZN(g23169), .A(II29960) );
  INV_X1 NOT_8317( .ZN(II29963), .A(g22639) );
  INV_X1 NOT_8318( .ZN(g23170), .A(II29963) );
  INV_X1 NOT_8319( .ZN(II29966), .A(g22613) );
  INV_X1 NOT_8320( .ZN(g23171), .A(II29966) );
  INV_X1 NOT_8321( .ZN(II29969), .A(g22640) );
  INV_X1 NOT_8322( .ZN(g23172), .A(II29969) );
  INV_X1 NOT_8323( .ZN(II29972), .A(g22669) );
  INV_X1 NOT_8324( .ZN(g23173), .A(II29972) );
  INV_X1 NOT_8325( .ZN(II29975), .A(g22641) );
  INV_X1 NOT_8326( .ZN(g23174), .A(II29975) );
  INV_X1 NOT_8327( .ZN(II29978), .A(g22670) );
  INV_X1 NOT_8328( .ZN(g23175), .A(II29978) );
  INV_X1 NOT_8329( .ZN(II29981), .A(g22702) );
  INV_X1 NOT_8330( .ZN(g23176), .A(II29981) );
  INV_X1 NOT_8331( .ZN(II29984), .A(g22671) );
  INV_X1 NOT_8332( .ZN(g23177), .A(II29984) );
  INV_X1 NOT_8333( .ZN(II29987), .A(g22703) );
  INV_X1 NOT_8334( .ZN(g23178), .A(II29987) );
  INV_X1 NOT_8335( .ZN(II29990), .A(g22728) );
  INV_X1 NOT_8336( .ZN(g23179), .A(II29990) );
  INV_X8 NOT_8337( .ZN(II29993), .A(g22704) );
  INV_X8 NOT_8338( .ZN(g23180), .A(II29993) );
  INV_X1 NOT_8339( .ZN(II29996), .A(g22729) );
  INV_X1 NOT_8340( .ZN(g23181), .A(II29996) );
  INV_X1 NOT_8341( .ZN(II29999), .A(g22756) );
  INV_X1 NOT_8342( .ZN(g23182), .A(II29999) );
  INV_X1 NOT_8343( .ZN(II30002), .A(g22730) );
  INV_X1 NOT_8344( .ZN(g23183), .A(II30002) );
  INV_X1 NOT_8345( .ZN(II30005), .A(g22757) );
  INV_X1 NOT_8346( .ZN(g23184), .A(II30005) );
  INV_X1 NOT_8347( .ZN(II30008), .A(g22785) );
  INV_X1 NOT_8348( .ZN(g23185), .A(II30008) );
  INV_X1 NOT_8349( .ZN(II30011), .A(g22758) );
  INV_X1 NOT_8350( .ZN(g23186), .A(II30011) );
  INV_X1 NOT_8351( .ZN(II30014), .A(g22786) );
  INV_X1 NOT_8352( .ZN(g23187), .A(II30014) );
  INV_X1 NOT_8353( .ZN(II30017), .A(g22824) );
  INV_X1 NOT_8354( .ZN(g23188), .A(II30017) );
  INV_X1 NOT_8355( .ZN(II30020), .A(g22519) );
  INV_X1 NOT_8356( .ZN(g23189), .A(II30020) );
  INV_X1 NOT_8357( .ZN(II30023), .A(g22550) );
  INV_X1 NOT_8358( .ZN(g23190), .A(II30023) );
  INV_X1 NOT_8359( .ZN(II30026), .A(g22586) );
  INV_X1 NOT_8360( .ZN(g23191), .A(II30026) );
  INV_X1 NOT_8361( .ZN(II30029), .A(g22642) );
  INV_X1 NOT_8362( .ZN(g23192), .A(II30029) );
  INV_X1 NOT_8363( .ZN(II30032), .A(g22672) );
  INV_X1 NOT_8364( .ZN(g23193), .A(II30032) );
  INV_X1 NOT_8365( .ZN(II30035), .A(g22705) );
  INV_X1 NOT_8366( .ZN(g23194), .A(II30035) );
  INV_X1 NOT_8367( .ZN(II30038), .A(g22673) );
  INV_X1 NOT_8368( .ZN(g23195), .A(II30038) );
  INV_X1 NOT_8369( .ZN(II30041), .A(g22706) );
  INV_X1 NOT_8370( .ZN(g23196), .A(II30041) );
  INV_X1 NOT_8371( .ZN(II30044), .A(g22731) );
  INV_X1 NOT_8372( .ZN(g23197), .A(II30044) );
  INV_X1 NOT_8373( .ZN(II30047), .A(g22107) );
  INV_X1 NOT_8374( .ZN(g23198), .A(II30047) );
  INV_X1 NOT_8375( .ZN(II30050), .A(g22619) );
  INV_X1 NOT_8376( .ZN(g23199), .A(II30050) );
  INV_X1 NOT_8377( .ZN(II30053), .A(g22558) );
  INV_X1 NOT_8378( .ZN(g23200), .A(II30053) );
  INV_X1 NOT_8379( .ZN(II30056), .A(g22589) );
  INV_X1 NOT_8380( .ZN(g23201), .A(II30056) );
  INV_X1 NOT_8381( .ZN(II30059), .A(g22620) );
  INV_X1 NOT_8382( .ZN(g23202), .A(II30059) );
  INV_X1 NOT_8383( .ZN(II30062), .A(g22590) );
  INV_X1 NOT_8384( .ZN(g23203), .A(II30062) );
  INV_X1 NOT_8385( .ZN(II30065), .A(g22621) );
  INV_X1 NOT_8386( .ZN(g23204), .A(II30065) );
  INV_X1 NOT_8387( .ZN(II30068), .A(g22647) );
  INV_X1 NOT_8388( .ZN(g23205), .A(II30068) );
  INV_X1 NOT_8389( .ZN(II30071), .A(g22622) );
  INV_X1 NOT_8390( .ZN(g23206), .A(II30071) );
  INV_X1 NOT_8391( .ZN(II30074), .A(g22648) );
  INV_X1 NOT_8392( .ZN(g23207), .A(II30074) );
  INV_X1 NOT_8393( .ZN(II30077), .A(g22675) );
  INV_X1 NOT_8394( .ZN(g23208), .A(II30077) );
  INV_X1 NOT_8395( .ZN(II30080), .A(g22649) );
  INV_X1 NOT_8396( .ZN(g23209), .A(II30080) );
  INV_X1 NOT_8397( .ZN(II30083), .A(g22676) );
  INV_X1 NOT_8398( .ZN(g23210), .A(II30083) );
  INV_X1 NOT_8399( .ZN(II30086), .A(g22709) );
  INV_X1 NOT_8400( .ZN(g23211), .A(II30086) );
  INV_X1 NOT_8401( .ZN(II30089), .A(g22677) );
  INV_X1 NOT_8402( .ZN(g23212), .A(II30089) );
  INV_X1 NOT_8403( .ZN(II30092), .A(g22710) );
  INV_X1 NOT_8404( .ZN(g23213), .A(II30092) );
  INV_X1 NOT_8405( .ZN(II30095), .A(g22733) );
  INV_X1 NOT_8406( .ZN(g23214), .A(II30095) );
  INV_X1 NOT_8407( .ZN(II30098), .A(g22711) );
  INV_X1 NOT_8408( .ZN(g23215), .A(II30098) );
  INV_X1 NOT_8409( .ZN(II30101), .A(g22734) );
  INV_X1 NOT_8410( .ZN(g23216), .A(II30101) );
  INV_X1 NOT_8411( .ZN(II30104), .A(g22760) );
  INV_X1 NOT_8412( .ZN(g23217), .A(II30104) );
  INV_X1 NOT_8413( .ZN(II30107), .A(g22735) );
  INV_X1 NOT_8414( .ZN(g23218), .A(II30107) );
  INV_X1 NOT_8415( .ZN(II30110), .A(g22761) );
  INV_X1 NOT_8416( .ZN(g23219), .A(II30110) );
  INV_X1 NOT_8417( .ZN(II30113), .A(g22790) );
  INV_X1 NOT_8418( .ZN(g23220), .A(II30113) );
  INV_X1 NOT_8419( .ZN(II30116), .A(g22762) );
  INV_X1 NOT_8420( .ZN(g23221), .A(II30116) );
  INV_X1 NOT_8421( .ZN(II30119), .A(g22791) );
  INV_X1 NOT_8422( .ZN(g23222), .A(II30119) );
  INV_X1 NOT_8423( .ZN(II30122), .A(g22827) );
  INV_X1 NOT_8424( .ZN(g23223), .A(II30122) );
  INV_X1 NOT_8425( .ZN(II30125), .A(g22792) );
  INV_X1 NOT_8426( .ZN(g23224), .A(II30125) );
  INV_X1 NOT_8427( .ZN(II30128), .A(g22828) );
  INV_X1 NOT_8428( .ZN(g23225), .A(II30128) );
  INV_X1 NOT_8429( .ZN(II30131), .A(g22864) );
  INV_X1 NOT_8430( .ZN(g23226), .A(II30131) );
  INV_X1 NOT_8431( .ZN(II30134), .A(g22559) );
  INV_X1 NOT_8432( .ZN(g23227), .A(II30134) );
  INV_X1 NOT_8433( .ZN(II30137), .A(g22591) );
  INV_X1 NOT_8434( .ZN(g23228), .A(II30137) );
  INV_X1 NOT_8435( .ZN(II30140), .A(g22623) );
  INV_X1 NOT_8436( .ZN(g23229), .A(II30140) );
  INV_X1 NOT_8437( .ZN(II30143), .A(g22678) );
  INV_X1 NOT_8438( .ZN(g23230), .A(II30143) );
  INV_X1 NOT_8439( .ZN(II30146), .A(g22712) );
  INV_X1 NOT_8440( .ZN(g23231), .A(II30146) );
  INV_X1 NOT_8441( .ZN(II30149), .A(g22736) );
  INV_X1 NOT_8442( .ZN(g23232), .A(II30149) );
  INV_X1 NOT_8443( .ZN(II30152), .A(g22713) );
  INV_X1 NOT_8444( .ZN(g23233), .A(II30152) );
  INV_X1 NOT_8445( .ZN(II30155), .A(g22737) );
  INV_X1 NOT_8446( .ZN(g23234), .A(II30155) );
  INV_X1 NOT_8447( .ZN(II30158), .A(g22763) );
  INV_X1 NOT_8448( .ZN(g23235), .A(II30158) );
  INV_X1 NOT_8449( .ZN(II30161), .A(g22133) );
  INV_X1 NOT_8450( .ZN(g23236), .A(II30161) );
  INV_X1 NOT_8451( .ZN(II30164), .A(g22655) );
  INV_X8 NOT_8452( .ZN(g23237), .A(II30164) );
  INV_X8 NOT_8453( .ZN(II30167), .A(g22598) );
  INV_X1 NOT_8454( .ZN(g23238), .A(II30167) );
  INV_X1 NOT_8455( .ZN(II30170), .A(g22626) );
  INV_X1 NOT_8456( .ZN(g23239), .A(II30170) );
  INV_X1 NOT_8457( .ZN(II30173), .A(g22656) );
  INV_X1 NOT_8458( .ZN(g23240), .A(II30173) );
  INV_X1 NOT_8459( .ZN(II30176), .A(g22627) );
  INV_X1 NOT_8460( .ZN(g23241), .A(II30176) );
  INV_X1 NOT_8461( .ZN(II30179), .A(g22657) );
  INV_X1 NOT_8462( .ZN(g23242), .A(II30179) );
  INV_X1 NOT_8463( .ZN(II30182), .A(g22683) );
  INV_X1 NOT_8464( .ZN(g23243), .A(II30182) );
  INV_X1 NOT_8465( .ZN(II30185), .A(g22658) );
  INV_X1 NOT_8466( .ZN(g23244), .A(II30185) );
  INV_X1 NOT_8467( .ZN(II30188), .A(g22684) );
  INV_X1 NOT_8468( .ZN(g23245), .A(II30188) );
  INV_X1 NOT_8469( .ZN(II30191), .A(g22715) );
  INV_X1 NOT_8470( .ZN(g23246), .A(II30191) );
  INV_X1 NOT_8471( .ZN(II30194), .A(g22685) );
  INV_X1 NOT_8472( .ZN(g23247), .A(II30194) );
  INV_X1 NOT_8473( .ZN(II30197), .A(g22716) );
  INV_X1 NOT_8474( .ZN(g23248), .A(II30197) );
  INV_X1 NOT_8475( .ZN(II30200), .A(g22740) );
  INV_X1 NOT_8476( .ZN(g23249), .A(II30200) );
  INV_X1 NOT_8477( .ZN(II30203), .A(g22717) );
  INV_X1 NOT_8478( .ZN(g23250), .A(II30203) );
  INV_X1 NOT_8479( .ZN(II30206), .A(g22741) );
  INV_X1 NOT_8480( .ZN(g23251), .A(II30206) );
  INV_X1 NOT_8481( .ZN(II30209), .A(g22765) );
  INV_X1 NOT_8482( .ZN(g23252), .A(II30209) );
  INV_X1 NOT_8483( .ZN(II30212), .A(g22742) );
  INV_X1 NOT_8484( .ZN(g23253), .A(II30212) );
  INV_X1 NOT_8485( .ZN(II30215), .A(g22766) );
  INV_X1 NOT_8486( .ZN(g23254), .A(II30215) );
  INV_X1 NOT_8487( .ZN(II30218), .A(g22794) );
  INV_X1 NOT_8488( .ZN(g23255), .A(II30218) );
  INV_X1 NOT_8489( .ZN(II30221), .A(g22767) );
  INV_X1 NOT_8490( .ZN(g23256), .A(II30221) );
  INV_X1 NOT_8491( .ZN(II30224), .A(g22795) );
  INV_X1 NOT_8492( .ZN(g23257), .A(II30224) );
  INV_X1 NOT_8493( .ZN(II30227), .A(g22832) );
  INV_X1 NOT_8494( .ZN(g23258), .A(II30227) );
  INV_X1 NOT_8495( .ZN(II30230), .A(g22796) );
  INV_X1 NOT_8496( .ZN(g23259), .A(II30230) );
  INV_X1 NOT_8497( .ZN(II30233), .A(g22833) );
  INV_X1 NOT_8498( .ZN(g23260), .A(II30233) );
  INV_X1 NOT_8499( .ZN(II30236), .A(g22866) );
  INV_X1 NOT_8500( .ZN(g23261), .A(II30236) );
  INV_X1 NOT_8501( .ZN(II30239), .A(g22834) );
  INV_X1 NOT_8502( .ZN(g23262), .A(II30239) );
  INV_X1 NOT_8503( .ZN(II30242), .A(g22867) );
  INV_X1 NOT_8504( .ZN(g23263), .A(II30242) );
  INV_X1 NOT_8505( .ZN(II30245), .A(g22899) );
  INV_X1 NOT_8506( .ZN(g23264), .A(II30245) );
  INV_X1 NOT_8507( .ZN(II30248), .A(g22599) );
  INV_X1 NOT_8508( .ZN(g23265), .A(II30248) );
  INV_X1 NOT_8509( .ZN(II30251), .A(g22628) );
  INV_X1 NOT_8510( .ZN(g23266), .A(II30251) );
  INV_X1 NOT_8511( .ZN(II30254), .A(g22659) );
  INV_X1 NOT_8512( .ZN(g23267), .A(II30254) );
  INV_X1 NOT_8513( .ZN(II30257), .A(g22718) );
  INV_X1 NOT_8514( .ZN(g23268), .A(II30257) );
  INV_X1 NOT_8515( .ZN(II30260), .A(g22743) );
  INV_X1 NOT_8516( .ZN(g23269), .A(II30260) );
  INV_X1 NOT_8517( .ZN(II30263), .A(g22768) );
  INV_X1 NOT_8518( .ZN(g23270), .A(II30263) );
  INV_X1 NOT_8519( .ZN(II30266), .A(g22744) );
  INV_X1 NOT_8520( .ZN(g23271), .A(II30266) );
  INV_X1 NOT_8521( .ZN(II30269), .A(g22769) );
  INV_X1 NOT_8522( .ZN(g23272), .A(II30269) );
  INV_X1 NOT_8523( .ZN(II30272), .A(g22797) );
  INV_X1 NOT_8524( .ZN(g23273), .A(II30272) );
  INV_X1 NOT_8525( .ZN(II30275), .A(g22156) );
  INV_X1 NOT_8526( .ZN(g23274), .A(II30275) );
  INV_X1 NOT_8527( .ZN(II30278), .A(g22691) );
  INV_X1 NOT_8528( .ZN(g23275), .A(II30278) );
  INV_X1 NOT_8529( .ZN(II30281), .A(g22635) );
  INV_X1 NOT_8530( .ZN(g23276), .A(II30281) );
  INV_X1 NOT_8531( .ZN(II30284), .A(g22662) );
  INV_X1 NOT_8532( .ZN(g23277), .A(II30284) );
  INV_X1 NOT_8533( .ZN(II30287), .A(g22692) );
  INV_X1 NOT_8534( .ZN(g23278), .A(II30287) );
  INV_X1 NOT_8535( .ZN(II30290), .A(g22663) );
  INV_X1 NOT_8536( .ZN(g23279), .A(II30290) );
  INV_X1 NOT_8537( .ZN(II30293), .A(g22693) );
  INV_X1 NOT_8538( .ZN(g23280), .A(II30293) );
  INV_X1 NOT_8539( .ZN(II30296), .A(g22723) );
  INV_X1 NOT_8540( .ZN(g23281), .A(II30296) );
  INV_X1 NOT_8541( .ZN(II30299), .A(g22694) );
  INV_X1 NOT_8542( .ZN(g23282), .A(II30299) );
  INV_X1 NOT_8543( .ZN(II30302), .A(g22724) );
  INV_X1 NOT_8544( .ZN(g23283), .A(II30302) );
  INV_X1 NOT_8545( .ZN(II30305), .A(g22746) );
  INV_X1 NOT_8546( .ZN(g23284), .A(II30305) );
  INV_X1 NOT_8547( .ZN(II30308), .A(g22725) );
  INV_X1 NOT_8548( .ZN(g23285), .A(II30308) );
  INV_X1 NOT_8549( .ZN(II30311), .A(g22747) );
  INV_X1 NOT_8550( .ZN(g23286), .A(II30311) );
  INV_X1 NOT_8551( .ZN(II30314), .A(g22772) );
  INV_X1 NOT_8552( .ZN(g23287), .A(II30314) );
  INV_X1 NOT_8553( .ZN(II30317), .A(g22748) );
  INV_X1 NOT_8554( .ZN(g23288), .A(II30317) );
  INV_X1 NOT_8555( .ZN(II30320), .A(g22773) );
  INV_X1 NOT_8556( .ZN(g23289), .A(II30320) );
  INV_X1 NOT_8557( .ZN(II30323), .A(g22799) );
  INV_X1 NOT_8558( .ZN(g23290), .A(II30323) );
  INV_X1 NOT_8559( .ZN(II30326), .A(g22774) );
  INV_X1 NOT_8560( .ZN(g23291), .A(II30326) );
  INV_X1 NOT_8561( .ZN(II30329), .A(g22800) );
  INV_X1 NOT_8562( .ZN(g23292), .A(II30329) );
  INV_X1 NOT_8563( .ZN(II30332), .A(g22836) );
  INV_X1 NOT_8564( .ZN(g23293), .A(II30332) );
  INV_X1 NOT_8565( .ZN(II30335), .A(g22801) );
  INV_X1 NOT_8566( .ZN(g23294), .A(II30335) );
  INV_X1 NOT_8567( .ZN(II30338), .A(g22837) );
  INV_X1 NOT_8568( .ZN(g23295), .A(II30338) );
  INV_X1 NOT_8569( .ZN(II30341), .A(g22871) );
  INV_X8 NOT_8570( .ZN(g23296), .A(II30341) );
  INV_X8 NOT_8571( .ZN(II30344), .A(g22838) );
  INV_X1 NOT_8572( .ZN(g23297), .A(II30344) );
  INV_X1 NOT_8573( .ZN(II30347), .A(g22872) );
  INV_X1 NOT_8574( .ZN(g23298), .A(II30347) );
  INV_X1 NOT_8575( .ZN(II30350), .A(g22901) );
  INV_X1 NOT_8576( .ZN(g23299), .A(II30350) );
  INV_X1 NOT_8577( .ZN(II30353), .A(g22873) );
  INV_X1 NOT_8578( .ZN(g23300), .A(II30353) );
  INV_X1 NOT_8579( .ZN(II30356), .A(g22902) );
  INV_X1 NOT_8580( .ZN(g23301), .A(II30356) );
  INV_X1 NOT_8581( .ZN(II30359), .A(g22934) );
  INV_X1 NOT_8582( .ZN(g23302), .A(II30359) );
  INV_X1 NOT_8583( .ZN(II30362), .A(g22636) );
  INV_X1 NOT_8584( .ZN(g23303), .A(II30362) );
  INV_X1 NOT_8585( .ZN(II30365), .A(g22664) );
  INV_X1 NOT_8586( .ZN(g23304), .A(II30365) );
  INV_X1 NOT_8587( .ZN(II30368), .A(g22695) );
  INV_X1 NOT_8588( .ZN(g23305), .A(II30368) );
  INV_X1 NOT_8589( .ZN(II30371), .A(g22749) );
  INV_X1 NOT_8590( .ZN(g23306), .A(II30371) );
  INV_X1 NOT_8591( .ZN(II30374), .A(g22775) );
  INV_X1 NOT_8592( .ZN(g23307), .A(II30374) );
  INV_X1 NOT_8593( .ZN(II30377), .A(g22802) );
  INV_X1 NOT_8594( .ZN(g23308), .A(II30377) );
  INV_X1 NOT_8595( .ZN(II30380), .A(g22776) );
  INV_X1 NOT_8596( .ZN(g23309), .A(II30380) );
  INV_X1 NOT_8597( .ZN(II30383), .A(g22803) );
  INV_X1 NOT_8598( .ZN(g23310), .A(II30383) );
  INV_X1 NOT_8599( .ZN(II30386), .A(g22839) );
  INV_X1 NOT_8600( .ZN(g23311), .A(II30386) );
  INV_X1 NOT_8601( .ZN(II30389), .A(g22225) );
  INV_X1 NOT_8602( .ZN(g23312), .A(II30389) );
  INV_X1 NOT_8603( .ZN(II30392), .A(g22226) );
  INV_X1 NOT_8604( .ZN(g23313), .A(II30392) );
  INV_X1 NOT_8605( .ZN(II30395), .A(g22253) );
  INV_X1 NOT_8606( .ZN(g23314), .A(II30395) );
  INV_X1 NOT_8607( .ZN(II30398), .A(g22840) );
  INV_X1 NOT_8608( .ZN(g23315), .A(II30398) );
  INV_X1 NOT_8609( .ZN(II30401), .A(g22444) );
  INV_X1 NOT_8610( .ZN(g23316), .A(II30401) );
  INV_X1 NOT_8611( .ZN(II30404), .A(g22948) );
  INV_X1 NOT_8612( .ZN(g23317), .A(II30404) );
  INV_X1 NOT_8613( .ZN(II30407), .A(g22970) );
  INV_X1 NOT_8614( .ZN(g23318), .A(II30407) );
  INV_X1 NOT_8615( .ZN(g23403), .A(g23052) );
  INV_X1 NOT_8616( .ZN(g23410), .A(g23071) );
  INV_X1 NOT_8617( .ZN(g23415), .A(g23084) );
  INV_X1 NOT_8618( .ZN(g23420), .A(g23089) );
  INV_X1 NOT_8619( .ZN(g23424), .A(g23100) );
  INV_X1 NOT_8620( .ZN(g23429), .A(g23107) );
  INV_X1 NOT_8621( .ZN(g23435), .A(g23120) );
  INV_X1 NOT_8622( .ZN(II30467), .A(g23000) );
  INV_X1 NOT_8623( .ZN(g23438), .A(II30467) );
  INV_X1 NOT_8624( .ZN(II30470), .A(g23117) );
  INV_X1 NOT_8625( .ZN(g23439), .A(II30470) );
  INV_X1 NOT_8626( .ZN(g23441), .A(g23129) );
  INV_X1 NOT_8627( .ZN(g23444), .A(g22945) );
  INV_X1 NOT_8628( .ZN(II30476), .A(g22876) );
  INV_X1 NOT_8629( .ZN(g23448), .A(II30476) );
  INV_X1 NOT_8630( .ZN(II30480), .A(g23014) );
  INV_X1 NOT_8631( .ZN(g23452), .A(II30480) );
  INV_X1 NOT_8632( .ZN(II30483), .A(g23126) );
  INV_X1 NOT_8633( .ZN(g23453), .A(II30483) );
  INV_X1 NOT_8634( .ZN(II30486), .A(g23022) );
  INV_X1 NOT_8635( .ZN(g23454), .A(II30486) );
  INV_X1 NOT_8636( .ZN(II30489), .A(g22911) );
  INV_X1 NOT_8637( .ZN(g23455), .A(II30489) );
  INV_X1 NOT_8638( .ZN(II30493), .A(g23030) );
  INV_X1 NOT_8639( .ZN(g23459), .A(II30493) );
  INV_X1 NOT_8640( .ZN(II30496), .A(g23137) );
  INV_X1 NOT_8641( .ZN(g23460), .A(II30496) );
  INV_X1 NOT_8642( .ZN(II30501), .A(g23039) );
  INV_X1 NOT_8643( .ZN(g23463), .A(II30501) );
  INV_X1 NOT_8644( .ZN(II30504), .A(g22936) );
  INV_X1 NOT_8645( .ZN(g23464), .A(II30504) );
  INV_X1 NOT_8646( .ZN(II30508), .A(g23047) );
  INV_X1 NOT_8647( .ZN(g23468), .A(II30508) );
  INV_X1 NOT_8648( .ZN(II30511), .A(g21970) );
  INV_X1 NOT_8649( .ZN(g23469), .A(II30511) );
  INV_X1 NOT_8650( .ZN(g23470), .A(g22188) );
  INV_X1 NOT_8651( .ZN(II30516), .A(g23058) );
  INV_X1 NOT_8652( .ZN(g23472), .A(II30516) );
  INV_X1 NOT_8653( .ZN(II30519), .A(g22942) );
  INV_X1 NOT_8654( .ZN(g23473), .A(II30519) );
  INV_X1 NOT_8655( .ZN(II30525), .A(g23067) );
  INV_X1 NOT_8656( .ZN(g23481), .A(II30525) );
  INV_X1 NOT_8657( .ZN(g23482), .A(g22197) );
  INV_X1 NOT_8658( .ZN(II30531), .A(g23076) );
  INV_X1 NOT_8659( .ZN(g23485), .A(II30531) );
  INV_X1 NOT_8660( .ZN(II30536), .A(g23081) );
  INV_X1 NOT_8661( .ZN(g23492), .A(II30536) );
  INV_X1 NOT_8662( .ZN(g23493), .A(g22203) );
  INV_X1 NOT_8663( .ZN(II30544), .A(g23092) );
  INV_X1 NOT_8664( .ZN(g23500), .A(II30544) );
  INV_X1 NOT_8665( .ZN(II30547), .A(g23093) );
  INV_X1 NOT_8666( .ZN(g23501), .A(II30547) );
  INV_X1 NOT_8667( .ZN(II30552), .A(g23097) );
  INV_X1 NOT_8668( .ZN(g23508), .A(II30552) );
  INV_X1 NOT_8669( .ZN(g23509), .A(g22209) );
  INV_X1 NOT_8670( .ZN(II30560), .A(g23110) );
  INV_X1 NOT_8671( .ZN(g23516), .A(II30560) );
  INV_X1 NOT_8672( .ZN(II30563), .A(g23111) );
  INV_X1 NOT_8673( .ZN(g23517), .A(II30563) );
  INV_X1 NOT_8674( .ZN(II30568), .A(g23114) );
  INV_X1 NOT_8675( .ZN(g23524), .A(II30568) );
  INV_X1 NOT_8676( .ZN(II30575), .A(g23123) );
  INV_X1 NOT_8677( .ZN(g23531), .A(II30575) );
  INV_X1 NOT_8678( .ZN(II30578), .A(g23124) );
  INV_X1 NOT_8679( .ZN(g23532), .A(II30578) );
  INV_X1 NOT_8680( .ZN(II30586), .A(g23132) );
  INV_X1 NOT_8681( .ZN(g23542), .A(II30586) );
  INV_X1 NOT_8682( .ZN(II30589), .A(g23133) );
  INV_X1 NOT_8683( .ZN(g23543), .A(II30589) );
  INV_X1 NOT_8684( .ZN(II30594), .A(g22025) );
  INV_X1 NOT_8685( .ZN(g23546), .A(II30594) );
  INV_X1 NOT_8686( .ZN(II30598), .A(g22027) );
  INV_X1 NOT_8687( .ZN(g23548), .A(II30598) );
  INV_X1 NOT_8688( .ZN(II30601), .A(g22028) );
  INV_X1 NOT_8689( .ZN(g23549), .A(II30601) );
  INV_X1 NOT_8690( .ZN(II30607), .A(g22029) );
  INV_X1 NOT_8691( .ZN(g23553), .A(II30607) );
  INV_X1 NOT_8692( .ZN(II30611), .A(g22030) );
  INV_X1 NOT_8693( .ZN(g23555), .A(II30611) );
  INV_X1 NOT_8694( .ZN(II30614), .A(g22031) );
  INV_X1 NOT_8695( .ZN(g23556), .A(II30614) );
  INV_X1 NOT_8696( .ZN(II30617), .A(g22032) );
  INV_X1 NOT_8697( .ZN(g23557), .A(II30617) );
  INV_X1 NOT_8698( .ZN(II30623), .A(g22033) );
  INV_X1 NOT_8699( .ZN(g23561), .A(II30623) );
  INV_X1 NOT_8700( .ZN(II30626), .A(g22034) );
  INV_X1 NOT_8701( .ZN(g23562), .A(II30626) );
  INV_X1 NOT_8702( .ZN(II30632), .A(g22035) );
  INV_X1 NOT_8703( .ZN(g23566), .A(II30632) );
  INV_X1 NOT_8704( .ZN(II30636), .A(g22037) );
  INV_X1 NOT_8705( .ZN(g23568), .A(II30636) );
  INV_X1 NOT_8706( .ZN(II30639), .A(g22038) );
  INV_X1 NOT_8707( .ZN(g23569), .A(II30639) );
  INV_X1 NOT_8708( .ZN(II30642), .A(g22039) );
  INV_X1 NOT_8709( .ZN(g23570), .A(II30642) );
  INV_X1 NOT_8710( .ZN(II30648), .A(g22040) );
  INV_X1 NOT_8711( .ZN(g23574), .A(II30648) );
  INV_X1 NOT_8712( .ZN(II30651), .A(g22041) );
  INV_X1 NOT_8713( .ZN(g23575), .A(II30651) );
  INV_X1 NOT_8714( .ZN(II30654), .A(g22042) );
  INV_X1 NOT_8715( .ZN(g23576), .A(II30654) );
  INV_X1 NOT_8716( .ZN(II30660), .A(g22043) );
  INV_X1 NOT_8717( .ZN(g23580), .A(II30660) );
  INV_X1 NOT_8718( .ZN(II30663), .A(g22044) );
  INV_X1 NOT_8719( .ZN(g23581), .A(II30663) );
  INV_X1 NOT_8720( .ZN(II30669), .A(g22045) );
  INV_X1 NOT_8721( .ZN(g23585), .A(II30669) );
  INV_X1 NOT_8722( .ZN(II30673), .A(g22047) );
  INV_X1 NOT_8723( .ZN(g23587), .A(II30673) );
  INV_X1 NOT_8724( .ZN(II30676), .A(g22048) );
  INV_X1 NOT_8725( .ZN(g23588), .A(II30676) );
  INV_X1 NOT_8726( .ZN(II30679), .A(g22049) );
  INV_X1 NOT_8727( .ZN(g23589), .A(II30679) );
  INV_X1 NOT_8728( .ZN(II30686), .A(g23136) );
  INV_X8 NOT_8729( .ZN(g23594), .A(II30686) );
  INV_X8 NOT_8730( .ZN(II30689), .A(g22054) );
  INV_X1 NOT_8731( .ZN(g23595), .A(II30689) );
  INV_X1 NOT_8732( .ZN(II30692), .A(g22055) );
  INV_X1 NOT_8733( .ZN(g23596), .A(II30692) );
  INV_X1 NOT_8734( .ZN(II30695), .A(g22056) );
  INV_X1 NOT_8735( .ZN(g23597), .A(II30695) );
  INV_X1 NOT_8736( .ZN(II30701), .A(g22057) );
  INV_X1 NOT_8737( .ZN(g23601), .A(II30701) );
  INV_X1 NOT_8738( .ZN(II30704), .A(g22058) );
  INV_X1 NOT_8739( .ZN(g23602), .A(II30704) );
  INV_X1 NOT_8740( .ZN(II30707), .A(g22059) );
  INV_X1 NOT_8741( .ZN(g23603), .A(II30707) );
  INV_X1 NOT_8742( .ZN(II30713), .A(g22060) );
  INV_X1 NOT_8743( .ZN(g23607), .A(II30713) );
  INV_X1 NOT_8744( .ZN(II30716), .A(g22061) );
  INV_X1 NOT_8745( .ZN(g23608), .A(II30716) );
  INV_X1 NOT_8746( .ZN(II30722), .A(g22063) );
  INV_X1 NOT_8747( .ZN(g23612), .A(II30722) );
  INV_X1 NOT_8748( .ZN(II30725), .A(g22064) );
  INV_X1 NOT_8749( .ZN(g23613), .A(II30725) );
  INV_X1 NOT_8750( .ZN(II30728), .A(g22065) );
  INV_X1 NOT_8751( .ZN(g23614), .A(II30728) );
  INV_X1 NOT_8752( .ZN(II30735), .A(g22066) );
  INV_X1 NOT_8753( .ZN(g23619), .A(II30735) );
  INV_X1 NOT_8754( .ZN(II30738), .A(g22067) );
  INV_X1 NOT_8755( .ZN(g23620), .A(II30738) );
  INV_X1 NOT_8756( .ZN(II30741), .A(g22068) );
  INV_X1 NOT_8757( .ZN(g23621), .A(II30741) );
  INV_X1 NOT_8758( .ZN(II30748), .A(g21969) );
  INV_X1 NOT_8759( .ZN(g23626), .A(II30748) );
  INV_X1 NOT_8760( .ZN(II30751), .A(g22073) );
  INV_X1 NOT_8761( .ZN(g23627), .A(II30751) );
  INV_X1 NOT_8762( .ZN(II30754), .A(g22074) );
  INV_X1 NOT_8763( .ZN(g23628), .A(II30754) );
  INV_X1 NOT_8764( .ZN(II30757), .A(g22075) );
  INV_X1 NOT_8765( .ZN(g23629), .A(II30757) );
  INV_X1 NOT_8766( .ZN(II30763), .A(g22076) );
  INV_X1 NOT_8767( .ZN(g23633), .A(II30763) );
  INV_X1 NOT_8768( .ZN(II30766), .A(g22077) );
  INV_X1 NOT_8769( .ZN(g23634), .A(II30766) );
  INV_X1 NOT_8770( .ZN(II30769), .A(g22078) );
  INV_X1 NOT_8771( .ZN(g23635), .A(II30769) );
  INV_X1 NOT_8772( .ZN(II30776), .A(g22079) );
  INV_X1 NOT_8773( .ZN(g23640), .A(II30776) );
  INV_X1 NOT_8774( .ZN(II30779), .A(g22080) );
  INV_X1 NOT_8775( .ZN(g23641), .A(II30779) );
  INV_X1 NOT_8776( .ZN(II30782), .A(g22081) );
  INV_X1 NOT_8777( .ZN(g23642), .A(II30782) );
  INV_X1 NOT_8778( .ZN(II30786), .A(g22454) );
  INV_X1 NOT_8779( .ZN(g23644), .A(II30786) );
  INV_X1 NOT_8780( .ZN(II30797), .A(g22087) );
  INV_X1 NOT_8781( .ZN(g23661), .A(II30797) );
  INV_X1 NOT_8782( .ZN(II30800), .A(g22088) );
  INV_X1 NOT_8783( .ZN(g23662), .A(II30800) );
  INV_X1 NOT_8784( .ZN(II30803), .A(g22089) );
  INV_X1 NOT_8785( .ZN(g23663), .A(II30803) );
  INV_X1 NOT_8786( .ZN(II30810), .A(g22090) );
  INV_X1 NOT_8787( .ZN(g23668), .A(II30810) );
  INV_X1 NOT_8788( .ZN(II30813), .A(g22091) );
  INV_X1 NOT_8789( .ZN(g23669), .A(II30813) );
  INV_X1 NOT_8790( .ZN(II30816), .A(g22092) );
  INV_X1 NOT_8791( .ZN(g23670), .A(II30816) );
  INV_X1 NOT_8792( .ZN(II30823), .A(g21972) );
  INV_X1 NOT_8793( .ZN(g23675), .A(II30823) );
  INV_X1 NOT_8794( .ZN(II30826), .A(g22097) );
  INV_X1 NOT_8795( .ZN(g23676), .A(II30826) );
  INV_X1 NOT_8796( .ZN(II30829), .A(g22098) );
  INV_X1 NOT_8797( .ZN(g23677), .A(II30829) );
  INV_X1 NOT_8798( .ZN(II30832), .A(g22099) );
  INV_X1 NOT_8799( .ZN(g23678), .A(II30832) );
  INV_X1 NOT_8800( .ZN(II30838), .A(g22100) );
  INV_X1 NOT_8801( .ZN(g23682), .A(II30838) );
  INV_X1 NOT_8802( .ZN(II30841), .A(g22101) );
  INV_X1 NOT_8803( .ZN(g23683), .A(II30841) );
  INV_X1 NOT_8804( .ZN(II30844), .A(g22102) );
  INV_X1 NOT_8805( .ZN(g23684), .A(II30844) );
  INV_X1 NOT_8806( .ZN(II30847), .A(g22103) );
  INV_X1 NOT_8807( .ZN(g23685), .A(II30847) );
  INV_X1 NOT_8808( .ZN(II30854), .A(g22104) );
  INV_X1 NOT_8809( .ZN(g23690), .A(II30854) );
  INV_X1 NOT_8810( .ZN(II30857), .A(g22105) );
  INV_X1 NOT_8811( .ZN(g23691), .A(II30857) );
  INV_X1 NOT_8812( .ZN(II30860), .A(g22106) );
  INV_X1 NOT_8813( .ZN(g23692), .A(II30860) );
  INV_X1 NOT_8814( .ZN(II30864), .A(g22493) );
  INV_X1 NOT_8815( .ZN(g23694), .A(II30864) );
  INV_X1 NOT_8816( .ZN(II30875), .A(g22112) );
  INV_X1 NOT_8817( .ZN(g23711), .A(II30875) );
  INV_X1 NOT_8818( .ZN(II30878), .A(g22113) );
  INV_X1 NOT_8819( .ZN(g23712), .A(II30878) );
  INV_X1 NOT_8820( .ZN(II30881), .A(g22114) );
  INV_X1 NOT_8821( .ZN(g23713), .A(II30881) );
  INV_X1 NOT_8822( .ZN(II30888), .A(g22115) );
  INV_X1 NOT_8823( .ZN(g23718), .A(II30888) );
  INV_X1 NOT_8824( .ZN(II30891), .A(g22116) );
  INV_X1 NOT_8825( .ZN(g23719), .A(II30891) );
  INV_X1 NOT_8826( .ZN(II30894), .A(g22117) );
  INV_X1 NOT_8827( .ZN(g23720), .A(II30894) );
  INV_X1 NOT_8828( .ZN(II30901), .A(g21974) );
  INV_X1 NOT_8829( .ZN(g23725), .A(II30901) );
  INV_X1 NOT_8830( .ZN(II30905), .A(g22122) );
  INV_X1 NOT_8831( .ZN(g23727), .A(II30905) );
  INV_X1 NOT_8832( .ZN(II30908), .A(g22123) );
  INV_X1 NOT_8833( .ZN(g23728), .A(II30908) );
  INV_X1 NOT_8834( .ZN(II30911), .A(g22124) );
  INV_X1 NOT_8835( .ZN(g23729), .A(II30911) );
  INV_X1 NOT_8836( .ZN(II30914), .A(g22125) );
  INV_X1 NOT_8837( .ZN(g23730), .A(II30914) );
  INV_X1 NOT_8838( .ZN(II30917), .A(g22806) );
  INV_X1 NOT_8839( .ZN(g23731), .A(II30917) );
  INV_X1 NOT_8840( .ZN(II30922), .A(g22126) );
  INV_X1 NOT_8841( .ZN(g23736), .A(II30922) );
  INV_X1 NOT_8842( .ZN(II30925), .A(g22127) );
  INV_X1 NOT_8843( .ZN(g23737), .A(II30925) );
  INV_X1 NOT_8844( .ZN(II30928), .A(g22128) );
  INV_X1 NOT_8845( .ZN(g23738), .A(II30928) );
  INV_X1 NOT_8846( .ZN(II30931), .A(g22129) );
  INV_X1 NOT_8847( .ZN(g23739), .A(II30931) );
  INV_X1 NOT_8848( .ZN(II30938), .A(g22130) );
  INV_X1 NOT_8849( .ZN(g23744), .A(II30938) );
  INV_X1 NOT_8850( .ZN(II30941), .A(g22131) );
  INV_X1 NOT_8851( .ZN(g23745), .A(II30941) );
  INV_X1 NOT_8852( .ZN(II30944), .A(g22132) );
  INV_X1 NOT_8853( .ZN(g23746), .A(II30944) );
  INV_X1 NOT_8854( .ZN(II30948), .A(g22536) );
  INV_X1 NOT_8855( .ZN(g23748), .A(II30948) );
  INV_X1 NOT_8856( .ZN(II30959), .A(g22138) );
  INV_X1 NOT_8857( .ZN(g23765), .A(II30959) );
  INV_X1 NOT_8858( .ZN(II30962), .A(g22139) );
  INV_X1 NOT_8859( .ZN(g23766), .A(II30962) );
  INV_X1 NOT_8860( .ZN(II30965), .A(g22140) );
  INV_X1 NOT_8861( .ZN(g23767), .A(II30965) );
  INV_X1 NOT_8862( .ZN(II30973), .A(g22141) );
  INV_X1 NOT_8863( .ZN(g23773), .A(II30973) );
  INV_X1 NOT_8864( .ZN(II30976), .A(g22142) );
  INV_X1 NOT_8865( .ZN(g23774), .A(II30976) );
  INV_X1 NOT_8866( .ZN(II30979), .A(g22143) );
  INV_X1 NOT_8867( .ZN(g23775), .A(II30979) );
  INV_X1 NOT_8868( .ZN(II30985), .A(g22992) );
  INV_X1 NOT_8869( .ZN(g23779), .A(II30985) );
  INV_X1 NOT_8870( .ZN(II30988), .A(g22145) );
  INV_X1 NOT_8871( .ZN(g23782), .A(II30988) );
  INV_X1 NOT_8872( .ZN(II30991), .A(g22146) );
  INV_X1 NOT_8873( .ZN(g23783), .A(II30991) );
  INV_X1 NOT_8874( .ZN(II30994), .A(g22147) );
  INV_X1 NOT_8875( .ZN(g23784), .A(II30994) );
  INV_X1 NOT_8876( .ZN(II30997), .A(g22148) );
  INV_X1 NOT_8877( .ZN(g23785), .A(II30997) );
  INV_X1 NOT_8878( .ZN(II31000), .A(g22847) );
  INV_X1 NOT_8879( .ZN(g23786), .A(II31000) );
  INV_X1 NOT_8880( .ZN(II31005), .A(g22149) );
  INV_X1 NOT_8881( .ZN(g23791), .A(II31005) );
  INV_X1 NOT_8882( .ZN(II31008), .A(g22150) );
  INV_X1 NOT_8883( .ZN(g23792), .A(II31008) );
  INV_X1 NOT_8884( .ZN(II31011), .A(g22151) );
  INV_X1 NOT_8885( .ZN(g23793), .A(II31011) );
  INV_X1 NOT_8886( .ZN(II31014), .A(g22152) );
  INV_X1 NOT_8887( .ZN(g23794), .A(II31014) );
  INV_X1 NOT_8888( .ZN(II31021), .A(g22153) );
  INV_X1 NOT_8889( .ZN(g23799), .A(II31021) );
  INV_X1 NOT_8890( .ZN(II31024), .A(g22154) );
  INV_X1 NOT_8891( .ZN(g23800), .A(II31024) );
  INV_X1 NOT_8892( .ZN(II31027), .A(g22155) );
  INV_X1 NOT_8893( .ZN(g23801), .A(II31027) );
  INV_X1 NOT_8894( .ZN(II31031), .A(g22576) );
  INV_X1 NOT_8895( .ZN(g23803), .A(II31031) );
  INV_X1 NOT_8896( .ZN(II31043), .A(g22161) );
  INV_X1 NOT_8897( .ZN(g23821), .A(II31043) );
  INV_X1 NOT_8898( .ZN(II31050), .A(g22162) );
  INV_X1 NOT_8899( .ZN(g23826), .A(II31050) );
  INV_X1 NOT_8900( .ZN(II31053), .A(g22163) );
  INV_X1 NOT_8901( .ZN(g23827), .A(II31053) );
  INV_X1 NOT_8902( .ZN(II31056), .A(g22164) );
  INV_X1 NOT_8903( .ZN(g23828), .A(II31056) );
  INV_X1 NOT_8904( .ZN(II31062), .A(g23003) );
  INV_X1 NOT_8905( .ZN(g23832), .A(II31062) );
  INV_X1 NOT_8906( .ZN(II31065), .A(g22166) );
  INV_X1 NOT_8907( .ZN(g23835), .A(II31065) );
  INV_X1 NOT_8908( .ZN(II31068), .A(g22167) );
  INV_X1 NOT_8909( .ZN(g23836), .A(II31068) );
  INV_X1 NOT_8910( .ZN(II31071), .A(g22168) );
  INV_X1 NOT_8911( .ZN(g23837), .A(II31071) );
  INV_X1 NOT_8912( .ZN(II31074), .A(g22169) );
  INV_X1 NOT_8913( .ZN(g23838), .A(II31074) );
  INV_X1 NOT_8914( .ZN(II31077), .A(g22882) );
  INV_X1 NOT_8915( .ZN(g23839), .A(II31077) );
  INV_X1 NOT_8916( .ZN(II31082), .A(g22170) );
  INV_X1 NOT_8917( .ZN(g23844), .A(II31082) );
  INV_X1 NOT_8918( .ZN(II31085), .A(g22171) );
  INV_X1 NOT_8919( .ZN(g23845), .A(II31085) );
  INV_X1 NOT_8920( .ZN(II31088), .A(g22172) );
  INV_X1 NOT_8921( .ZN(g23846), .A(II31088) );
  INV_X1 NOT_8922( .ZN(II31091), .A(g22173) );
  INV_X1 NOT_8923( .ZN(g23847), .A(II31091) );
  INV_X1 NOT_8924( .ZN(g23853), .A(g22300) );
  INV_X1 NOT_8925( .ZN(II31102), .A(g22177) );
  INV_X1 NOT_8926( .ZN(g23856), .A(II31102) );
  INV_X1 NOT_8927( .ZN(II31109), .A(g22178) );
  INV_X1 NOT_8928( .ZN(g23861), .A(II31109) );
  INV_X1 NOT_8929( .ZN(II31112), .A(g22179) );
  INV_X1 NOT_8930( .ZN(g23862), .A(II31112) );
  INV_X1 NOT_8931( .ZN(II31115), .A(g22180) );
  INV_X1 NOT_8932( .ZN(g23863), .A(II31115) );
  INV_X1 NOT_8933( .ZN(II31121), .A(g23017) );
  INV_X1 NOT_8934( .ZN(g23867), .A(II31121) );
  INV_X1 NOT_8935( .ZN(II31124), .A(g22182) );
  INV_X1 NOT_8936( .ZN(g23870), .A(II31124) );
  INV_X1 NOT_8937( .ZN(II31127), .A(g22183) );
  INV_X1 NOT_8938( .ZN(g23871), .A(II31127) );
  INV_X1 NOT_8939( .ZN(II31130), .A(g22184) );
  INV_X1 NOT_8940( .ZN(g23872), .A(II31130) );
  INV_X1 NOT_8941( .ZN(II31133), .A(g22185) );
  INV_X1 NOT_8942( .ZN(g23873), .A(II31133) );
  INV_X1 NOT_8943( .ZN(II31136), .A(g22917) );
  INV_X1 NOT_8944( .ZN(g23874), .A(II31136) );
  INV_X1 NOT_8945( .ZN(II31141), .A(g22777) );
  INV_X1 NOT_8946( .ZN(g23879), .A(II31141) );
  INV_X1 NOT_8947( .ZN(II31144), .A(g22935) );
  INV_X1 NOT_8948( .ZN(g23882), .A(II31144) );
  INV_X1 NOT_8949( .ZN(g23885), .A(g22062) );
  INV_X1 NOT_8950( .ZN(g23887), .A(g22328) );
  INV_X1 NOT_8951( .ZN(II31152), .A(g22191) );
  INV_X1 NOT_8952( .ZN(g23890), .A(II31152) );
  INV_X1 NOT_8953( .ZN(II31159), .A(g22192) );
  INV_X1 NOT_8954( .ZN(g23895), .A(II31159) );
  INV_X1 NOT_8955( .ZN(II31162), .A(g22193) );
  INV_X1 NOT_8956( .ZN(g23896), .A(II31162) );
  INV_X1 NOT_8957( .ZN(II31165), .A(g22194) );
  INV_X8 NOT_8958( .ZN(g23897), .A(II31165) );
  INV_X1 NOT_8959( .ZN(II31171), .A(g23033) );
  INV_X1 NOT_8960( .ZN(g23901), .A(II31171) );
  INV_X1 NOT_8961( .ZN(g23905), .A(g22046) );
  INV_X1 NOT_8962( .ZN(g23908), .A(g22353) );
  INV_X1 NOT_8963( .ZN(II31181), .A(g22200) );
  INV_X1 NOT_8964( .ZN(g23911), .A(II31181) );
  INV_X1 NOT_8965( .ZN(II31188), .A(g21989) );
  INV_X1 NOT_8966( .ZN(g23916), .A(II31188) );
  INV_X1 NOT_8967( .ZN(g23918), .A(g22036) );
  INV_X1 NOT_8968( .ZN(II31195), .A(g22578) );
  INV_X1 NOT_8969( .ZN(g23923), .A(II31195) );
  INV_X1 NOT_8970( .ZN(g23940), .A(g22376) );
  INV_X1 NOT_8971( .ZN(II31205), .A(g22002) );
  INV_X1 NOT_8972( .ZN(g23943), .A(II31205) );
  INV_X1 NOT_8973( .ZN(II31213), .A(g22615) );
  INV_X1 NOT_8974( .ZN(g23955), .A(II31213) );
  INV_X1 NOT_8975( .ZN(II31226), .A(g22651) );
  INV_X1 NOT_8976( .ZN(g23984), .A(II31226) );
  INV_X1 NOT_8977( .ZN(II31232), .A(g22026) );
  INV_X1 NOT_8978( .ZN(g24000), .A(II31232) );
  INV_X1 NOT_8979( .ZN(II31235), .A(g22218) );
  INV_X1 NOT_8980( .ZN(g24001), .A(II31235) );
  INV_X1 NOT_8981( .ZN(II31244), .A(g22687) );
  INV_X1 NOT_8982( .ZN(g24014), .A(II31244) );
  INV_X1 NOT_8983( .ZN(II31250), .A(g22953) );
  INV_X1 NOT_8984( .ZN(g24030), .A(II31250) );
  INV_X1 NOT_8985( .ZN(II31253), .A(g22231) );
  INV_X1 NOT_8986( .ZN(g24033), .A(II31253) );
  INV_X1 NOT_8987( .ZN(II31257), .A(g22234) );
  INV_X1 NOT_8988( .ZN(g24035), .A(II31257) );
  INV_X1 NOT_8989( .ZN(g24047), .A(g23023) );
  INV_X1 NOT_8990( .ZN(II31266), .A(g22242) );
  INV_X1 NOT_8991( .ZN(g24051), .A(II31266) );
  INV_X1 NOT_8992( .ZN(II31270), .A(g22247) );
  INV_X1 NOT_8993( .ZN(g24053), .A(II31270) );
  INV_X1 NOT_8994( .ZN(II31274), .A(g22249) );
  INV_X1 NOT_8995( .ZN(g24055), .A(II31274) );
  INV_X1 NOT_8996( .ZN(g24060), .A(g23040) );
  INV_X1 NOT_8997( .ZN(II31282), .A(g22263) );
  INV_X1 NOT_8998( .ZN(g24064), .A(II31282) );
  INV_X1 NOT_8999( .ZN(II31286), .A(g22267) );
  INV_X1 NOT_9000( .ZN(g24066), .A(II31286) );
  INV_X1 NOT_9001( .ZN(II31290), .A(g22269) );
  INV_X1 NOT_9002( .ZN(g24068), .A(II31290) );
  INV_X1 NOT_9003( .ZN(g24073), .A(g23059) );
  INV_X1 NOT_9004( .ZN(II31298), .A(g22280) );
  INV_X1 NOT_9005( .ZN(g24077), .A(II31298) );
  INV_X1 NOT_9006( .ZN(II31302), .A(g22284) );
  INV_X1 NOT_9007( .ZN(g24079), .A(II31302) );
  INV_X1 NOT_9008( .ZN(g24084), .A(g23077) );
  INV_X1 NOT_9009( .ZN(II31310), .A(g22299) );
  INV_X1 NOT_9010( .ZN(g24088), .A(II31310) );
  INV_X1 NOT_9011( .ZN(g24094), .A(g22339) );
  INV_X1 NOT_9012( .ZN(g24095), .A(g22362) );
  INV_X1 NOT_9013( .ZN(g24096), .A(g22405) );
  INV_X1 NOT_9014( .ZN(g24097), .A(g22382) );
  INV_X1 NOT_9015( .ZN(g24098), .A(g22409) );
  INV_X1 NOT_9016( .ZN(g24099), .A(g22412) );
  INV_X1 NOT_9017( .ZN(g24101), .A(g22415) );
  INV_X1 NOT_9018( .ZN(g24102), .A(g22418) );
  INV_X1 NOT_9019( .ZN(g24103), .A(g22397) );
  INV_X1 NOT_9020( .ZN(g24104), .A(g22422) );
  INV_X1 NOT_9021( .ZN(g24105), .A(g22425) );
  INV_X1 NOT_9022( .ZN(g24106), .A(g22428) );
  INV_X1 NOT_9023( .ZN(g24107), .A(g22431) );
  INV_X1 NOT_9024( .ZN(g24108), .A(g22434) );
  INV_X1 NOT_9025( .ZN(g24110), .A(g22437) );
  INV_X1 NOT_9026( .ZN(g24111), .A(g22440) );
  INV_X1 NOT_9027( .ZN(g24112), .A(g22445) );
  INV_X1 NOT_9028( .ZN(g24113), .A(g22448) );
  INV_X1 NOT_9029( .ZN(g24114), .A(g22451) );
  INV_X1 NOT_9030( .ZN(g24115), .A(g22381) );
  INV_X1 NOT_9031( .ZN(g24121), .A(g22455) );
  INV_X1 NOT_9032( .ZN(g24122), .A(g22458) );
  INV_X1 NOT_9033( .ZN(g24123), .A(g22461) );
  INV_X1 NOT_9034( .ZN(g24124), .A(g22464) );
  INV_X1 NOT_9035( .ZN(g24125), .A(g22467) );
  INV_X1 NOT_9036( .ZN(g24127), .A(g22470) );
  INV_X1 NOT_9037( .ZN(g24128), .A(g22473) );
  INV_X1 NOT_9038( .ZN(g24129), .A(g22477) );
  INV_X1 NOT_9039( .ZN(g24130), .A(g22480) );
  INV_X1 NOT_9040( .ZN(g24131), .A(g22484) );
  INV_X1 NOT_9041( .ZN(g24132), .A(g22487) );
  INV_X1 NOT_9042( .ZN(g24133), .A(g22490) );
  INV_X1 NOT_9043( .ZN(g24134), .A(g22396) );
  INV_X1 NOT_9044( .ZN(g24140), .A(g22494) );
  INV_X1 NOT_9045( .ZN(g24141), .A(g22497) );
  INV_X1 NOT_9046( .ZN(g24142), .A(g22500) );
  INV_X1 NOT_9047( .ZN(g24143), .A(g22503) );
  INV_X1 NOT_9048( .ZN(g24144), .A(g22506) );
  INV_X1 NOT_9049( .ZN(g24146), .A(g22509) );
  INV_X1 NOT_9050( .ZN(g24147), .A(g22512) );
  INV_X1 NOT_9051( .ZN(g24148), .A(g22520) );
  INV_X1 NOT_9052( .ZN(g24149), .A(g22523) );
  INV_X1 NOT_9053( .ZN(g24150), .A(g22527) );
  INV_X1 NOT_9054( .ZN(g24151), .A(g22530) );
  INV_X1 NOT_9055( .ZN(g24152), .A(g22533) );
  INV_X1 NOT_9056( .ZN(g24153), .A(g22399) );
  INV_X1 NOT_9057( .ZN(g24159), .A(g22537) );
  INV_X1 NOT_9058( .ZN(g24160), .A(g22540) );
  INV_X1 NOT_9059( .ZN(g24161), .A(g22543) );
  INV_X1 NOT_9060( .ZN(g24162), .A(g22552) );
  INV_X1 NOT_9061( .ZN(g24163), .A(g22560) );
  INV_X1 NOT_9062( .ZN(g24164), .A(g22563) );
  INV_X1 NOT_9063( .ZN(g24165), .A(g22567) );
  INV_X1 NOT_9064( .ZN(g24166), .A(g22570) );
  INV_X1 NOT_9065( .ZN(g24167), .A(g22573) );
  INV_X1 NOT_9066( .ZN(g24168), .A(g22400) );
  INV_X1 NOT_9067( .ZN(g24175), .A(g22592) );
  INV_X1 NOT_9068( .ZN(g24176), .A(g22600) );
  INV_X1 NOT_9069( .ZN(g24177), .A(g22603) );
  INV_X1 NOT_9070( .ZN(g24180), .A(g22629) );
  INV_X1 NOT_9071( .ZN(II31387), .A(g22811) );
  INV_X1 NOT_9072( .ZN(g24183), .A(II31387) );
  INV_X1 NOT_9073( .ZN(g24210), .A(g22696) );
  INV_X1 NOT_9074( .ZN(g24220), .A(g22750) );
  INV_X1 NOT_9075( .ZN(II31417), .A(g22578) );
  INV_X1 NOT_9076( .ZN(g24233), .A(II31417) );
  INV_X1 NOT_9077( .ZN(II31426), .A(g22615) );
  INV_X1 NOT_9078( .ZN(g24240), .A(II31426) );
  INV_X1 NOT_9079( .ZN(II31436), .A(g22651) );
  INV_X1 NOT_9080( .ZN(g24248), .A(II31436) );
  INV_X1 NOT_9081( .ZN(g24251), .A(g22903) );
  INV_X1 NOT_9082( .ZN(II31445), .A(g22687) );
  INV_X1 NOT_9083( .ZN(g24255), .A(II31445) );
  INV_X1 NOT_9084( .ZN(II31451), .A(g23682) );
  INV_X1 NOT_9085( .ZN(g24259), .A(II31451) );
  INV_X1 NOT_9086( .ZN(II31454), .A(g23727) );
  INV_X1 NOT_9087( .ZN(g24260), .A(II31454) );
  INV_X1 NOT_9088( .ZN(II31457), .A(g23773) );
  INV_X1 NOT_9089( .ZN(g24261), .A(II31457) );
  INV_X1 NOT_9090( .ZN(II31460), .A(g23728) );
  INV_X1 NOT_9091( .ZN(g24262), .A(II31460) );
  INV_X1 NOT_9092( .ZN(II31463), .A(g23774) );
  INV_X1 NOT_9093( .ZN(g24263), .A(II31463) );
  INV_X1 NOT_9094( .ZN(II31466), .A(g23821) );
  INV_X1 NOT_9095( .ZN(g24264), .A(II31466) );
  INV_X1 NOT_9096( .ZN(II31469), .A(g23546) );
  INV_X1 NOT_9097( .ZN(g24265), .A(II31469) );
  INV_X1 NOT_9098( .ZN(II31472), .A(g23548) );
  INV_X1 NOT_9099( .ZN(g24266), .A(II31472) );
  INV_X1 NOT_9100( .ZN(II31475), .A(g23555) );
  INV_X1 NOT_9101( .ZN(g24267), .A(II31475) );
  INV_X1 NOT_9102( .ZN(II31478), .A(g23549) );
  INV_X1 NOT_9103( .ZN(g24268), .A(II31478) );
  INV_X1 NOT_9104( .ZN(II31481), .A(g23556) );
  INV_X1 NOT_9105( .ZN(g24269), .A(II31481) );
  INV_X1 NOT_9106( .ZN(II31484), .A(g23568) );
  INV_X1 NOT_9107( .ZN(g24270), .A(II31484) );
  INV_X1 NOT_9108( .ZN(II31487), .A(g23557) );
  INV_X1 NOT_9109( .ZN(g24271), .A(II31487) );
  INV_X1 NOT_9110( .ZN(II31490), .A(g23569) );
  INV_X1 NOT_9111( .ZN(g24272), .A(II31490) );
  INV_X1 NOT_9112( .ZN(II31493), .A(g23587) );
  INV_X1 NOT_9113( .ZN(g24273), .A(II31493) );
  INV_X1 NOT_9114( .ZN(II31496), .A(g23570) );
  INV_X1 NOT_9115( .ZN(g24274), .A(II31496) );
  INV_X1 NOT_9116( .ZN(II31499), .A(g23588) );
  INV_X1 NOT_9117( .ZN(g24275), .A(II31499) );
  INV_X1 NOT_9118( .ZN(II31502), .A(g23612) );
  INV_X1 NOT_9119( .ZN(g24276), .A(II31502) );
  INV_X1 NOT_9120( .ZN(II31505), .A(g23589) );
  INV_X1 NOT_9121( .ZN(g24277), .A(II31505) );
  INV_X1 NOT_9122( .ZN(II31508), .A(g23613) );
  INV_X1 NOT_9123( .ZN(g24278), .A(II31508) );
  INV_X1 NOT_9124( .ZN(II31511), .A(g23640) );
  INV_X1 NOT_9125( .ZN(g24279), .A(II31511) );
  INV_X1 NOT_9126( .ZN(II31514), .A(g23614) );
  INV_X1 NOT_9127( .ZN(g24280), .A(II31514) );
  INV_X1 NOT_9128( .ZN(II31517), .A(g23641) );
  INV_X1 NOT_9129( .ZN(g24281), .A(II31517) );
  INV_X1 NOT_9130( .ZN(II31520), .A(g23683) );
  INV_X1 NOT_9131( .ZN(g24282), .A(II31520) );
  INV_X1 NOT_9132( .ZN(II31523), .A(g23642) );
  INV_X8 NOT_9133( .ZN(g24283), .A(II31523) );
  INV_X8 NOT_9134( .ZN(II31526), .A(g23684) );
  INV_X8 NOT_9135( .ZN(g24284), .A(II31526) );
  INV_X1 NOT_9136( .ZN(II31529), .A(g23729) );
  INV_X1 NOT_9137( .ZN(g24285), .A(II31529) );
  INV_X1 NOT_9138( .ZN(II31532), .A(g23685) );
  INV_X1 NOT_9139( .ZN(g24286), .A(II31532) );
  INV_X1 NOT_9140( .ZN(II31535), .A(g23730) );
  INV_X1 NOT_9141( .ZN(g24287), .A(II31535) );
  INV_X1 NOT_9142( .ZN(II31538), .A(g23775) );
  INV_X1 NOT_9143( .ZN(g24288), .A(II31538) );
  INV_X1 NOT_9144( .ZN(II31541), .A(g23500) );
  INV_X1 NOT_9145( .ZN(g24289), .A(II31541) );
  INV_X1 NOT_9146( .ZN(II31544), .A(g23438) );
  INV_X1 NOT_9147( .ZN(g24290), .A(II31544) );
  INV_X1 NOT_9148( .ZN(II31547), .A(g23454) );
  INV_X1 NOT_9149( .ZN(g24291), .A(II31547) );
  INV_X1 NOT_9150( .ZN(II31550), .A(g23481) );
  INV_X1 NOT_9151( .ZN(g24292), .A(II31550) );
  INV_X1 NOT_9152( .ZN(II31553), .A(g23501) );
  INV_X1 NOT_9153( .ZN(g24293), .A(II31553) );
  INV_X1 NOT_9154( .ZN(II31556), .A(g23439) );
  INV_X1 NOT_9155( .ZN(g24294), .A(II31556) );
  INV_X1 NOT_9156( .ZN(II31559), .A(g24233) );
  INV_X1 NOT_9157( .ZN(g24295), .A(II31559) );
  INV_X1 NOT_9158( .ZN(II31562), .A(g23594) );
  INV_X1 NOT_9159( .ZN(g24296), .A(II31562) );
  INV_X1 NOT_9160( .ZN(II31565), .A(g24001) );
  INV_X1 NOT_9161( .ZN(g24297), .A(II31565) );
  INV_X1 NOT_9162( .ZN(II31568), .A(g24033) );
  INV_X1 NOT_9163( .ZN(g24298), .A(II31568) );
  INV_X1 NOT_9164( .ZN(II31571), .A(g24051) );
  INV_X1 NOT_9165( .ZN(g24299), .A(II31571) );
  INV_X1 NOT_9166( .ZN(II31574), .A(g23736) );
  INV_X1 NOT_9167( .ZN(g24300), .A(II31574) );
  INV_X1 NOT_9168( .ZN(II31577), .A(g23782) );
  INV_X1 NOT_9169( .ZN(g24301), .A(II31577) );
  INV_X1 NOT_9170( .ZN(II31580), .A(g23826) );
  INV_X1 NOT_9171( .ZN(g24302), .A(II31580) );
  INV_X1 NOT_9172( .ZN(II31583), .A(g23783) );
  INV_X1 NOT_9173( .ZN(g24303), .A(II31583) );
  INV_X1 NOT_9174( .ZN(II31586), .A(g23827) );
  INV_X1 NOT_9175( .ZN(g24304), .A(II31586) );
  INV_X1 NOT_9176( .ZN(II31589), .A(g23856) );
  INV_X1 NOT_9177( .ZN(g24305), .A(II31589) );
  INV_X1 NOT_9178( .ZN(II31592), .A(g23553) );
  INV_X1 NOT_9179( .ZN(g24306), .A(II31592) );
  INV_X1 NOT_9180( .ZN(II31595), .A(g23561) );
  INV_X1 NOT_9181( .ZN(g24307), .A(II31595) );
  INV_X1 NOT_9182( .ZN(II31598), .A(g23574) );
  INV_X1 NOT_9183( .ZN(g24308), .A(II31598) );
  INV_X1 NOT_9184( .ZN(II31601), .A(g23562) );
  INV_X1 NOT_9185( .ZN(g24309), .A(II31601) );
  INV_X1 NOT_9186( .ZN(II31604), .A(g23575) );
  INV_X1 NOT_9187( .ZN(g24310), .A(II31604) );
  INV_X1 NOT_9188( .ZN(II31607), .A(g23595) );
  INV_X1 NOT_9189( .ZN(g24311), .A(II31607) );
  INV_X1 NOT_9190( .ZN(II31610), .A(g23576) );
  INV_X1 NOT_9191( .ZN(g24312), .A(II31610) );
  INV_X1 NOT_9192( .ZN(II31613), .A(g23596) );
  INV_X1 NOT_9193( .ZN(g24313), .A(II31613) );
  INV_X1 NOT_9194( .ZN(II31616), .A(g23619) );
  INV_X1 NOT_9195( .ZN(g24314), .A(II31616) );
  INV_X1 NOT_9196( .ZN(II31619), .A(g23597) );
  INV_X1 NOT_9197( .ZN(g24315), .A(II31619) );
  INV_X1 NOT_9198( .ZN(II31622), .A(g23620) );
  INV_X1 NOT_9199( .ZN(g24316), .A(II31622) );
  INV_X1 NOT_9200( .ZN(II31625), .A(g23661) );
  INV_X1 NOT_9201( .ZN(g24317), .A(II31625) );
  INV_X1 NOT_9202( .ZN(II31628), .A(g23621) );
  INV_X1 NOT_9203( .ZN(g24318), .A(II31628) );
  INV_X1 NOT_9204( .ZN(II31631), .A(g23662) );
  INV_X1 NOT_9205( .ZN(g24319), .A(II31631) );
  INV_X1 NOT_9206( .ZN(II31634), .A(g23690) );
  INV_X1 NOT_9207( .ZN(g24320), .A(II31634) );
  INV_X1 NOT_9208( .ZN(II31637), .A(g23663) );
  INV_X1 NOT_9209( .ZN(g24321), .A(II31637) );
  INV_X1 NOT_9210( .ZN(II31640), .A(g23691) );
  INV_X1 NOT_9211( .ZN(g24322), .A(II31640) );
  INV_X1 NOT_9212( .ZN(II31643), .A(g23737) );
  INV_X1 NOT_9213( .ZN(g24323), .A(II31643) );
  INV_X1 NOT_9214( .ZN(II31646), .A(g23692) );
  INV_X1 NOT_9215( .ZN(g24324), .A(II31646) );
  INV_X1 NOT_9216( .ZN(II31649), .A(g23738) );
  INV_X1 NOT_9217( .ZN(g24325), .A(II31649) );
  INV_X1 NOT_9218( .ZN(II31652), .A(g23784) );
  INV_X1 NOT_9219( .ZN(g24326), .A(II31652) );
  INV_X1 NOT_9220( .ZN(II31655), .A(g23739) );
  INV_X1 NOT_9221( .ZN(g24327), .A(II31655) );
  INV_X1 NOT_9222( .ZN(II31658), .A(g23785) );
  INV_X1 NOT_9223( .ZN(g24328), .A(II31658) );
  INV_X1 NOT_9224( .ZN(II31661), .A(g23828) );
  INV_X1 NOT_9225( .ZN(g24329), .A(II31661) );
  INV_X1 NOT_9226( .ZN(II31664), .A(g23516) );
  INV_X1 NOT_9227( .ZN(g24330), .A(II31664) );
  INV_X1 NOT_9228( .ZN(II31667), .A(g23452) );
  INV_X1 NOT_9229( .ZN(g24331), .A(II31667) );
  INV_X1 NOT_9230( .ZN(II31670), .A(g23463) );
  INV_X1 NOT_9231( .ZN(g24332), .A(II31670) );
  INV_X1 NOT_9232( .ZN(II31673), .A(g23492) );
  INV_X1 NOT_9233( .ZN(g24333), .A(II31673) );
  INV_X1 NOT_9234( .ZN(II31676), .A(g23517) );
  INV_X1 NOT_9235( .ZN(g24334), .A(II31676) );
  INV_X1 NOT_9236( .ZN(II31679), .A(g23453) );
  INV_X1 NOT_9237( .ZN(g24335), .A(II31679) );
  INV_X1 NOT_9238( .ZN(II31682), .A(g24240) );
  INV_X1 NOT_9239( .ZN(g24336), .A(II31682) );
  INV_X1 NOT_9240( .ZN(II31685), .A(g23626) );
  INV_X1 NOT_9241( .ZN(g24337), .A(II31685) );
  INV_X1 NOT_9242( .ZN(II31688), .A(g24035) );
  INV_X1 NOT_9243( .ZN(g24338), .A(II31688) );
  INV_X1 NOT_9244( .ZN(II31691), .A(g24053) );
  INV_X1 NOT_9245( .ZN(g24339), .A(II31691) );
  INV_X1 NOT_9246( .ZN(II31694), .A(g24064) );
  INV_X1 NOT_9247( .ZN(g24340), .A(II31694) );
  INV_X1 NOT_9248( .ZN(II31697), .A(g23791) );
  INV_X1 NOT_9249( .ZN(g24341), .A(II31697) );
  INV_X1 NOT_9250( .ZN(II31700), .A(g23835) );
  INV_X1 NOT_9251( .ZN(g24342), .A(II31700) );
  INV_X1 NOT_9252( .ZN(II31703), .A(g23861) );
  INV_X1 NOT_9253( .ZN(g24343), .A(II31703) );
  INV_X1 NOT_9254( .ZN(II31706), .A(g23836) );
  INV_X1 NOT_9255( .ZN(g24344), .A(II31706) );
  INV_X1 NOT_9256( .ZN(II31709), .A(g23862) );
  INV_X1 NOT_9257( .ZN(g24345), .A(II31709) );
  INV_X1 NOT_9258( .ZN(II31712), .A(g23890) );
  INV_X1 NOT_9259( .ZN(g24346), .A(II31712) );
  INV_X1 NOT_9260( .ZN(II31715), .A(g23566) );
  INV_X1 NOT_9261( .ZN(g24347), .A(II31715) );
  INV_X1 NOT_9262( .ZN(II31718), .A(g23580) );
  INV_X1 NOT_9263( .ZN(g24348), .A(II31718) );
  INV_X1 NOT_9264( .ZN(II31721), .A(g23601) );
  INV_X1 NOT_9265( .ZN(g24349), .A(II31721) );
  INV_X1 NOT_9266( .ZN(II31724), .A(g23581) );
  INV_X1 NOT_9267( .ZN(g24350), .A(II31724) );
  INV_X1 NOT_9268( .ZN(II31727), .A(g23602) );
  INV_X1 NOT_9269( .ZN(g24351), .A(II31727) );
  INV_X1 NOT_9270( .ZN(II31730), .A(g23627) );
  INV_X1 NOT_9271( .ZN(g24352), .A(II31730) );
  INV_X1 NOT_9272( .ZN(II31733), .A(g23603) );
  INV_X1 NOT_9273( .ZN(g24353), .A(II31733) );
  INV_X1 NOT_9274( .ZN(II31736), .A(g23628) );
  INV_X1 NOT_9275( .ZN(g24354), .A(II31736) );
  INV_X1 NOT_9276( .ZN(II31739), .A(g23668) );
  INV_X1 NOT_9277( .ZN(g24355), .A(II31739) );
  INV_X1 NOT_9278( .ZN(II31742), .A(g23629) );
  INV_X1 NOT_9279( .ZN(g24356), .A(II31742) );
  INV_X1 NOT_9280( .ZN(II31745), .A(g23669) );
  INV_X1 NOT_9281( .ZN(g24357), .A(II31745) );
  INV_X1 NOT_9282( .ZN(II31748), .A(g23711) );
  INV_X1 NOT_9283( .ZN(g24358), .A(II31748) );
  INV_X1 NOT_9284( .ZN(II31751), .A(g23670) );
  INV_X1 NOT_9285( .ZN(g24359), .A(II31751) );
  INV_X1 NOT_9286( .ZN(II31754), .A(g23712) );
  INV_X1 NOT_9287( .ZN(g24360), .A(II31754) );
  INV_X1 NOT_9288( .ZN(II31757), .A(g23744) );
  INV_X1 NOT_9289( .ZN(g24361), .A(II31757) );
  INV_X1 NOT_9290( .ZN(II31760), .A(g23713) );
  INV_X1 NOT_9291( .ZN(g24362), .A(II31760) );
  INV_X1 NOT_9292( .ZN(II31763), .A(g23745) );
  INV_X1 NOT_9293( .ZN(g24363), .A(II31763) );
  INV_X1 NOT_9294( .ZN(II31766), .A(g23792) );
  INV_X1 NOT_9295( .ZN(g24364), .A(II31766) );
  INV_X1 NOT_9296( .ZN(II31769), .A(g23746) );
  INV_X1 NOT_9297( .ZN(g24365), .A(II31769) );
  INV_X1 NOT_9298( .ZN(II31772), .A(g23793) );
  INV_X1 NOT_9299( .ZN(g24366), .A(II31772) );
  INV_X1 NOT_9300( .ZN(II31775), .A(g23837) );
  INV_X1 NOT_9301( .ZN(g24367), .A(II31775) );
  INV_X1 NOT_9302( .ZN(II31778), .A(g23794) );
  INV_X1 NOT_9303( .ZN(g24368), .A(II31778) );
  INV_X1 NOT_9304( .ZN(II31781), .A(g23838) );
  INV_X1 NOT_9305( .ZN(g24369), .A(II31781) );
  INV_X1 NOT_9306( .ZN(II31784), .A(g23863) );
  INV_X1 NOT_9307( .ZN(g24370), .A(II31784) );
  INV_X1 NOT_9308( .ZN(II31787), .A(g23531) );
  INV_X1 NOT_9309( .ZN(g24371), .A(II31787) );
  INV_X8 NOT_9310( .ZN(II31790), .A(g23459) );
  INV_X1 NOT_9311( .ZN(g24372), .A(II31790) );
  INV_X1 NOT_9312( .ZN(II31793), .A(g23472) );
  INV_X1 NOT_9313( .ZN(g24373), .A(II31793) );
  INV_X1 NOT_9314( .ZN(II31796), .A(g23508) );
  INV_X1 NOT_9315( .ZN(g24374), .A(II31796) );
  INV_X1 NOT_9316( .ZN(II31799), .A(g23532) );
  INV_X1 NOT_9317( .ZN(g24375), .A(II31799) );
  INV_X1 NOT_9318( .ZN(II31802), .A(g23460) );
  INV_X1 NOT_9319( .ZN(g24376), .A(II31802) );
  INV_X1 NOT_9320( .ZN(II31805), .A(g24248) );
  INV_X1 NOT_9321( .ZN(g24377), .A(II31805) );
  INV_X1 NOT_9322( .ZN(II31808), .A(g23675) );
  INV_X1 NOT_9323( .ZN(g24378), .A(II31808) );
  INV_X1 NOT_9324( .ZN(II31811), .A(g24055) );
  INV_X1 NOT_9325( .ZN(g24379), .A(II31811) );
  INV_X1 NOT_9326( .ZN(II31814), .A(g24066) );
  INV_X1 NOT_9327( .ZN(g24380), .A(II31814) );
  INV_X1 NOT_9328( .ZN(II31817), .A(g24077) );
  INV_X1 NOT_9329( .ZN(g24381), .A(II31817) );
  INV_X1 NOT_9330( .ZN(II31820), .A(g23844) );
  INV_X1 NOT_9331( .ZN(g24382), .A(II31820) );
  INV_X1 NOT_9332( .ZN(II31823), .A(g23870) );
  INV_X1 NOT_9333( .ZN(g24383), .A(II31823) );
  INV_X1 NOT_9334( .ZN(II31826), .A(g23895) );
  INV_X1 NOT_9335( .ZN(g24384), .A(II31826) );
  INV_X1 NOT_9336( .ZN(II31829), .A(g23871) );
  INV_X1 NOT_9337( .ZN(g24385), .A(II31829) );
  INV_X1 NOT_9338( .ZN(II31832), .A(g23896) );
  INV_X1 NOT_9339( .ZN(g24386), .A(II31832) );
  INV_X1 NOT_9340( .ZN(II31835), .A(g23911) );
  INV_X1 NOT_9341( .ZN(g24387), .A(II31835) );
  INV_X1 NOT_9342( .ZN(II31838), .A(g23585) );
  INV_X1 NOT_9343( .ZN(g24388), .A(II31838) );
  INV_X1 NOT_9344( .ZN(II31841), .A(g23607) );
  INV_X1 NOT_9345( .ZN(g24389), .A(II31841) );
  INV_X1 NOT_9346( .ZN(II31844), .A(g23633) );
  INV_X1 NOT_9347( .ZN(g24390), .A(II31844) );
  INV_X1 NOT_9348( .ZN(II31847), .A(g23608) );
  INV_X1 NOT_9349( .ZN(g24391), .A(II31847) );
  INV_X1 NOT_9350( .ZN(II31850), .A(g23634) );
  INV_X1 NOT_9351( .ZN(g24392), .A(II31850) );
  INV_X1 NOT_9352( .ZN(II31853), .A(g23676) );
  INV_X1 NOT_9353( .ZN(g24393), .A(II31853) );
  INV_X1 NOT_9354( .ZN(II31856), .A(g23635) );
  INV_X1 NOT_9355( .ZN(g24394), .A(II31856) );
  INV_X1 NOT_9356( .ZN(II31859), .A(g23677) );
  INV_X1 NOT_9357( .ZN(g24395), .A(II31859) );
  INV_X1 NOT_9358( .ZN(II31862), .A(g23718) );
  INV_X1 NOT_9359( .ZN(g24396), .A(II31862) );
  INV_X1 NOT_9360( .ZN(II31865), .A(g23678) );
  INV_X1 NOT_9361( .ZN(g24397), .A(II31865) );
  INV_X1 NOT_9362( .ZN(II31868), .A(g23719) );
  INV_X1 NOT_9363( .ZN(g24398), .A(II31868) );
  INV_X1 NOT_9364( .ZN(II31871), .A(g23765) );
  INV_X1 NOT_9365( .ZN(g24399), .A(II31871) );
  INV_X1 NOT_9366( .ZN(II31874), .A(g23720) );
  INV_X1 NOT_9367( .ZN(g24400), .A(II31874) );
  INV_X1 NOT_9368( .ZN(II31877), .A(g23766) );
  INV_X1 NOT_9369( .ZN(g24401), .A(II31877) );
  INV_X1 NOT_9370( .ZN(II31880), .A(g23799) );
  INV_X1 NOT_9371( .ZN(g24402), .A(II31880) );
  INV_X1 NOT_9372( .ZN(II31883), .A(g23767) );
  INV_X1 NOT_9373( .ZN(g24403), .A(II31883) );
  INV_X1 NOT_9374( .ZN(II31886), .A(g23800) );
  INV_X1 NOT_9375( .ZN(g24404), .A(II31886) );
  INV_X1 NOT_9376( .ZN(II31889), .A(g23845) );
  INV_X1 NOT_9377( .ZN(g24405), .A(II31889) );
  INV_X1 NOT_9378( .ZN(II31892), .A(g23801) );
  INV_X1 NOT_9379( .ZN(g24406), .A(II31892) );
  INV_X1 NOT_9380( .ZN(II31895), .A(g23846) );
  INV_X1 NOT_9381( .ZN(g24407), .A(II31895) );
  INV_X1 NOT_9382( .ZN(II31898), .A(g23872) );
  INV_X1 NOT_9383( .ZN(g24408), .A(II31898) );
  INV_X1 NOT_9384( .ZN(II31901), .A(g23847) );
  INV_X1 NOT_9385( .ZN(g24409), .A(II31901) );
  INV_X1 NOT_9386( .ZN(II31904), .A(g23873) );
  INV_X1 NOT_9387( .ZN(g24410), .A(II31904) );
  INV_X1 NOT_9388( .ZN(II31907), .A(g23897) );
  INV_X1 NOT_9389( .ZN(g24411), .A(II31907) );
  INV_X1 NOT_9390( .ZN(II31910), .A(g23542) );
  INV_X1 NOT_9391( .ZN(g24412), .A(II31910) );
  INV_X1 NOT_9392( .ZN(II31913), .A(g23468) );
  INV_X1 NOT_9393( .ZN(g24413), .A(II31913) );
  INV_X1 NOT_9394( .ZN(II31916), .A(g23485) );
  INV_X1 NOT_9395( .ZN(g24414), .A(II31916) );
  INV_X1 NOT_9396( .ZN(II31919), .A(g23524) );
  INV_X1 NOT_9397( .ZN(g24415), .A(II31919) );
  INV_X1 NOT_9398( .ZN(II31922), .A(g23543) );
  INV_X1 NOT_9399( .ZN(g24416), .A(II31922) );
  INV_X1 NOT_9400( .ZN(II31925), .A(g23469) );
  INV_X1 NOT_9401( .ZN(g24417), .A(II31925) );
  INV_X1 NOT_9402( .ZN(II31928), .A(g24255) );
  INV_X1 NOT_9403( .ZN(g24418), .A(II31928) );
  INV_X1 NOT_9404( .ZN(II31931), .A(g23725) );
  INV_X1 NOT_9405( .ZN(g24419), .A(II31931) );
  INV_X1 NOT_9406( .ZN(II31934), .A(g24068) );
  INV_X1 NOT_9407( .ZN(g24420), .A(II31934) );
  INV_X1 NOT_9408( .ZN(II31937), .A(g24079) );
  INV_X1 NOT_9409( .ZN(g24421), .A(II31937) );
  INV_X1 NOT_9410( .ZN(II31940), .A(g24088) );
  INV_X1 NOT_9411( .ZN(g24422), .A(II31940) );
  INV_X1 NOT_9412( .ZN(II31943), .A(g24000) );
  INV_X1 NOT_9413( .ZN(g24423), .A(II31943) );
  INV_X1 NOT_9414( .ZN(II31946), .A(g23916) );
  INV_X1 NOT_9415( .ZN(g24424), .A(II31946) );
  INV_X1 NOT_9416( .ZN(II31949), .A(g23943) );
  INV_X1 NOT_9417( .ZN(g24425), .A(II31949) );
  INV_X1 NOT_9418( .ZN(g24482), .A(g24183) );
  INV_X1 NOT_9419( .ZN(II32042), .A(g23399) );
  INV_X1 NOT_9420( .ZN(g24518), .A(II32042) );
  INV_X1 NOT_9421( .ZN(II32057), .A(g23406) );
  INV_X1 NOT_9422( .ZN(g24531), .A(II32057) );
  INV_X1 NOT_9423( .ZN(II32067), .A(g24174) );
  INV_X8 NOT_9424( .ZN(g24539), .A(II32067) );
  INV_X8 NOT_9425( .ZN(II32074), .A(g23413) );
  INV_X1 NOT_9426( .ZN(g24544), .A(II32074) );
  INV_X1 NOT_9427( .ZN(II32081), .A(g24178) );
  INV_X1 NOT_9428( .ZN(g24549), .A(II32081) );
  INV_X1 NOT_9429( .ZN(II32085), .A(g24179) );
  INV_X1 NOT_9430( .ZN(g24551), .A(II32085) );
  INV_X1 NOT_9431( .ZN(II32092), .A(g23418) );
  INV_X1 NOT_9432( .ZN(g24556), .A(II32092) );
  INV_X1 NOT_9433( .ZN(II32098), .A(g24181) );
  INV_X1 NOT_9434( .ZN(g24560), .A(II32098) );
  INV_X1 NOT_9435( .ZN(II32102), .A(g24182) );
  INV_X1 NOT_9436( .ZN(g24562), .A(II32102) );
  INV_X1 NOT_9437( .ZN(II32109), .A(g24206) );
  INV_X1 NOT_9438( .ZN(g24567), .A(II32109) );
  INV_X1 NOT_9439( .ZN(II32112), .A(g24207) );
  INV_X1 NOT_9440( .ZN(g24568), .A(II32112) );
  INV_X1 NOT_9441( .ZN(II32116), .A(g24208) );
  INV_X1 NOT_9442( .ZN(g24570), .A(II32116) );
  INV_X1 NOT_9443( .ZN(II32120), .A(g24209) );
  INV_X1 NOT_9444( .ZN(g24572), .A(II32120) );
  INV_X1 NOT_9445( .ZN(II32126), .A(g24212) );
  INV_X1 NOT_9446( .ZN(g24576), .A(II32126) );
  INV_X1 NOT_9447( .ZN(II32129), .A(g24213) );
  INV_X1 NOT_9448( .ZN(g24577), .A(II32129) );
  INV_X1 NOT_9449( .ZN(II32133), .A(g24214) );
  INV_X1 NOT_9450( .ZN(g24579), .A(II32133) );
  INV_X1 NOT_9451( .ZN(II32137), .A(g24215) );
  INV_X1 NOT_9452( .ZN(g24581), .A(II32137) );
  INV_X1 NOT_9453( .ZN(II32140), .A(g24216) );
  INV_X1 NOT_9454( .ZN(g24582), .A(II32140) );
  INV_X1 NOT_9455( .ZN(II32143), .A(g24218) );
  INV_X1 NOT_9456( .ZN(g24583), .A(II32143) );
  INV_X1 NOT_9457( .ZN(II32146), .A(g24219) );
  INV_X1 NOT_9458( .ZN(g24584), .A(II32146) );
  INV_X1 NOT_9459( .ZN(II32150), .A(g24222) );
  INV_X1 NOT_9460( .ZN(g24586), .A(II32150) );
  INV_X1 NOT_9461( .ZN(II32153), .A(g24223) );
  INV_X1 NOT_9462( .ZN(g24587), .A(II32153) );
  INV_X1 NOT_9463( .ZN(II32156), .A(g24225) );
  INV_X1 NOT_9464( .ZN(g24588), .A(II32156) );
  INV_X1 NOT_9465( .ZN(II32159), .A(g24226) );
  INV_X1 NOT_9466( .ZN(g24589), .A(II32159) );
  INV_X1 NOT_9467( .ZN(II32164), .A(g24228) );
  INV_X1 NOT_9468( .ZN(g24592), .A(II32164) );
  INV_X1 NOT_9469( .ZN(II32167), .A(g24230) );
  INV_X1 NOT_9470( .ZN(g24593), .A(II32167) );
  INV_X1 NOT_9471( .ZN(II32170), .A(g24231) );
  INV_X1 NOT_9472( .ZN(g24594), .A(II32170) );
  INV_X1 NOT_9473( .ZN(II32175), .A(g24235) );
  INV_X1 NOT_9474( .ZN(g24597), .A(II32175) );
  INV_X1 NOT_9475( .ZN(II32178), .A(g24237) );
  INV_X1 NOT_9476( .ZN(g24598), .A(II32178) );
  INV_X1 NOT_9477( .ZN(II32181), .A(g24238) );
  INV_X1 NOT_9478( .ZN(g24599), .A(II32181) );
  INV_X1 NOT_9479( .ZN(II32184), .A(g23497) );
  INV_X1 NOT_9480( .ZN(g24600), .A(II32184) );
  INV_X1 NOT_9481( .ZN(II32189), .A(g24243) );
  INV_X1 NOT_9482( .ZN(g24605), .A(II32189) );
  INV_X8 NOT_9483( .ZN(II32193), .A(g23513) );
  INV_X1 NOT_9484( .ZN(g24607), .A(II32193) );
  INV_X1 NOT_9485( .ZN(II32198), .A(g24250) );
  INV_X1 NOT_9486( .ZN(g24612), .A(II32198) );
  INV_X1 NOT_9487( .ZN(II32203), .A(g23528) );
  INV_X1 NOT_9488( .ZN(g24619), .A(II32203) );
  INV_X1 NOT_9489( .ZN(II32210), .A(g23539) );
  INV_X1 NOT_9490( .ZN(g24630), .A(II32210) );
  INV_X1 NOT_9491( .ZN(g24648), .A(g23470) );
  INV_X1 NOT_9492( .ZN(g24668), .A(g23482) );
  INV_X1 NOT_9493( .ZN(g24687), .A(g23493) );
  INV_X1 NOT_9494( .ZN(g24704), .A(g23509) );
  INV_X1 NOT_9495( .ZN(II32248), .A(g23919) );
  INV_X1 NOT_9496( .ZN(g24734), .A(II32248) );
  INV_X1 NOT_9497( .ZN(II32251), .A(g23919) );
  INV_X1 NOT_9498( .ZN(g24735), .A(II32251) );
  INV_X1 NOT_9499( .ZN(II32281), .A(g23950) );
  INV_X1 NOT_9500( .ZN(g24763), .A(II32281) );
  INV_X1 NOT_9501( .ZN(II32320), .A(g23979) );
  INV_X1 NOT_9502( .ZN(g24784), .A(II32320) );
  INV_X1 NOT_9503( .ZN(II32365), .A(g24009) );
  INV_X1 NOT_9504( .ZN(g24805), .A(II32365) );
  INV_X1 NOT_9505( .ZN(g24815), .A(g23448) );
  INV_X1 NOT_9506( .ZN(II32388), .A(g23385) );
  INV_X1 NOT_9507( .ZN(g24816), .A(II32388) );
  INV_X1 NOT_9508( .ZN(II32419), .A(g24043) );
  INV_X1 NOT_9509( .ZN(g24827), .A(II32419) );
  INV_X1 NOT_9510( .ZN(g24834), .A(g23455) );
  INV_X1 NOT_9511( .ZN(II32439), .A(g23392) );
  INV_X1 NOT_9512( .ZN(g24835), .A(II32439) );
  INV_X1 NOT_9513( .ZN(g24850), .A(g23464) );
  INV_X1 NOT_9514( .ZN(II32487), .A(g23400) );
  INV_X1 NOT_9515( .ZN(g24851), .A(II32487) );
  INV_X1 NOT_9516( .ZN(II32506), .A(g23324) );
  INV_X1 NOT_9517( .ZN(g24856), .A(II32506) );
  INV_X1 NOT_9518( .ZN(g24864), .A(g23473) );
  INV_X1 NOT_9519( .ZN(II32535), .A(g23407) );
  INV_X1 NOT_9520( .ZN(g24865), .A(II32535) );
  INV_X1 NOT_9521( .ZN(II32556), .A(g23329) );
  INV_X1 NOT_9522( .ZN(g24872), .A(II32556) );
  INV_X1 NOT_9523( .ZN(II32583), .A(g23330) );
  INV_X1 NOT_9524( .ZN(g24879), .A(II32583) );
  INV_X1 NOT_9525( .ZN(II32604), .A(g23339) );
  INV_X1 NOT_9526( .ZN(g24886), .A(II32604) );
  INV_X1 NOT_9527( .ZN(g24893), .A(g23486) );
  INV_X1 NOT_9528( .ZN(II32642), .A(g23348) );
  INV_X1 NOT_9529( .ZN(g24903), .A(II32642) );
  INV_X1 NOT_9530( .ZN(g24912), .A(g23495) );
  INV_X1 NOT_9531( .ZN(g24916), .A(g23502) );
  INV_X1 NOT_9532( .ZN(g24929), .A(g23511) );
  INV_X1 NOT_9533( .ZN(g24933), .A(g23518) );
  INV_X1 NOT_9534( .ZN(g24939), .A(g23660) );
  INV_X1 NOT_9535( .ZN(g24941), .A(g23526) );
  INV_X1 NOT_9536( .ZN(g24945), .A(g23533) );
  INV_X1 NOT_9537( .ZN(II32704), .A(g23357) );
  INV_X1 NOT_9538( .ZN(g24949), .A(II32704) );
  INV_X1 NOT_9539( .ZN(g24950), .A(g23710) );
  INV_X1 NOT_9540( .ZN(g24952), .A(g23537) );
  INV_X1 NOT_9541( .ZN(II32716), .A(g23358) );
  INV_X1 NOT_9542( .ZN(g24956), .A(II32716) );
  INV_X1 NOT_9543( .ZN(II32719), .A(g23359) );
  INV_X1 NOT_9544( .ZN(g24957), .A(II32719) );
  INV_X1 NOT_9545( .ZN(g24958), .A(g23478) );
  INV_X1 NOT_9546( .ZN(g24962), .A(g23764) );
  INV_X1 NOT_9547( .ZN(g24969), .A(g23489) );
  INV_X1 NOT_9548( .ZN(g24973), .A(g23819) );
  INV_X1 NOT_9549( .ZN(g24982), .A(g23505) );
  INV_X1 NOT_9550( .ZN(g24993), .A(g23521) );
  INV_X1 NOT_9551( .ZN(g25087), .A(g23731) );
  INV_X1 NOT_9552( .ZN(g25094), .A(g23779) );
  INV_X1 NOT_9553( .ZN(g25095), .A(g23786) );
  INV_X1 NOT_9554( .ZN(II32829), .A(g24059) );
  INV_X1 NOT_9555( .ZN(g25103), .A(II32829) );
  INV_X1 NOT_9556( .ZN(g25104), .A(g23832) );
  INV_X1 NOT_9557( .ZN(g25105), .A(g23839) );
  INV_X1 NOT_9558( .ZN(II32835), .A(g24072) );
  INV_X1 NOT_9559( .ZN(g25109), .A(II32835) );
  INV_X1 NOT_9560( .ZN(g25110), .A(g23867) );
  INV_X1 NOT_9561( .ZN(g25111), .A(g23874) );
  INV_X1 NOT_9562( .ZN(g25115), .A(g23879) );
  INV_X1 NOT_9563( .ZN(g25116), .A(g23882) );
  INV_X1 NOT_9564( .ZN(II32844), .A(g23644) );
  INV_X1 NOT_9565( .ZN(g25118), .A(II32844) );
  INV_X1 NOT_9566( .ZN(II32847), .A(g24083) );
  INV_X1 NOT_9567( .ZN(g25119), .A(II32847) );
  INV_X1 NOT_9568( .ZN(g25120), .A(g23901) );
  INV_X1 NOT_9569( .ZN(II32851), .A(g23694) );
  INV_X1 NOT_9570( .ZN(g25121), .A(II32851) );
  INV_X1 NOT_9571( .ZN(II32854), .A(g24092) );
  INV_X1 NOT_9572( .ZN(g25122), .A(II32854) );
  INV_X1 NOT_9573( .ZN(II32857), .A(g23748) );
  INV_X1 NOT_9574( .ZN(g25123), .A(II32857) );
  INV_X1 NOT_9575( .ZN(II32860), .A(g23803) );
  INV_X1 NOT_9576( .ZN(g25124), .A(II32860) );
  INV_X1 NOT_9577( .ZN(g25126), .A(g24030) );
  INV_X1 NOT_9578( .ZN(II32868), .A(g25118) );
  INV_X1 NOT_9579( .ZN(g25130), .A(II32868) );
  INV_X1 NOT_9580( .ZN(II32871), .A(g24518) );
  INV_X1 NOT_9581( .ZN(g25131), .A(II32871) );
  INV_X1 NOT_9582( .ZN(II32874), .A(g24539) );
  INV_X1 NOT_9583( .ZN(g25132), .A(II32874) );
  INV_X1 NOT_9584( .ZN(II32877), .A(g24567) );
  INV_X1 NOT_9585( .ZN(g25133), .A(II32877) );
  INV_X1 NOT_9586( .ZN(II32880), .A(g24581) );
  INV_X1 NOT_9587( .ZN(g25134), .A(II32880) );
  INV_X1 NOT_9588( .ZN(II32883), .A(g24592) );
  INV_X1 NOT_9589( .ZN(g25135), .A(II32883) );
  INV_X1 NOT_9590( .ZN(II32886), .A(g24549) );
  INV_X1 NOT_9591( .ZN(g25136), .A(II32886) );
  INV_X1 NOT_9592( .ZN(II32889), .A(g24568) );
  INV_X1 NOT_9593( .ZN(g25137), .A(II32889) );
  INV_X1 NOT_9594( .ZN(II32892), .A(g24582) );
  INV_X1 NOT_9595( .ZN(g25138), .A(II32892) );
  INV_X1 NOT_9596( .ZN(II32895), .A(g24816) );
  INV_X1 NOT_9597( .ZN(g25139), .A(II32895) );
  INV_X1 NOT_9598( .ZN(II32898), .A(g24856) );
  INV_X1 NOT_9599( .ZN(g25140), .A(II32898) );
  INV_X1 NOT_9600( .ZN(II32901), .A(g25121) );
  INV_X8 NOT_9601( .ZN(g25141), .A(II32901) );
  INV_X8 NOT_9602( .ZN(II32904), .A(g24531) );
  INV_X1 NOT_9603( .ZN(g25142), .A(II32904) );
  INV_X1 NOT_9604( .ZN(II32907), .A(g24551) );
  INV_X1 NOT_9605( .ZN(g25143), .A(II32907) );
  INV_X1 NOT_9606( .ZN(II32910), .A(g24576) );
  INV_X1 NOT_9607( .ZN(g25144), .A(II32910) );
  INV_X1 NOT_9608( .ZN(II32913), .A(g24586) );
  INV_X1 NOT_9609( .ZN(g25145), .A(II32913) );
  INV_X1 NOT_9610( .ZN(II32916), .A(g24597) );
  INV_X1 NOT_9611( .ZN(g25146), .A(II32916) );
  INV_X1 NOT_9612( .ZN(II32919), .A(g24560) );
  INV_X1 NOT_9613( .ZN(g25147), .A(II32919) );
  INV_X1 NOT_9614( .ZN(II32922), .A(g24577) );
  INV_X1 NOT_9615( .ZN(g25148), .A(II32922) );
  INV_X1 NOT_9616( .ZN(II32925), .A(g24587) );
  INV_X1 NOT_9617( .ZN(g25149), .A(II32925) );
  INV_X1 NOT_9618( .ZN(II32928), .A(g24835) );
  INV_X1 NOT_9619( .ZN(g25150), .A(II32928) );
  INV_X1 NOT_9620( .ZN(II32931), .A(g24872) );
  INV_X1 NOT_9621( .ZN(g25151), .A(II32931) );
  INV_X1 NOT_9622( .ZN(II32934), .A(g25123) );
  INV_X1 NOT_9623( .ZN(g25152), .A(II32934) );
  INV_X1 NOT_9624( .ZN(II32937), .A(g24544) );
  INV_X1 NOT_9625( .ZN(g25153), .A(II32937) );
  INV_X1 NOT_9626( .ZN(II32940), .A(g24562) );
  INV_X1 NOT_9627( .ZN(g25154), .A(II32940) );
  INV_X1 NOT_9628( .ZN(II32943), .A(g24583) );
  INV_X1 NOT_9629( .ZN(g25155), .A(II32943) );
  INV_X1 NOT_9630( .ZN(II32946), .A(g24593) );
  INV_X1 NOT_9631( .ZN(g25156), .A(II32946) );
  INV_X1 NOT_9632( .ZN(II32949), .A(g24605) );
  INV_X1 NOT_9633( .ZN(g25157), .A(II32949) );
  INV_X1 NOT_9634( .ZN(II32952), .A(g24570) );
  INV_X1 NOT_9635( .ZN(g25158), .A(II32952) );
  INV_X1 NOT_9636( .ZN(II32955), .A(g24584) );
  INV_X1 NOT_9637( .ZN(g25159), .A(II32955) );
  INV_X1 NOT_9638( .ZN(II32958), .A(g24594) );
  INV_X1 NOT_9639( .ZN(g25160), .A(II32958) );
  INV_X1 NOT_9640( .ZN(II32961), .A(g24851) );
  INV_X1 NOT_9641( .ZN(g25161), .A(II32961) );
  INV_X1 NOT_9642( .ZN(II32964), .A(g24886) );
  INV_X1 NOT_9643( .ZN(g25162), .A(II32964) );
  INV_X1 NOT_9644( .ZN(II32967), .A(g25124) );
  INV_X1 NOT_9645( .ZN(g25163), .A(II32967) );
  INV_X1 NOT_9646( .ZN(II32970), .A(g24556) );
  INV_X1 NOT_9647( .ZN(g25164), .A(II32970) );
  INV_X1 NOT_9648( .ZN(II32973), .A(g24572) );
  INV_X1 NOT_9649( .ZN(g25165), .A(II32973) );
  INV_X1 NOT_9650( .ZN(II32976), .A(g24588) );
  INV_X1 NOT_9651( .ZN(g25166), .A(II32976) );
  INV_X1 NOT_9652( .ZN(II32979), .A(g24598) );
  INV_X1 NOT_9653( .ZN(g25167), .A(II32979) );
  INV_X1 NOT_9654( .ZN(II32982), .A(g24612) );
  INV_X1 NOT_9655( .ZN(g25168), .A(II32982) );
  INV_X1 NOT_9656( .ZN(II32985), .A(g24579) );
  INV_X1 NOT_9657( .ZN(g25169), .A(II32985) );
  INV_X1 NOT_9658( .ZN(II32988), .A(g24589) );
  INV_X1 NOT_9659( .ZN(g25170), .A(II32988) );
  INV_X1 NOT_9660( .ZN(II32991), .A(g24599) );
  INV_X1 NOT_9661( .ZN(g25171), .A(II32991) );
  INV_X1 NOT_9662( .ZN(II32994), .A(g24865) );
  INV_X1 NOT_9663( .ZN(g25172), .A(II32994) );
  INV_X1 NOT_9664( .ZN(II32997), .A(g24903) );
  INV_X1 NOT_9665( .ZN(g25173), .A(II32997) );
  INV_X1 NOT_9666( .ZN(II33000), .A(g24949) );
  INV_X1 NOT_9667( .ZN(g25174), .A(II33000) );
  INV_X1 NOT_9668( .ZN(II33003), .A(g24956) );
  INV_X1 NOT_9669( .ZN(g25175), .A(II33003) );
  INV_X1 NOT_9670( .ZN(II33006), .A(g24957) );
  INV_X1 NOT_9671( .ZN(g25176), .A(II33006) );
  INV_X1 NOT_9672( .ZN(II33009), .A(g24879) );
  INV_X1 NOT_9673( .ZN(g25177), .A(II33009) );
  INV_X1 NOT_9674( .ZN(II33013), .A(g25119) );
  INV_X1 NOT_9675( .ZN(g25179), .A(II33013) );
  INV_X1 NOT_9676( .ZN(II33016), .A(g25122) );
  INV_X1 NOT_9677( .ZN(g25180), .A(II33016) );
  INV_X1 NOT_9678( .ZN(g25274), .A(g24912) );
  INV_X1 NOT_9679( .ZN(g25283), .A(g24929) );
  INV_X1 NOT_9680( .ZN(g25291), .A(g24941) );
  INV_X1 NOT_9681( .ZN(II33128), .A(g24975) );
  INV_X1 NOT_9682( .ZN(g25296), .A(II33128) );
  INV_X1 NOT_9683( .ZN(g25301), .A(g24952) );
  INV_X1 NOT_9684( .ZN(g25305), .A(g24880) );
  INV_X1 NOT_9685( .ZN(II33136), .A(g24986) );
  INV_X1 NOT_9686( .ZN(g25306), .A(II33136) );
  INV_X1 NOT_9687( .ZN(g25313), .A(g24868) );
  INV_X1 NOT_9688( .ZN(g25314), .A(g24897) );
  INV_X1 NOT_9689( .ZN(II33145), .A(g24997) );
  INV_X1 NOT_9690( .ZN(g25315), .A(II33145) );
  INV_X1 NOT_9691( .ZN(g25319), .A(g24857) );
  INV_X1 NOT_9692( .ZN(g25322), .A(g24883) );
  INV_X1 NOT_9693( .ZN(g25323), .A(g24920) );
  INV_X1 NOT_9694( .ZN(II33154), .A(g25005) );
  INV_X1 NOT_9695( .ZN(g25324), .A(II33154) );
  INV_X1 NOT_9696( .ZN(II33157), .A(g25027) );
  INV_X1 NOT_9697( .ZN(g25327), .A(II33157) );
  INV_X1 NOT_9698( .ZN(g25329), .A(g24844) );
  INV_X1 NOT_9699( .ZN(g25330), .A(g24873) );
  INV_X1 NOT_9700( .ZN(g25332), .A(g24900) );
  INV_X1 NOT_9701( .ZN(g25333), .A(g24937) );
  INV_X1 NOT_9702( .ZN(g25335), .A(g24832) );
  INV_X1 NOT_9703( .ZN(II33168), .A(g25042) );
  INV_X1 NOT_9704( .ZN(g25336), .A(II33168) );
  INV_X1 NOT_9705( .ZN(g25338), .A(g24860) );
  INV_X1 NOT_9706( .ZN(g25339), .A(g24887) );
  INV_X1 NOT_9707( .ZN(g25341), .A(g24923) );
  INV_X1 NOT_9708( .ZN(g25347), .A(g24817) );
  INV_X1 NOT_9709( .ZN(g25349), .A(g24848) );
  INV_X1 NOT_9710( .ZN(II33182), .A(g25056) );
  INV_X1 NOT_9711( .ZN(g25350), .A(II33182) );
  INV_X1 NOT_9712( .ZN(g25352), .A(g24875) );
  INV_X1 NOT_9713( .ZN(g25353), .A(g24904) );
  INV_X1 NOT_9714( .ZN(II33188), .A(g24814) );
  INV_X1 NOT_9715( .ZN(g25354), .A(II33188) );
  INV_X1 NOT_9716( .ZN(g25355), .A(g24797) );
  INV_X1 NOT_9717( .ZN(g25361), .A(g24837) );
  INV_X1 NOT_9718( .ZN(g25363), .A(g24862) );
  INV_X1 NOT_9719( .ZN(II33198), .A(g25067) );
  INV_X1 NOT_9720( .ZN(g25364), .A(II33198) );
  INV_X1 NOT_9721( .ZN(g25366), .A(g24889) );
  INV_X1 NOT_9722( .ZN(g25367), .A(g24676) );
  INV_X1 NOT_9723( .ZN(g25368), .A(g24778) );
  INV_X1 NOT_9724( .ZN(II33205), .A(g24833) );
  INV_X1 NOT_9725( .ZN(g25369), .A(II33205) );
  INV_X1 NOT_9726( .ZN(g25370), .A(g24820) );
  INV_X1 NOT_9727( .ZN(g25376), .A(g24852) );
  INV_X1 NOT_9728( .ZN(g25378), .A(g24877) );
  INV_X1 NOT_9729( .ZN(g25379), .A(g24893) );
  INV_X1 NOT_9730( .ZN(g25383), .A(g24766) );
  INV_X1 NOT_9731( .ZN(g25384), .A(g24695) );
  INV_X1 NOT_9732( .ZN(g25385), .A(g24801) );
  INV_X1 NOT_9733( .ZN(II33219), .A(g24849) );
  INV_X1 NOT_9734( .ZN(g25386), .A(II33219) );
  INV_X1 NOT_9735( .ZN(g25387), .A(g24839) );
  INV_X1 NOT_9736( .ZN(g25393), .A(g24866) );
  INV_X1 NOT_9737( .ZN(g25394), .A(g24753) );
  INV_X1 NOT_9738( .ZN(g25395), .A(g24916) );
  INV_X1 NOT_9739( .ZN(g25399), .A(g24787) );
  INV_X1 NOT_9740( .ZN(g25400), .A(g24712) );
  INV_X1 NOT_9741( .ZN(g25401), .A(g24823) );
  INV_X1 NOT_9742( .ZN(II33232), .A(g24863) );
  INV_X1 NOT_9743( .ZN(g25402), .A(II33232) );
  INV_X1 NOT_9744( .ZN(g25403), .A(g24854) );
  INV_X1 NOT_9745( .ZN(g25404), .A(g24771) );
  INV_X1 NOT_9746( .ZN(g25405), .A(g24933) );
  INV_X1 NOT_9747( .ZN(g25409), .A(g24808) );
  INV_X1 NOT_9748( .ZN(g25410), .A(g24723) );
  INV_X1 NOT_9749( .ZN(g25411), .A(g24842) );
  INV_X1 NOT_9750( .ZN(g25412), .A(g24791) );
  INV_X1 NOT_9751( .ZN(g25413), .A(g24945) );
  INV_X1 NOT_9752( .ZN(g25417), .A(g24830) );
  INV_X1 NOT_9753( .ZN(g25419), .A(g24812) );
  INV_X1 NOT_9754( .ZN(II33246), .A(g24890) );
  INV_X1 NOT_9755( .ZN(g25420), .A(II33246) );
  INV_X1 NOT_9756( .ZN(II33249), .A(g24890) );
  INV_X1 NOT_9757( .ZN(g25421), .A(II33249) );
  INV_X1 NOT_9758( .ZN(g25422), .A(g24958) );
  INV_X1 NOT_9759( .ZN(g25430), .A(g24616) );
  INV_X1 NOT_9760( .ZN(g25431), .A(g24969) );
  INV_X1 NOT_9761( .ZN(II33257), .A(g24909) );
  INV_X1 NOT_9762( .ZN(g25435), .A(II33257) );
  INV_X1 NOT_9763( .ZN(II33260), .A(g24909) );
  INV_X1 NOT_9764( .ZN(g25436), .A(II33260) );
  INV_X1 NOT_9765( .ZN(g25437), .A(g24627) );
  INV_X1 NOT_9766( .ZN(g25438), .A(g24982) );
  INV_X1 NOT_9767( .ZN(II33265), .A(g24925) );
  INV_X1 NOT_9768( .ZN(g25442), .A(II33265) );
  INV_X1 NOT_9769( .ZN(II33268), .A(g24925) );
  INV_X1 NOT_9770( .ZN(g25443), .A(II33268) );
  INV_X1 NOT_9771( .ZN(g25444), .A(g24641) );
  INV_X4 NOT_9772( .ZN(g25445), .A(g24993) );
  INV_X4 NOT_9773( .ZN(g25449), .A(g24660) );
  INV_X4 NOT_9774( .ZN(II33278), .A(g25088) );
  INV_X1 NOT_9775( .ZN(g25454), .A(II33278) );
  INV_X1 NOT_9776( .ZN(II33282), .A(g25096) );
  INV_X1 NOT_9777( .ZN(g25458), .A(II33282) );
  INV_X1 NOT_9778( .ZN(II33286), .A(g24426) );
  INV_X1 NOT_9779( .ZN(g25462), .A(II33286) );
  INV_X1 NOT_9780( .ZN(II33289), .A(g25106) );
  INV_X1 NOT_9781( .ZN(g25463), .A(II33289) );
  INV_X1 NOT_9782( .ZN(II33293), .A(g25008) );
  INV_X1 NOT_9783( .ZN(g25467), .A(II33293) );
  INV_X1 NOT_9784( .ZN(II33297), .A(g24430) );
  INV_X1 NOT_9785( .ZN(g25471), .A(II33297) );
  INV_X1 NOT_9786( .ZN(II33300), .A(g25112) );
  INV_X1 NOT_9787( .ZN(g25472), .A(II33300) );
  INV_X1 NOT_9788( .ZN(II33304), .A(g25004) );
  INV_X1 NOT_9789( .ZN(g25476), .A(II33304) );
  INV_X1 NOT_9790( .ZN(II33307), .A(g25011) );
  INV_X1 NOT_9791( .ZN(g25479), .A(II33307) );
  INV_X1 NOT_9792( .ZN(II33312), .A(g25014) );
  INV_X1 NOT_9793( .ZN(g25484), .A(II33312) );
  INV_X1 NOT_9794( .ZN(II33316), .A(g24434) );
  INV_X1 NOT_9795( .ZN(g25488), .A(II33316) );
  INV_X1 NOT_9796( .ZN(II33321), .A(g24442) );
  INV_X1 NOT_9797( .ZN(g25493), .A(II33321) );
  INV_X1 NOT_9798( .ZN(II33324), .A(g25009) );
  INV_X1 NOT_9799( .ZN(g25496), .A(II33324) );
  INV_X1 NOT_9800( .ZN(II33327), .A(g25017) );
  INV_X1 NOT_9801( .ZN(g25499), .A(II33327) );
  INV_X1 NOT_9802( .ZN(II33330), .A(g25019) );
  INV_X1 NOT_9803( .ZN(g25502), .A(II33330) );
  INV_X1 NOT_9804( .ZN(II33335), .A(g25010) );
  INV_X1 NOT_9805( .ZN(g25507), .A(II33335) );
  INV_X1 NOT_9806( .ZN(II33338), .A(g25021) );
  INV_X1 NOT_9807( .ZN(g25510), .A(II33338) );
  INV_X1 NOT_9808( .ZN(II33343), .A(g25024) );
  INV_X1 NOT_9809( .ZN(g25515), .A(II33343) );
  INV_X1 NOT_9810( .ZN(II33347), .A(g24438) );
  INV_X1 NOT_9811( .ZN(g25519), .A(II33347) );
  INV_X1 NOT_9812( .ZN(II33352), .A(g24443) );
  INV_X1 NOT_9813( .ZN(g25524), .A(II33352) );
  INV_X1 NOT_9814( .ZN(II33355), .A(g25012) );
  INV_X1 NOT_9815( .ZN(g25527), .A(II33355) );
  INV_X1 NOT_9816( .ZN(II33358), .A(g25028) );
  INV_X1 NOT_9817( .ZN(g25530), .A(II33358) );
  INV_X1 NOT_9818( .ZN(II33361), .A(g25013) );
  INV_X1 NOT_9819( .ZN(g25533), .A(II33361) );
  INV_X1 NOT_9820( .ZN(II33364), .A(g25029) );
  INV_X1 NOT_9821( .ZN(g25536), .A(II33364) );
  INV_X1 NOT_9822( .ZN(II33368), .A(g24444) );
  INV_X1 NOT_9823( .ZN(g25540), .A(II33368) );
  INV_X1 NOT_9824( .ZN(II33371), .A(g25015) );
  INV_X1 NOT_9825( .ZN(g25543), .A(II33371) );
  INV_X1 NOT_9826( .ZN(II33374), .A(g25031) );
  INV_X1 NOT_9827( .ZN(g25546), .A(II33374) );
  INV_X1 NOT_9828( .ZN(II33377), .A(g25033) );
  INV_X1 NOT_9829( .ZN(g25549), .A(II33377) );
  INV_X1 NOT_9830( .ZN(II33382), .A(g25016) );
  INV_X1 NOT_9831( .ZN(g25554), .A(II33382) );
  INV_X1 NOT_9832( .ZN(II33385), .A(g25035) );
  INV_X1 NOT_9833( .ZN(g25557), .A(II33385) );
  INV_X1 NOT_9834( .ZN(II33390), .A(g25038) );
  INV_X1 NOT_9835( .ZN(g25562), .A(II33390) );
  INV_X1 NOT_9836( .ZN(II33396), .A(g24447) );
  INV_X1 NOT_9837( .ZN(g25573), .A(II33396) );
  INV_X1 NOT_9838( .ZN(II33399), .A(g25018) );
  INV_X1 NOT_9839( .ZN(g25576), .A(II33399) );
  INV_X1 NOT_9840( .ZN(II33402), .A(g24448) );
  INV_X1 NOT_9841( .ZN(g25579), .A(II33402) );
  INV_X1 NOT_9842( .ZN(II33405), .A(g25020) );
  INV_X1 NOT_9843( .ZN(g25582), .A(II33405) );
  INV_X1 NOT_9844( .ZN(II33408), .A(g25040) );
  INV_X1 NOT_9845( .ZN(g25585), .A(II33408) );
  INV_X1 NOT_9846( .ZN(II33411), .A(g24491) );
  INV_X1 NOT_9847( .ZN(g25588), .A(II33411) );
  INV_X1 NOT_9848( .ZN(II33415), .A(g24449) );
  INV_X1 NOT_9849( .ZN(g25590), .A(II33415) );
  INV_X1 NOT_9850( .ZN(II33418), .A(g25022) );
  INV_X1 NOT_9851( .ZN(g25593), .A(II33418) );
  INV_X1 NOT_9852( .ZN(II33421), .A(g25043) );
  INV_X1 NOT_9853( .ZN(g25596), .A(II33421) );
  INV_X1 NOT_9854( .ZN(II33424), .A(g25023) );
  INV_X1 NOT_9855( .ZN(g25599), .A(II33424) );
  INV_X1 NOT_9856( .ZN(II33427), .A(g25044) );
  INV_X1 NOT_9857( .ZN(g25602), .A(II33427) );
  INV_X1 NOT_9858( .ZN(II33431), .A(g24450) );
  INV_X1 NOT_9859( .ZN(g25606), .A(II33431) );
  INV_X1 NOT_9860( .ZN(II33434), .A(g25025) );
  INV_X1 NOT_9861( .ZN(g25609), .A(II33434) );
  INV_X1 NOT_9862( .ZN(II33437), .A(g25046) );
  INV_X1 NOT_9863( .ZN(g25612), .A(II33437) );
  INV_X1 NOT_9864( .ZN(II33440), .A(g25048) );
  INV_X1 NOT_9865( .ZN(g25615), .A(II33440) );
  INV_X1 NOT_9866( .ZN(II33445), .A(g25026) );
  INV_X1 NOT_9867( .ZN(g25620), .A(II33445) );
  INV_X1 NOT_9868( .ZN(II33448), .A(g25050) );
  INV_X1 NOT_9869( .ZN(g25623), .A(II33448) );
  INV_X1 NOT_9870( .ZN(g25630), .A(g24478) );
  INV_X1 NOT_9871( .ZN(II33457), .A(g24451) );
  INV_X1 NOT_9872( .ZN(g25634), .A(II33457) );
  INV_X1 NOT_9873( .ZN(II33460), .A(g24452) );
  INV_X1 NOT_9874( .ZN(g25637), .A(II33460) );
  INV_X1 NOT_9875( .ZN(II33463), .A(g25030) );
  INV_X1 NOT_9876( .ZN(g25640), .A(II33463) );
  INV_X1 NOT_9877( .ZN(II33466), .A(g25053) );
  INV_X1 NOT_9878( .ZN(g25643), .A(II33466) );
  INV_X1 NOT_9879( .ZN(II33469), .A(g24498) );
  INV_X1 NOT_9880( .ZN(g25646), .A(II33469) );
  INV_X1 NOT_9881( .ZN(II33472), .A(g24499) );
  INV_X1 NOT_9882( .ZN(g25647), .A(II33472) );
  INV_X1 NOT_9883( .ZN(II33476), .A(g24453) );
  INV_X1 NOT_9884( .ZN(g25652), .A(II33476) );
  INV_X1 NOT_9885( .ZN(II33479), .A(g25032) );
  INV_X1 NOT_9886( .ZN(g25655), .A(II33479) );
  INV_X1 NOT_9887( .ZN(II33482), .A(g24454) );
  INV_X4 NOT_9888( .ZN(g25658), .A(II33482) );
  INV_X1 NOT_9889( .ZN(II33485), .A(g25034) );
  INV_X1 NOT_9890( .ZN(g25661), .A(II33485) );
  INV_X1 NOT_9891( .ZN(II33488), .A(g25054) );
  INV_X1 NOT_9892( .ZN(g25664), .A(II33488) );
  INV_X1 NOT_9893( .ZN(II33491), .A(g24501) );
  INV_X1 NOT_9894( .ZN(g25667), .A(II33491) );
  INV_X1 NOT_9895( .ZN(II33495), .A(g24455) );
  INV_X1 NOT_9896( .ZN(g25669), .A(II33495) );
  INV_X1 NOT_9897( .ZN(II33498), .A(g25036) );
  INV_X1 NOT_9898( .ZN(g25672), .A(II33498) );
  INV_X1 NOT_9899( .ZN(II33501), .A(g25057) );
  INV_X1 NOT_9900( .ZN(g25675), .A(II33501) );
  INV_X1 NOT_9901( .ZN(II33504), .A(g25037) );
  INV_X1 NOT_9902( .ZN(g25678), .A(II33504) );
  INV_X1 NOT_9903( .ZN(II33507), .A(g25058) );
  INV_X1 NOT_9904( .ZN(g25681), .A(II33507) );
  INV_X1 NOT_9905( .ZN(II33511), .A(g24456) );
  INV_X1 NOT_9906( .ZN(g25685), .A(II33511) );
  INV_X1 NOT_9907( .ZN(II33514), .A(g25039) );
  INV_X1 NOT_9908( .ZN(g25688), .A(II33514) );
  INV_X1 NOT_9909( .ZN(II33517), .A(g25060) );
  INV_X1 NOT_9910( .ZN(g25691), .A(II33517) );
  INV_X1 NOT_9911( .ZN(II33520), .A(g25062) );
  INV_X1 NOT_9912( .ZN(g25694), .A(II33520) );
  INV_X1 NOT_9913( .ZN(g25698), .A(g24600) );
  INV_X1 NOT_9914( .ZN(II33526), .A(g24457) );
  INV_X1 NOT_9915( .ZN(g25700), .A(II33526) );
  INV_X1 NOT_9916( .ZN(II33529), .A(g25041) );
  INV_X1 NOT_9917( .ZN(g25703), .A(II33529) );
  INV_X1 NOT_9918( .ZN(II33532), .A(g24507) );
  INV_X1 NOT_9919( .ZN(g25706), .A(II33532) );
  INV_X1 NOT_9920( .ZN(II33535), .A(g24508) );
  INV_X1 NOT_9921( .ZN(g25707), .A(II33535) );
  INV_X1 NOT_9922( .ZN(II33539), .A(g24458) );
  INV_X1 NOT_9923( .ZN(g25711), .A(II33539) );
  INV_X1 NOT_9924( .ZN(II33542), .A(g24459) );
  INV_X1 NOT_9925( .ZN(g25714), .A(II33542) );
  INV_X1 NOT_9926( .ZN(II33545), .A(g25045) );
  INV_X1 NOT_9927( .ZN(g25717), .A(II33545) );
  INV_X1 NOT_9928( .ZN(II33548), .A(g25064) );
  INV_X1 NOT_9929( .ZN(g25720), .A(II33548) );
  INV_X1 NOT_9930( .ZN(II33551), .A(g24510) );
  INV_X1 NOT_9931( .ZN(g25723), .A(II33551) );
  INV_X1 NOT_9932( .ZN(II33554), .A(g24511) );
  INV_X1 NOT_9933( .ZN(g25724), .A(II33554) );
  INV_X1 NOT_9934( .ZN(II33558), .A(g24460) );
  INV_X1 NOT_9935( .ZN(g25729), .A(II33558) );
  INV_X1 NOT_9936( .ZN(II33561), .A(g25047) );
  INV_X1 NOT_9937( .ZN(g25732), .A(II33561) );
  INV_X1 NOT_9938( .ZN(II33564), .A(g24461) );
  INV_X1 NOT_9939( .ZN(g25735), .A(II33564) );
  INV_X1 NOT_9940( .ZN(II33567), .A(g25049) );
  INV_X1 NOT_9941( .ZN(g25738), .A(II33567) );
  INV_X1 NOT_9942( .ZN(II33570), .A(g25065) );
  INV_X1 NOT_9943( .ZN(g25741), .A(II33570) );
  INV_X1 NOT_9944( .ZN(II33573), .A(g24513) );
  INV_X1 NOT_9945( .ZN(g25744), .A(II33573) );
  INV_X1 NOT_9946( .ZN(II33577), .A(g24462) );
  INV_X1 NOT_9947( .ZN(g25746), .A(II33577) );
  INV_X1 NOT_9948( .ZN(II33580), .A(g25051) );
  INV_X1 NOT_9949( .ZN(g25749), .A(II33580) );
  INV_X1 NOT_9950( .ZN(II33583), .A(g25068) );
  INV_X1 NOT_9951( .ZN(g25752), .A(II33583) );
  INV_X1 NOT_9952( .ZN(II33586), .A(g25052) );
  INV_X1 NOT_9953( .ZN(g25755), .A(II33586) );
  INV_X1 NOT_9954( .ZN(II33589), .A(g25069) );
  INV_X1 NOT_9955( .ZN(g25758), .A(II33589) );
  INV_X1 NOT_9956( .ZN(II33593), .A(g24445) );
  INV_X1 NOT_9957( .ZN(g25762), .A(II33593) );
  INV_X1 NOT_9958( .ZN(II33596), .A(g24446) );
  INV_X1 NOT_9959( .ZN(g25763), .A(II33596) );
  INV_X1 NOT_9960( .ZN(II33600), .A(g24463) );
  INV_X1 NOT_9961( .ZN(g25767), .A(II33600) );
  INV_X1 NOT_9962( .ZN(II33603), .A(g24519) );
  INV_X1 NOT_9963( .ZN(g25770), .A(II33603) );
  INV_X1 NOT_9964( .ZN(g25771), .A(g24607) );
  INV_X1 NOT_9965( .ZN(II33608), .A(g24464) );
  INV_X1 NOT_9966( .ZN(g25773), .A(II33608) );
  INV_X1 NOT_9967( .ZN(II33611), .A(g25055) );
  INV_X1 NOT_9968( .ZN(g25776), .A(II33611) );
  INV_X1 NOT_9969( .ZN(II33614), .A(g24521) );
  INV_X1 NOT_9970( .ZN(g25779), .A(II33614) );
  INV_X1 NOT_9971( .ZN(II33617), .A(g24522) );
  INV_X1 NOT_9972( .ZN(g25780), .A(II33617) );
  INV_X1 NOT_9973( .ZN(II33621), .A(g24465) );
  INV_X1 NOT_9974( .ZN(g25784), .A(II33621) );
  INV_X1 NOT_9975( .ZN(II33624), .A(g24466) );
  INV_X1 NOT_9976( .ZN(g25787), .A(II33624) );
  INV_X1 NOT_9977( .ZN(II33627), .A(g25059) );
  INV_X1 NOT_9978( .ZN(g25790), .A(II33627) );
  INV_X1 NOT_9979( .ZN(II33630), .A(g25071) );
  INV_X1 NOT_9980( .ZN(g25793), .A(II33630) );
  INV_X1 NOT_9981( .ZN(II33633), .A(g24524) );
  INV_X1 NOT_9982( .ZN(g25796), .A(II33633) );
  INV_X1 NOT_9983( .ZN(II33636), .A(g24525) );
  INV_X1 NOT_9984( .ZN(g25797), .A(II33636) );
  INV_X1 NOT_9985( .ZN(II33640), .A(g24467) );
  INV_X1 NOT_9986( .ZN(g25802), .A(II33640) );
  INV_X1 NOT_9987( .ZN(II33643), .A(g25061) );
  INV_X1 NOT_9988( .ZN(g25805), .A(II33643) );
  INV_X1 NOT_9989( .ZN(II33646), .A(g24468) );
  INV_X1 NOT_9990( .ZN(g25808), .A(II33646) );
  INV_X1 NOT_9991( .ZN(II33649), .A(g25063) );
  INV_X1 NOT_9992( .ZN(g25811), .A(II33649) );
  INV_X1 NOT_9993( .ZN(II33652), .A(g25072) );
  INV_X1 NOT_9994( .ZN(g25814), .A(II33652) );
  INV_X1 NOT_9995( .ZN(II33655), .A(g24527) );
  INV_X1 NOT_9996( .ZN(g25817), .A(II33655) );
  INV_X1 NOT_9997( .ZN(II33659), .A(g24469) );
  INV_X1 NOT_9998( .ZN(g25821), .A(II33659) );
  INV_X1 NOT_9999( .ZN(II33662), .A(g24532) );
  INV_X1 NOT_10000( .ZN(g25824), .A(II33662) );
  INV_X1 NOT_10001( .ZN(g25825), .A(g24619) );
  INV_X1 NOT_10002( .ZN(II33667), .A(g24470) );
  INV_X4 NOT_10003( .ZN(g25827), .A(II33667) );
  INV_X4 NOT_10004( .ZN(II33670), .A(g25066) );
  INV_X1 NOT_10005( .ZN(g25830), .A(II33670) );
  INV_X1 NOT_10006( .ZN(II33673), .A(g24534) );
  INV_X1 NOT_10007( .ZN(g25833), .A(II33673) );
  INV_X1 NOT_10008( .ZN(II33676), .A(g24535) );
  INV_X1 NOT_10009( .ZN(g25834), .A(II33676) );
  INV_X1 NOT_10010( .ZN(II33680), .A(g24471) );
  INV_X1 NOT_10011( .ZN(g25838), .A(II33680) );
  INV_X1 NOT_10012( .ZN(II33683), .A(g24472) );
  INV_X1 NOT_10013( .ZN(g25841), .A(II33683) );
  INV_X1 NOT_10014( .ZN(II33686), .A(g25070) );
  INV_X1 NOT_10015( .ZN(g25844), .A(II33686) );
  INV_X1 NOT_10016( .ZN(II33689), .A(g25074) );
  INV_X1 NOT_10017( .ZN(g25847), .A(II33689) );
  INV_X1 NOT_10018( .ZN(II33692), .A(g24537) );
  INV_X1 NOT_10019( .ZN(g25850), .A(II33692) );
  INV_X1 NOT_10020( .ZN(II33695), .A(g24538) );
  INV_X1 NOT_10021( .ZN(g25851), .A(II33695) );
  INV_X1 NOT_10022( .ZN(II33700), .A(g24474) );
  INV_X1 NOT_10023( .ZN(g25856), .A(II33700) );
  INV_X1 NOT_10024( .ZN(II33703), .A(g24545) );
  INV_X1 NOT_10025( .ZN(g25859), .A(II33703) );
  INV_X1 NOT_10026( .ZN(g25860), .A(g24630) );
  INV_X1 NOT_10027( .ZN(II33708), .A(g24475) );
  INV_X1 NOT_10028( .ZN(g25862), .A(II33708) );
  INV_X1 NOT_10029( .ZN(II33711), .A(g25073) );
  INV_X1 NOT_10030( .ZN(g25865), .A(II33711) );
  INV_X1 NOT_10031( .ZN(II33714), .A(g24547) );
  INV_X1 NOT_10032( .ZN(g25868), .A(II33714) );
  INV_X1 NOT_10033( .ZN(II33717), .A(g24548) );
  INV_X1 NOT_10034( .ZN(g25869), .A(II33717) );
  INV_X1 NOT_10035( .ZN(II33723), .A(g24477) );
  INV_X1 NOT_10036( .ZN(g25877), .A(II33723) );
  INV_X1 NOT_10037( .ZN(II33726), .A(g24557) );
  INV_X1 NOT_10038( .ZN(g25880), .A(II33726) );
  INV_X1 NOT_10039( .ZN(II33732), .A(g24473) );
  INV_X1 NOT_10040( .ZN(g25886), .A(II33732) );
  INV_X1 NOT_10041( .ZN(II33737), .A(g24476) );
  INV_X1 NOT_10042( .ZN(g25891), .A(II33737) );
  INV_X1 NOT_10043( .ZN(g25895), .A(g24939) );
  INV_X1 NOT_10044( .ZN(g25899), .A(g24928) );
  INV_X1 NOT_10045( .ZN(g25903), .A(g24950) );
  INV_X1 NOT_10046( .ZN(g25907), .A(g24940) );
  INV_X1 NOT_10047( .ZN(g25911), .A(g24962) );
  INV_X1 NOT_10048( .ZN(g25915), .A(g24951) );
  INV_X1 NOT_10049( .ZN(g25919), .A(g24973) );
  INV_X1 NOT_10050( .ZN(g25923), .A(g24963) );
  INV_X1 NOT_10051( .ZN(g25937), .A(g24763) );
  INV_X1 NOT_10052( .ZN(g25939), .A(g24784) );
  INV_X1 NOT_10053( .ZN(g25942), .A(g24805) );
  INV_X1 NOT_10054( .ZN(g25945), .A(g24827) );
  INV_X1 NOT_10055( .ZN(g25952), .A(g24735) );
  INV_X1 NOT_10056( .ZN(II33790), .A(g25103) );
  INV_X1 NOT_10057( .ZN(g25976), .A(II33790) );
  INV_X1 NOT_10058( .ZN(II33798), .A(g25109) );
  INV_X1 NOT_10059( .ZN(g25982), .A(II33798) );
  INV_X1 NOT_10060( .ZN(II33801), .A(g25327) );
  INV_X1 NOT_10061( .ZN(g25983), .A(II33801) );
  INV_X1 NOT_10062( .ZN(II33804), .A(g25976) );
  INV_X1 NOT_10063( .ZN(g25984), .A(II33804) );
  INV_X1 NOT_10064( .ZN(II33807), .A(g25588) );
  INV_X1 NOT_10065( .ZN(g25985), .A(II33807) );
  INV_X1 NOT_10066( .ZN(II33810), .A(g25646) );
  INV_X1 NOT_10067( .ZN(g25986), .A(II33810) );
  INV_X1 NOT_10068( .ZN(II33813), .A(g25706) );
  INV_X1 NOT_10069( .ZN(g25987), .A(II33813) );
  INV_X1 NOT_10070( .ZN(II33816), .A(g25647) );
  INV_X1 NOT_10071( .ZN(g25988), .A(II33816) );
  INV_X1 NOT_10072( .ZN(II33819), .A(g25707) );
  INV_X1 NOT_10073( .ZN(g25989), .A(II33819) );
  INV_X1 NOT_10074( .ZN(II33822), .A(g25770) );
  INV_X1 NOT_10075( .ZN(g25990), .A(II33822) );
  INV_X1 NOT_10076( .ZN(II33825), .A(g25462) );
  INV_X1 NOT_10077( .ZN(g25991), .A(II33825) );
  INV_X1 NOT_10078( .ZN(II33828), .A(g25336) );
  INV_X1 NOT_10079( .ZN(g25992), .A(II33828) );
  INV_X1 NOT_10080( .ZN(II33831), .A(g25982) );
  INV_X1 NOT_10081( .ZN(g25993), .A(II33831) );
  INV_X1 NOT_10082( .ZN(II33834), .A(g25667) );
  INV_X1 NOT_10083( .ZN(g25994), .A(II33834) );
  INV_X1 NOT_10084( .ZN(II33837), .A(g25723) );
  INV_X1 NOT_10085( .ZN(g25995), .A(II33837) );
  INV_X1 NOT_10086( .ZN(II33840), .A(g25779) );
  INV_X1 NOT_10087( .ZN(g25996), .A(II33840) );
  INV_X1 NOT_10088( .ZN(II33843), .A(g25724) );
  INV_X1 NOT_10089( .ZN(g25997), .A(II33843) );
  INV_X1 NOT_10090( .ZN(II33846), .A(g25780) );
  INV_X1 NOT_10091( .ZN(g25998), .A(II33846) );
  INV_X1 NOT_10092( .ZN(II33849), .A(g25824) );
  INV_X1 NOT_10093( .ZN(g25999), .A(II33849) );
  INV_X1 NOT_10094( .ZN(II33852), .A(g25471) );
  INV_X1 NOT_10095( .ZN(g26000), .A(II33852) );
  INV_X1 NOT_10096( .ZN(II33855), .A(g25350) );
  INV_X1 NOT_10097( .ZN(g26001), .A(II33855) );
  INV_X1 NOT_10098( .ZN(II33858), .A(g25179) );
  INV_X1 NOT_10099( .ZN(g26002), .A(II33858) );
  INV_X1 NOT_10100( .ZN(II33861), .A(g25744) );
  INV_X1 NOT_10101( .ZN(g26003), .A(II33861) );
  INV_X1 NOT_10102( .ZN(II33864), .A(g25796) );
  INV_X1 NOT_10103( .ZN(g26004), .A(II33864) );
  INV_X1 NOT_10104( .ZN(II33867), .A(g25833) );
  INV_X1 NOT_10105( .ZN(g26005), .A(II33867) );
  INV_X1 NOT_10106( .ZN(II33870), .A(g25797) );
  INV_X1 NOT_10107( .ZN(g26006), .A(II33870) );
  INV_X1 NOT_10108( .ZN(II33873), .A(g25834) );
  INV_X1 NOT_10109( .ZN(g26007), .A(II33873) );
  INV_X1 NOT_10110( .ZN(II33876), .A(g25859) );
  INV_X1 NOT_10111( .ZN(g26008), .A(II33876) );
  INV_X1 NOT_10112( .ZN(II33879), .A(g25488) );
  INV_X1 NOT_10113( .ZN(g26009), .A(II33879) );
  INV_X1 NOT_10114( .ZN(II33882), .A(g25364) );
  INV_X1 NOT_10115( .ZN(g26010), .A(II33882) );
  INV_X1 NOT_10116( .ZN(II33885), .A(g25180) );
  INV_X1 NOT_10117( .ZN(g26011), .A(II33885) );
  INV_X4 NOT_10118( .ZN(II33888), .A(g25817) );
  INV_X4 NOT_10119( .ZN(g26012), .A(II33888) );
  INV_X1 NOT_10120( .ZN(II33891), .A(g25850) );
  INV_X1 NOT_10121( .ZN(g26013), .A(II33891) );
  INV_X1 NOT_10122( .ZN(II33894), .A(g25868) );
  INV_X1 NOT_10123( .ZN(g26014), .A(II33894) );
  INV_X1 NOT_10124( .ZN(II33897), .A(g25851) );
  INV_X1 NOT_10125( .ZN(g26015), .A(II33897) );
  INV_X1 NOT_10126( .ZN(II33900), .A(g25869) );
  INV_X1 NOT_10127( .ZN(g26016), .A(II33900) );
  INV_X1 NOT_10128( .ZN(II33903), .A(g25880) );
  INV_X1 NOT_10129( .ZN(g26017), .A(II33903) );
  INV_X1 NOT_10130( .ZN(II33906), .A(g25519) );
  INV_X1 NOT_10131( .ZN(g26018), .A(II33906) );
  INV_X1 NOT_10132( .ZN(II33909), .A(g25886) );
  INV_X1 NOT_10133( .ZN(g26019), .A(II33909) );
  INV_X1 NOT_10134( .ZN(II33912), .A(g25891) );
  INV_X1 NOT_10135( .ZN(g26020), .A(II33912) );
  INV_X1 NOT_10136( .ZN(II33915), .A(g25762) );
  INV_X1 NOT_10137( .ZN(g26021), .A(II33915) );
  INV_X1 NOT_10138( .ZN(II33918), .A(g25763) );
  INV_X1 NOT_10139( .ZN(g26022), .A(II33918) );
  INV_X1 NOT_10140( .ZN(II33954), .A(g25343) );
  INV_X1 NOT_10141( .ZN(g26056), .A(II33954) );
  INV_X1 NOT_10142( .ZN(II33961), .A(g25357) );
  INV_X1 NOT_10143( .ZN(g26063), .A(II33961) );
  INV_X1 NOT_10144( .ZN(II33968), .A(g25372) );
  INV_X1 NOT_10145( .ZN(g26070), .A(II33968) );
  INV_X1 NOT_10146( .ZN(II33974), .A(g25389) );
  INV_X1 NOT_10147( .ZN(g26076), .A(II33974) );
  INV_X1 NOT_10148( .ZN(II33984), .A(g25932) );
  INV_X1 NOT_10149( .ZN(g26086), .A(II33984) );
  INV_X1 NOT_10150( .ZN(II33990), .A(g25870) );
  INV_X1 NOT_10151( .ZN(g26092), .A(II33990) );
  INV_X1 NOT_10152( .ZN(II33995), .A(g25935) );
  INV_X1 NOT_10153( .ZN(g26102), .A(II33995) );
  INV_X1 NOT_10154( .ZN(II33999), .A(g25490) );
  INV_X1 NOT_10155( .ZN(g26104), .A(II33999) );
  INV_X1 NOT_10156( .ZN(II34002), .A(g25490) );
  INV_X1 NOT_10157( .ZN(g26105), .A(II34002) );
  INV_X1 NOT_10158( .ZN(II34009), .A(g25882) );
  INV_X1 NOT_10159( .ZN(g26114), .A(II34009) );
  INV_X1 NOT_10160( .ZN(II34012), .A(g25938) );
  INV_X1 NOT_10161( .ZN(g26118), .A(II34012) );
  INV_X1 NOT_10162( .ZN(II34017), .A(g25887) );
  INV_X1 NOT_10163( .ZN(g26121), .A(II34017) );
  INV_X1 NOT_10164( .ZN(II34020), .A(g25940) );
  INV_X1 NOT_10165( .ZN(g26125), .A(II34020) );
  INV_X1 NOT_10166( .ZN(II34026), .A(g25892) );
  INV_X1 NOT_10167( .ZN(g26131), .A(II34026) );
  INV_X1 NOT_10168( .ZN(II34029), .A(g25520) );
  INV_X1 NOT_10169( .ZN(g26135), .A(II34029) );
  INV_X1 NOT_10170( .ZN(II34032), .A(g25520) );
  INV_X1 NOT_10171( .ZN(g26136), .A(II34032) );
  INV_X1 NOT_10172( .ZN(II34041), .A(g25566) );
  INV_X1 NOT_10173( .ZN(g26149), .A(II34041) );
  INV_X1 NOT_10174( .ZN(II34044), .A(g25566) );
  INV_X1 NOT_10175( .ZN(g26150), .A(II34044) );
  INV_X1 NOT_10176( .ZN(II34051), .A(g25204) );
  INV_X1 NOT_10177( .ZN(g26159), .A(II34051) );
  INV_X1 NOT_10178( .ZN(II34056), .A(g25206) );
  INV_X1 NOT_10179( .ZN(g26164), .A(II34056) );
  INV_X1 NOT_10180( .ZN(II34059), .A(g25207) );
  INV_X1 NOT_10181( .ZN(g26165), .A(II34059) );
  INV_X1 NOT_10182( .ZN(II34063), .A(g25209) );
  INV_X1 NOT_10183( .ZN(g26167), .A(II34063) );
  INV_X1 NOT_10184( .ZN(II34068), .A(g25211) );
  INV_X1 NOT_10185( .ZN(g26172), .A(II34068) );
  INV_X1 NOT_10186( .ZN(II34071), .A(g25212) );
  INV_X1 NOT_10187( .ZN(g26173), .A(II34071) );
  INV_X1 NOT_10188( .ZN(II34074), .A(g25213) );
  INV_X1 NOT_10189( .ZN(g26174), .A(II34074) );
  INV_X1 NOT_10190( .ZN(II34077), .A(g25954) );
  INV_X1 NOT_10191( .ZN(g26175), .A(II34077) );
  INV_X1 NOT_10192( .ZN(II34080), .A(g25539) );
  INV_X1 NOT_10193( .ZN(g26178), .A(II34080) );
  INV_X1 NOT_10194( .ZN(II34083), .A(g25214) );
  INV_X1 NOT_10195( .ZN(g26181), .A(II34083) );
  INV_X1 NOT_10196( .ZN(II34086), .A(g25215) );
  INV_X1 NOT_10197( .ZN(g26182), .A(II34086) );
  INV_X1 NOT_10198( .ZN(II34091), .A(g25217) );
  INV_X1 NOT_10199( .ZN(g26187), .A(II34091) );
  INV_X1 NOT_10200( .ZN(g26189), .A(g25952) );
  INV_X1 NOT_10201( .ZN(II34096), .A(g25218) );
  INV_X1 NOT_10202( .ZN(g26190), .A(II34096) );
  INV_X1 NOT_10203( .ZN(II34099), .A(g25219) );
  INV_X1 NOT_10204( .ZN(g26191), .A(II34099) );
  INV_X1 NOT_10205( .ZN(II34102), .A(g25220) );
  INV_X1 NOT_10206( .ZN(g26192), .A(II34102) );
  INV_X1 NOT_10207( .ZN(II34105), .A(g25221) );
  INV_X1 NOT_10208( .ZN(g26193), .A(II34105) );
  INV_X1 NOT_10209( .ZN(II34108), .A(g25222) );
  INV_X1 NOT_10210( .ZN(g26194), .A(II34108) );
  INV_X1 NOT_10211( .ZN(II34111), .A(g25223) );
  INV_X1 NOT_10212( .ZN(g26195), .A(II34111) );
  INV_X1 NOT_10213( .ZN(II34114), .A(g25958) );
  INV_X1 NOT_10214( .ZN(g26196), .A(II34114) );
  INV_X1 NOT_10215( .ZN(II34118), .A(g25605) );
  INV_X1 NOT_10216( .ZN(g26202), .A(II34118) );
  INV_X1 NOT_10217( .ZN(II34121), .A(g25224) );
  INV_X1 NOT_10218( .ZN(g26205), .A(II34121) );
  INV_X1 NOT_10219( .ZN(II34124), .A(g25225) );
  INV_X1 NOT_10220( .ZN(g26206), .A(II34124) );
  INV_X1 NOT_10221( .ZN(II34128), .A(g25227) );
  INV_X1 NOT_10222( .ZN(g26208), .A(II34128) );
  INV_X1 NOT_10223( .ZN(g26209), .A(g25296) );
  INV_X1 NOT_10224( .ZN(II34132), .A(g25228) );
  INV_X1 NOT_10225( .ZN(g26210), .A(II34132) );
  INV_X1 NOT_10226( .ZN(II34135), .A(g25229) );
  INV_X1 NOT_10227( .ZN(g26211), .A(II34135) );
  INV_X1 NOT_10228( .ZN(II34140), .A(g25230) );
  INV_X1 NOT_10229( .ZN(g26214), .A(II34140) );
  INV_X1 NOT_10230( .ZN(II34143), .A(g25231) );
  INV_X1 NOT_10231( .ZN(g26215), .A(II34143) );
  INV_X1 NOT_10232( .ZN(II34146), .A(g25232) );
  INV_X1 NOT_10233( .ZN(g26216), .A(II34146) );
  INV_X1 NOT_10234( .ZN(II34150), .A(g25233) );
  INV_X4 NOT_10235( .ZN(g26220), .A(II34150) );
  INV_X4 NOT_10236( .ZN(II34153), .A(g25234) );
  INV_X1 NOT_10237( .ZN(g26221), .A(II34153) );
  INV_X1 NOT_10238( .ZN(II34156), .A(g25235) );
  INV_X1 NOT_10239( .ZN(g26222), .A(II34156) );
  INV_X1 NOT_10240( .ZN(II34159), .A(g25964) );
  INV_X1 NOT_10241( .ZN(g26223), .A(II34159) );
  INV_X1 NOT_10242( .ZN(II34162), .A(g25684) );
  INV_X1 NOT_10243( .ZN(g26226), .A(II34162) );
  INV_X1 NOT_10244( .ZN(II34165), .A(g25236) );
  INV_X1 NOT_10245( .ZN(g26229), .A(II34165) );
  INV_X1 NOT_10246( .ZN(II34168), .A(g25237) );
  INV_X1 NOT_10247( .ZN(g26230), .A(II34168) );
  INV_X1 NOT_10248( .ZN(II34172), .A(g25239) );
  INV_X1 NOT_10249( .ZN(g26232), .A(II34172) );
  INV_X1 NOT_10250( .ZN(g26237), .A(g25306) );
  INV_X1 NOT_10251( .ZN(II34180), .A(g25240) );
  INV_X1 NOT_10252( .ZN(g26238), .A(II34180) );
  INV_X1 NOT_10253( .ZN(II34183), .A(g25241) );
  INV_X1 NOT_10254( .ZN(g26239), .A(II34183) );
  INV_X1 NOT_10255( .ZN(II34189), .A(g25242) );
  INV_X1 NOT_10256( .ZN(g26245), .A(II34189) );
  INV_X1 NOT_10257( .ZN(II34192), .A(g25243) );
  INV_X1 NOT_10258( .ZN(g26246), .A(II34192) );
  INV_X1 NOT_10259( .ZN(II34195), .A(g25244) );
  INV_X1 NOT_10260( .ZN(g26247), .A(II34195) );
  INV_X1 NOT_10261( .ZN(II34198), .A(g25245) );
  INV_X1 NOT_10262( .ZN(g26248), .A(II34198) );
  INV_X1 NOT_10263( .ZN(II34201), .A(g25246) );
  INV_X1 NOT_10264( .ZN(g26249), .A(II34201) );
  INV_X1 NOT_10265( .ZN(II34204), .A(g25247) );
  INV_X1 NOT_10266( .ZN(g26250), .A(II34204) );
  INV_X1 NOT_10267( .ZN(II34207), .A(g25969) );
  INV_X1 NOT_10268( .ZN(g26251), .A(II34207) );
  INV_X1 NOT_10269( .ZN(II34210), .A(g25761) );
  INV_X1 NOT_10270( .ZN(g26254), .A(II34210) );
  INV_X1 NOT_10271( .ZN(II34220), .A(g25248) );
  INV_X1 NOT_10272( .ZN(g26264), .A(II34220) );
  INV_X1 NOT_10273( .ZN(g26275), .A(g25315) );
  INV_X1 NOT_10274( .ZN(II34230), .A(g25249) );
  INV_X1 NOT_10275( .ZN(g26276), .A(II34230) );
  INV_X1 NOT_10276( .ZN(II34233), .A(g25250) );
  INV_X1 NOT_10277( .ZN(g26277), .A(II34233) );
  INV_X1 NOT_10278( .ZN(II34238), .A(g25251) );
  INV_X1 NOT_10279( .ZN(g26280), .A(II34238) );
  INV_X1 NOT_10280( .ZN(II34241), .A(g25252) );
  INV_X1 NOT_10281( .ZN(g26281), .A(II34241) );
  INV_X1 NOT_10282( .ZN(II34244), .A(g25253) );
  INV_X1 NOT_10283( .ZN(g26282), .A(II34244) );
  INV_X1 NOT_10284( .ZN(II34254), .A(g25185) );
  INV_X1 NOT_10285( .ZN(g26294), .A(II34254) );
  INV_X1 NOT_10286( .ZN(II34266), .A(g25255) );
  INV_X1 NOT_10287( .ZN(g26308), .A(II34266) );
  INV_X1 NOT_10288( .ZN(g26313), .A(g25324) );
  INV_X1 NOT_10289( .ZN(II34274), .A(g25256) );
  INV_X1 NOT_10290( .ZN(g26314), .A(II34274) );
  INV_X1 NOT_10291( .ZN(II34277), .A(g25257) );
  INV_X1 NOT_10292( .ZN(g26315), .A(II34277) );
  INV_X1 NOT_10293( .ZN(II34296), .A(g25189) );
  INV_X1 NOT_10294( .ZN(g26341), .A(II34296) );
  INV_X1 NOT_10295( .ZN(II34306), .A(g25259) );
  INV_X1 NOT_10296( .ZN(g26349), .A(II34306) );
  INV_X1 NOT_10297( .ZN(II34313), .A(g25265) );
  INV_X1 NOT_10298( .ZN(g26354), .A(II34313) );
  INV_X1 NOT_10299( .ZN(II34316), .A(g25191) );
  INV_X1 NOT_10300( .ZN(g26355), .A(II34316) );
  INV_X1 NOT_10301( .ZN(II34321), .A(g25928) );
  INV_X1 NOT_10302( .ZN(g26358), .A(II34321) );
  INV_X1 NOT_10303( .ZN(II34327), .A(g25260) );
  INV_X1 NOT_10304( .ZN(g26364), .A(II34327) );
  INV_X1 NOT_10305( .ZN(II34343), .A(g25194) );
  INV_X1 NOT_10306( .ZN(g26385), .A(II34343) );
  INV_X1 NOT_10307( .ZN(II34353), .A(g25927) );
  INV_X1 NOT_10308( .ZN(g26393), .A(II34353) );
  INV_X1 NOT_10309( .ZN(II34358), .A(g25262) );
  INV_X1 NOT_10310( .ZN(g26398), .A(II34358) );
  INV_X1 NOT_10311( .ZN(II34363), .A(g25930) );
  INV_X1 NOT_10312( .ZN(g26401), .A(II34363) );
  INV_X1 NOT_10313( .ZN(II34369), .A(g25263) );
  INV_X1 NOT_10314( .ZN(g26407), .A(II34369) );
  INV_X1 NOT_10315( .ZN(II34385), .A(g25197) );
  INV_X1 NOT_10316( .ZN(g26428), .A(II34385) );
  INV_X1 NOT_10317( .ZN(II34388), .A(g25200) );
  INV_X1 NOT_10318( .ZN(g26429), .A(II34388) );
  INV_X1 NOT_10319( .ZN(II34392), .A(g25266) );
  INV_X1 NOT_10320( .ZN(g26433), .A(II34392) );
  INV_X1 NOT_10321( .ZN(II34395), .A(g25929) );
  INV_X1 NOT_10322( .ZN(g26434), .A(II34395) );
  INV_X1 NOT_10323( .ZN(II34400), .A(g25267) );
  INV_X1 NOT_10324( .ZN(g26439), .A(II34400) );
  INV_X1 NOT_10325( .ZN(II34405), .A(g25933) );
  INV_X1 NOT_10326( .ZN(g26442), .A(II34405) );
  INV_X1 NOT_10327( .ZN(II34411), .A(g25268) );
  INV_X1 NOT_10328( .ZN(g26448), .A(II34411) );
  INV_X1 NOT_10329( .ZN(II34421), .A(g25203) );
  INV_X1 NOT_10330( .ZN(g26461), .A(II34421) );
  INV_X1 NOT_10331( .ZN(II34425), .A(g25270) );
  INV_X1 NOT_10332( .ZN(g26465), .A(II34425) );
  INV_X1 NOT_10333( .ZN(II34428), .A(g25931) );
  INV_X1 NOT_10334( .ZN(g26466), .A(II34428) );
  INV_X1 NOT_10335( .ZN(II34433), .A(g25271) );
  INV_X1 NOT_10336( .ZN(g26471), .A(II34433) );
  INV_X1 NOT_10337( .ZN(II34438), .A(g25936) );
  INV_X1 NOT_10338( .ZN(g26474), .A(II34438) );
  INV_X1 NOT_10339( .ZN(II34444), .A(g25272) );
  INV_X1 NOT_10340( .ZN(g26480), .A(II34444) );
  INV_X1 NOT_10341( .ZN(g26481), .A(g25764) );
  INV_X1 NOT_10342( .ZN(II34449), .A(g25205) );
  INV_X1 NOT_10343( .ZN(g26485), .A(II34449) );
  INV_X1 NOT_10344( .ZN(II34453), .A(g25279) );
  INV_X1 NOT_10345( .ZN(g26489), .A(II34453) );
  INV_X4 NOT_10346( .ZN(II34456), .A(g25934) );
  INV_X4 NOT_10347( .ZN(g26490), .A(II34456) );
  INV_X1 NOT_10348( .ZN(II34461), .A(g25280) );
  INV_X1 NOT_10349( .ZN(g26495), .A(II34461) );
  INV_X1 NOT_10350( .ZN(II34464), .A(g25199) );
  INV_X1 NOT_10351( .ZN(g26496), .A(II34464) );
  INV_X1 NOT_10352( .ZN(g26497), .A(g25818) );
  INV_X1 NOT_10353( .ZN(II34469), .A(g25210) );
  INV_X1 NOT_10354( .ZN(g26501), .A(II34469) );
  INV_X1 NOT_10355( .ZN(II34473), .A(g25288) );
  INV_X1 NOT_10356( .ZN(g26505), .A(II34473) );
  INV_X1 NOT_10357( .ZN(II34476), .A(g25201) );
  INV_X1 NOT_10358( .ZN(g26506), .A(II34476) );
  INV_X1 NOT_10359( .ZN(II34479), .A(g25202) );
  INV_X1 NOT_10360( .ZN(g26507), .A(II34479) );
  INV_X1 NOT_10361( .ZN(g26508), .A(g25312) );
  INV_X1 NOT_10362( .ZN(g26512), .A(g25853) );
  INV_X1 NOT_10363( .ZN(g26516), .A(g25320) );
  INV_X1 NOT_10364( .ZN(g26520), .A(g25874) );
  INV_X1 NOT_10365( .ZN(g26521), .A(g25331) );
  INV_X1 NOT_10366( .ZN(g26525), .A(g25340) );
  INV_X1 NOT_10367( .ZN(g26533), .A(g25454) );
  INV_X1 NOT_10368( .ZN(g26538), .A(g25458) );
  INV_X1 NOT_10369( .ZN(g26539), .A(g25463) );
  INV_X1 NOT_10370( .ZN(g26540), .A(g25467) );
  INV_X1 NOT_10371( .ZN(g26542), .A(g25472) );
  INV_X1 NOT_10372( .ZN(g26543), .A(g25476) );
  INV_X1 NOT_10373( .ZN(g26544), .A(g25479) );
  INV_X1 NOT_10374( .ZN(g26546), .A(g25484) );
  INV_X1 NOT_10375( .ZN(II34505), .A(g25450) );
  INV_X1 NOT_10376( .ZN(g26548), .A(II34505) );
  INV_X1 NOT_10377( .ZN(g26549), .A(g25421) );
  INV_X1 NOT_10378( .ZN(g26550), .A(g25493) );
  INV_X1 NOT_10379( .ZN(g26551), .A(g25496) );
  INV_X1 NOT_10380( .ZN(g26552), .A(g25499) );
  INV_X1 NOT_10381( .ZN(g26554), .A(g25502) );
  INV_X1 NOT_10382( .ZN(g26555), .A(g25507) );
  INV_X1 NOT_10383( .ZN(g26556), .A(g25510) );
  INV_X1 NOT_10384( .ZN(g26558), .A(g25515) );
  INV_X1 NOT_10385( .ZN(g26561), .A(g25524) );
  INV_X1 NOT_10386( .ZN(g26562), .A(g25527) );
  INV_X1 NOT_10387( .ZN(g26563), .A(g25530) );
  INV_X1 NOT_10388( .ZN(g26564), .A(g25533) );
  INV_X1 NOT_10389( .ZN(g26565), .A(g25536) );
  INV_X1 NOT_10390( .ZN(g26566), .A(g25540) );
  INV_X1 NOT_10391( .ZN(g26567), .A(g25543) );
  INV_X1 NOT_10392( .ZN(g26568), .A(g25546) );
  INV_X1 NOT_10393( .ZN(g26570), .A(g25549) );
  INV_X1 NOT_10394( .ZN(g26571), .A(g25554) );
  INV_X1 NOT_10395( .ZN(g26572), .A(g25557) );
  INV_X1 NOT_10396( .ZN(g26574), .A(g25562) );
  INV_X1 NOT_10397( .ZN(II34535), .A(g25451) );
  INV_X1 NOT_10398( .ZN(g26576), .A(II34535) );
  INV_X1 NOT_10399( .ZN(g26577), .A(g25436) );
  INV_X1 NOT_10400( .ZN(g26578), .A(g25573) );
  INV_X1 NOT_10401( .ZN(g26579), .A(g25576) );
  INV_X1 NOT_10402( .ZN(g26580), .A(g25579) );
  INV_X1 NOT_10403( .ZN(g26581), .A(g25582) );
  INV_X1 NOT_10404( .ZN(g26582), .A(g25585) );
  INV_X1 NOT_10405( .ZN(g26584), .A(g25590) );
  INV_X1 NOT_10406( .ZN(g26585), .A(g25593) );
  INV_X1 NOT_10407( .ZN(g26586), .A(g25596) );
  INV_X1 NOT_10408( .ZN(g26587), .A(g25599) );
  INV_X1 NOT_10409( .ZN(g26588), .A(g25602) );
  INV_X1 NOT_10410( .ZN(g26589), .A(g25606) );
  INV_X1 NOT_10411( .ZN(g26590), .A(g25609) );
  INV_X1 NOT_10412( .ZN(g26591), .A(g25612) );
  INV_X1 NOT_10413( .ZN(g26593), .A(g25615) );
  INV_X1 NOT_10414( .ZN(g26594), .A(g25620) );
  INV_X1 NOT_10415( .ZN(g26595), .A(g25623) );
  INV_X1 NOT_10416( .ZN(g26597), .A(g25443) );
  INV_X1 NOT_10417( .ZN(g26598), .A(g25634) );
  INV_X1 NOT_10418( .ZN(g26599), .A(g25637) );
  INV_X1 NOT_10419( .ZN(g26600), .A(g25640) );
  INV_X1 NOT_10420( .ZN(g26601), .A(g25643) );
  INV_X1 NOT_10421( .ZN(g26602), .A(g25652) );
  INV_X1 NOT_10422( .ZN(g26603), .A(g25655) );
  INV_X1 NOT_10423( .ZN(g26604), .A(g25658) );
  INV_X1 NOT_10424( .ZN(g26605), .A(g25661) );
  INV_X1 NOT_10425( .ZN(g26606), .A(g25664) );
  INV_X1 NOT_10426( .ZN(g26608), .A(g25669) );
  INV_X1 NOT_10427( .ZN(g26609), .A(g25672) );
  INV_X1 NOT_10428( .ZN(g26610), .A(g25675) );
  INV_X1 NOT_10429( .ZN(g26611), .A(g25678) );
  INV_X1 NOT_10430( .ZN(g26612), .A(g25681) );
  INV_X1 NOT_10431( .ZN(g26613), .A(g25685) );
  INV_X1 NOT_10432( .ZN(g26614), .A(g25688) );
  INV_X1 NOT_10433( .ZN(g26615), .A(g25691) );
  INV_X1 NOT_10434( .ZN(g26617), .A(g25694) );
  INV_X1 NOT_10435( .ZN(II34579), .A(g25452) );
  INV_X1 NOT_10436( .ZN(g26618), .A(II34579) );
  INV_X1 NOT_10437( .ZN(g26619), .A(g25700) );
  INV_X1 NOT_10438( .ZN(g26620), .A(g25703) );
  INV_X1 NOT_10439( .ZN(g26621), .A(g25711) );
  INV_X1 NOT_10440( .ZN(g26622), .A(g25714) );
  INV_X1 NOT_10441( .ZN(g26623), .A(g25717) );
  INV_X1 NOT_10442( .ZN(g26624), .A(g25720) );
  INV_X1 NOT_10443( .ZN(g26625), .A(g25729) );
  INV_X1 NOT_10444( .ZN(g26626), .A(g25732) );
  INV_X1 NOT_10445( .ZN(g26627), .A(g25735) );
  INV_X1 NOT_10446( .ZN(g26628), .A(g25738) );
  INV_X1 NOT_10447( .ZN(g26629), .A(g25741) );
  INV_X1 NOT_10448( .ZN(g26631), .A(g25746) );
  INV_X1 NOT_10449( .ZN(g26632), .A(g25749) );
  INV_X1 NOT_10450( .ZN(g26633), .A(g25752) );
  INV_X1 NOT_10451( .ZN(g26634), .A(g25755) );
  INV_X1 NOT_10452( .ZN(g26635), .A(g25758) );
  INV_X1 NOT_10453( .ZN(g26636), .A(g25767) );
  INV_X1 NOT_10454( .ZN(g26637), .A(g25773) );
  INV_X1 NOT_10455( .ZN(g26638), .A(g25776) );
  INV_X1 NOT_10456( .ZN(g26639), .A(g25784) );
  INV_X1 NOT_10457( .ZN(g26640), .A(g25787) );
  INV_X1 NOT_10458( .ZN(g26641), .A(g25790) );
  INV_X1 NOT_10459( .ZN(g26642), .A(g25793) );
  INV_X1 NOT_10460( .ZN(g26643), .A(g25802) );
  INV_X1 NOT_10461( .ZN(g26644), .A(g25805) );
  INV_X4 NOT_10462( .ZN(g26645), .A(g25808) );
  INV_X4 NOT_10463( .ZN(g26646), .A(g25811) );
  INV_X4 NOT_10464( .ZN(g26647), .A(g25814) );
  INV_X1 NOT_10465( .ZN(g26648), .A(g25821) );
  INV_X1 NOT_10466( .ZN(g26649), .A(g25827) );
  INV_X1 NOT_10467( .ZN(g26650), .A(g25830) );
  INV_X1 NOT_10468( .ZN(g26651), .A(g25838) );
  INV_X1 NOT_10469( .ZN(g26652), .A(g25841) );
  INV_X1 NOT_10470( .ZN(g26653), .A(g25844) );
  INV_X1 NOT_10471( .ZN(g26654), .A(g25847) );
  INV_X1 NOT_10472( .ZN(g26656), .A(g25856) );
  INV_X1 NOT_10473( .ZN(g26657), .A(g25862) );
  INV_X1 NOT_10474( .ZN(g26658), .A(g25865) );
  INV_X1 NOT_10475( .ZN(g26662), .A(g25877) );
  INV_X1 NOT_10476( .ZN(II34641), .A(g26086) );
  INV_X1 NOT_10477( .ZN(g26678), .A(II34641) );
  INV_X1 NOT_10478( .ZN(II34644), .A(g26159) );
  INV_X1 NOT_10479( .ZN(g26679), .A(II34644) );
  INV_X1 NOT_10480( .ZN(II34647), .A(g26164) );
  INV_X1 NOT_10481( .ZN(g26680), .A(II34647) );
  INV_X1 NOT_10482( .ZN(II34650), .A(g26172) );
  INV_X1 NOT_10483( .ZN(g26681), .A(II34650) );
  INV_X1 NOT_10484( .ZN(II34653), .A(g26165) );
  INV_X1 NOT_10485( .ZN(g26682), .A(II34653) );
  INV_X1 NOT_10486( .ZN(II34656), .A(g26173) );
  INV_X1 NOT_10487( .ZN(g26683), .A(II34656) );
  INV_X1 NOT_10488( .ZN(II34659), .A(g26190) );
  INV_X1 NOT_10489( .ZN(g26684), .A(II34659) );
  INV_X1 NOT_10490( .ZN(II34662), .A(g26174) );
  INV_X1 NOT_10491( .ZN(g26685), .A(II34662) );
  INV_X1 NOT_10492( .ZN(II34665), .A(g26191) );
  INV_X1 NOT_10493( .ZN(g26686), .A(II34665) );
  INV_X1 NOT_10494( .ZN(II34668), .A(g26210) );
  INV_X1 NOT_10495( .ZN(g26687), .A(II34668) );
  INV_X1 NOT_10496( .ZN(II34671), .A(g26192) );
  INV_X1 NOT_10497( .ZN(g26688), .A(II34671) );
  INV_X1 NOT_10498( .ZN(II34674), .A(g26211) );
  INV_X1 NOT_10499( .ZN(g26689), .A(II34674) );
  INV_X1 NOT_10500( .ZN(II34677), .A(g26232) );
  INV_X1 NOT_10501( .ZN(g26690), .A(II34677) );
  INV_X1 NOT_10502( .ZN(II34680), .A(g26294) );
  INV_X1 NOT_10503( .ZN(g26691), .A(II34680) );
  INV_X1 NOT_10504( .ZN(II34683), .A(g26364) );
  INV_X1 NOT_10505( .ZN(g26692), .A(II34683) );
  INV_X1 NOT_10506( .ZN(II34686), .A(g26398) );
  INV_X1 NOT_10507( .ZN(g26693), .A(II34686) );
  INV_X1 NOT_10508( .ZN(II34689), .A(g26433) );
  INV_X1 NOT_10509( .ZN(g26694), .A(II34689) );
  INV_X1 NOT_10510( .ZN(II34692), .A(g26102) );
  INV_X1 NOT_10511( .ZN(g26695), .A(II34692) );
  INV_X1 NOT_10512( .ZN(II34695), .A(g26167) );
  INV_X1 NOT_10513( .ZN(g26696), .A(II34695) );
  INV_X1 NOT_10514( .ZN(II34698), .A(g26181) );
  INV_X1 NOT_10515( .ZN(g26697), .A(II34698) );
  INV_X1 NOT_10516( .ZN(II34701), .A(g26193) );
  INV_X1 NOT_10517( .ZN(g26698), .A(II34701) );
  INV_X1 NOT_10518( .ZN(II34704), .A(g26182) );
  INV_X1 NOT_10519( .ZN(g26699), .A(II34704) );
  INV_X1 NOT_10520( .ZN(II34707), .A(g26194) );
  INV_X1 NOT_10521( .ZN(g26700), .A(II34707) );
  INV_X1 NOT_10522( .ZN(II34710), .A(g26214) );
  INV_X1 NOT_10523( .ZN(g26701), .A(II34710) );
  INV_X1 NOT_10524( .ZN(II34713), .A(g26195) );
  INV_X1 NOT_10525( .ZN(g26702), .A(II34713) );
  INV_X1 NOT_10526( .ZN(II34716), .A(g26215) );
  INV_X1 NOT_10527( .ZN(g26703), .A(II34716) );
  INV_X1 NOT_10528( .ZN(II34719), .A(g26238) );
  INV_X1 NOT_10529( .ZN(g26704), .A(II34719) );
  INV_X1 NOT_10530( .ZN(II34722), .A(g26216) );
  INV_X1 NOT_10531( .ZN(g26705), .A(II34722) );
  INV_X1 NOT_10532( .ZN(II34725), .A(g26239) );
  INV_X1 NOT_10533( .ZN(g26706), .A(II34725) );
  INV_X1 NOT_10534( .ZN(II34728), .A(g26264) );
  INV_X1 NOT_10535( .ZN(g26707), .A(II34728) );
  INV_X1 NOT_10536( .ZN(II34731), .A(g26341) );
  INV_X1 NOT_10537( .ZN(g26708), .A(II34731) );
  INV_X1 NOT_10538( .ZN(II34734), .A(g26407) );
  INV_X1 NOT_10539( .ZN(g26709), .A(II34734) );
  INV_X1 NOT_10540( .ZN(II34737), .A(g26439) );
  INV_X1 NOT_10541( .ZN(g26710), .A(II34737) );
  INV_X1 NOT_10542( .ZN(II34740), .A(g26465) );
  INV_X1 NOT_10543( .ZN(g26711), .A(II34740) );
  INV_X1 NOT_10544( .ZN(II34743), .A(g26118) );
  INV_X1 NOT_10545( .ZN(g26712), .A(II34743) );
  INV_X1 NOT_10546( .ZN(II34746), .A(g26187) );
  INV_X1 NOT_10547( .ZN(g26713), .A(II34746) );
  INV_X1 NOT_10548( .ZN(II34749), .A(g26205) );
  INV_X1 NOT_10549( .ZN(g26714), .A(II34749) );
  INV_X1 NOT_10550( .ZN(II34752), .A(g26220) );
  INV_X1 NOT_10551( .ZN(g26715), .A(II34752) );
  INV_X1 NOT_10552( .ZN(II34755), .A(g26206) );
  INV_X1 NOT_10553( .ZN(g26716), .A(II34755) );
  INV_X1 NOT_10554( .ZN(II34758), .A(g26221) );
  INV_X1 NOT_10555( .ZN(g26717), .A(II34758) );
  INV_X1 NOT_10556( .ZN(II34761), .A(g26245) );
  INV_X1 NOT_10557( .ZN(g26718), .A(II34761) );
  INV_X1 NOT_10558( .ZN(II34764), .A(g26222) );
  INV_X1 NOT_10559( .ZN(g26719), .A(II34764) );
  INV_X1 NOT_10560( .ZN(II34767), .A(g26246) );
  INV_X1 NOT_10561( .ZN(g26720), .A(II34767) );
  INV_X1 NOT_10562( .ZN(II34770), .A(g26276) );
  INV_X1 NOT_10563( .ZN(g26721), .A(II34770) );
  INV_X1 NOT_10564( .ZN(II34773), .A(g26247) );
  INV_X1 NOT_10565( .ZN(g26722), .A(II34773) );
  INV_X1 NOT_10566( .ZN(II34776), .A(g26277) );
  INV_X1 NOT_10567( .ZN(g26723), .A(II34776) );
  INV_X1 NOT_10568( .ZN(II34779), .A(g26308) );
  INV_X1 NOT_10569( .ZN(g26724), .A(II34779) );
  INV_X1 NOT_10570( .ZN(II34782), .A(g26385) );
  INV_X1 NOT_10571( .ZN(g26725), .A(II34782) );
  INV_X1 NOT_10572( .ZN(II34785), .A(g26448) );
  INV_X1 NOT_10573( .ZN(g26726), .A(II34785) );
  INV_X1 NOT_10574( .ZN(II34788), .A(g26471) );
  INV_X1 NOT_10575( .ZN(g26727), .A(II34788) );
  INV_X1 NOT_10576( .ZN(II34791), .A(g26489) );
  INV_X1 NOT_10577( .ZN(g26728), .A(II34791) );
  INV_X1 NOT_10578( .ZN(II34794), .A(g26125) );
  INV_X1 NOT_10579( .ZN(g26729), .A(II34794) );
  INV_X1 NOT_10580( .ZN(II34797), .A(g26208) );
  INV_X1 NOT_10581( .ZN(g26730), .A(II34797) );
  INV_X1 NOT_10582( .ZN(II34800), .A(g26229) );
  INV_X1 NOT_10583( .ZN(g26731), .A(II34800) );
  INV_X1 NOT_10584( .ZN(II34803), .A(g26248) );
  INV_X1 NOT_10585( .ZN(g26732), .A(II34803) );
  INV_X1 NOT_10586( .ZN(II34806), .A(g26230) );
  INV_X1 NOT_10587( .ZN(g26733), .A(II34806) );
  INV_X1 NOT_10588( .ZN(II34809), .A(g26249) );
  INV_X1 NOT_10589( .ZN(g26734), .A(II34809) );
  INV_X1 NOT_10590( .ZN(II34812), .A(g26280) );
  INV_X1 NOT_10591( .ZN(g26735), .A(II34812) );
  INV_X1 NOT_10592( .ZN(II34815), .A(g26250) );
  INV_X1 NOT_10593( .ZN(g26736), .A(II34815) );
  INV_X1 NOT_10594( .ZN(II34818), .A(g26281) );
  INV_X1 NOT_10595( .ZN(g26737), .A(II34818) );
  INV_X1 NOT_10596( .ZN(II34821), .A(g26314) );
  INV_X1 NOT_10597( .ZN(g26738), .A(II34821) );
  INV_X1 NOT_10598( .ZN(II34824), .A(g26282) );
  INV_X1 NOT_10599( .ZN(g26739), .A(II34824) );
  INV_X1 NOT_10600( .ZN(II34827), .A(g26315) );
  INV_X1 NOT_10601( .ZN(g26740), .A(II34827) );
  INV_X1 NOT_10602( .ZN(II34830), .A(g26349) );
  INV_X1 NOT_10603( .ZN(g26741), .A(II34830) );
  INV_X1 NOT_10604( .ZN(II34833), .A(g26428) );
  INV_X1 NOT_10605( .ZN(g26742), .A(II34833) );
  INV_X1 NOT_10606( .ZN(II34836), .A(g26480) );
  INV_X1 NOT_10607( .ZN(g26743), .A(II34836) );
  INV_X1 NOT_10608( .ZN(II34839), .A(g26495) );
  INV_X1 NOT_10609( .ZN(g26744), .A(II34839) );
  INV_X1 NOT_10610( .ZN(II34842), .A(g26505) );
  INV_X1 NOT_10611( .ZN(g26745), .A(II34842) );
  INV_X1 NOT_10612( .ZN(II34845), .A(g26496) );
  INV_X1 NOT_10613( .ZN(g26746), .A(II34845) );
  INV_X1 NOT_10614( .ZN(II34848), .A(g26506) );
  INV_X1 NOT_10615( .ZN(g26747), .A(II34848) );
  INV_X1 NOT_10616( .ZN(II34851), .A(g26354) );
  INV_X1 NOT_10617( .ZN(g26748), .A(II34851) );
  INV_X1 NOT_10618( .ZN(II34854), .A(g26507) );
  INV_X1 NOT_10619( .ZN(g26749), .A(II34854) );
  INV_X1 NOT_10620( .ZN(II34857), .A(g26355) );
  INV_X1 NOT_10621( .ZN(g26750), .A(II34857) );
  INV_X1 NOT_10622( .ZN(II34860), .A(g26548) );
  INV_X1 NOT_10623( .ZN(g26751), .A(II34860) );
  INV_X1 NOT_10624( .ZN(II34863), .A(g26576) );
  INV_X1 NOT_10625( .ZN(g26752), .A(II34863) );
  INV_X1 NOT_10626( .ZN(II34866), .A(g26618) );
  INV_X1 NOT_10627( .ZN(g26753), .A(II34866) );
  INV_X1 NOT_10628( .ZN(II34872), .A(g26217) );
  INV_X1 NOT_10629( .ZN(g26757), .A(II34872) );
  INV_X1 NOT_10630( .ZN(II34879), .A(g26240) );
  INV_X1 NOT_10631( .ZN(g26762), .A(II34879) );
  INV_X1 NOT_10632( .ZN(II34901), .A(g26295) );
  INV_X1 NOT_10633( .ZN(g26782), .A(II34901) );
  INV_X1 NOT_10634( .ZN(II34909), .A(g26265) );
  INV_X1 NOT_10635( .ZN(g26788), .A(II34909) );
  INV_X1 NOT_10636( .ZN(II34916), .A(g26240) );
  INV_X1 NOT_10637( .ZN(g26793), .A(II34916) );
  INV_X1 NOT_10638( .ZN(II34921), .A(g26217) );
  INV_X4 NOT_10639( .ZN(g26796), .A(II34921) );
  INV_X4 NOT_10640( .ZN(II34946), .A(g26534) );
  INV_X1 NOT_10641( .ZN(g26819), .A(II34946) );
  INV_X1 NOT_10642( .ZN(II34957), .A(g26541) );
  INV_X1 NOT_10643( .ZN(g26828), .A(II34957) );
  INV_X1 NOT_10644( .ZN(II34961), .A(g26545) );
  INV_X1 NOT_10645( .ZN(g26830), .A(II34961) );
  INV_X1 NOT_10646( .ZN(II34964), .A(g26547) );
  INV_X1 NOT_10647( .ZN(g26831), .A(II34964) );
  INV_X1 NOT_10648( .ZN(II34967), .A(g26553) );
  INV_X1 NOT_10649( .ZN(g26832), .A(II34967) );
  INV_X1 NOT_10650( .ZN(II34971), .A(g26557) );
  INV_X1 NOT_10651( .ZN(g26834), .A(II34971) );
  INV_X1 NOT_10652( .ZN(II34974), .A(g26168) );
  INV_X1 NOT_10653( .ZN(g26835), .A(II34974) );
  INV_X1 NOT_10654( .ZN(II34977), .A(g26559) );
  INV_X1 NOT_10655( .ZN(g26836), .A(II34977) );
  INV_X1 NOT_10656( .ZN(II34980), .A(g26458) );
  INV_X1 NOT_10657( .ZN(g26837), .A(II34980) );
  INV_X1 NOT_10658( .ZN(II34983), .A(g26569) );
  INV_X1 NOT_10659( .ZN(g26840), .A(II34983) );
  INV_X1 NOT_10660( .ZN(II34986), .A(g26160) );
  INV_X1 NOT_10661( .ZN(g26841), .A(II34986) );
  INV_X1 NOT_10662( .ZN(II34990), .A(g26573) );
  INV_X1 NOT_10663( .ZN(g26843), .A(II34990) );
  INV_X1 NOT_10664( .ZN(II34993), .A(g26575) );
  INV_X1 NOT_10665( .ZN(g26844), .A(II34993) );
  INV_X1 NOT_10666( .ZN(II34997), .A(g26482) );
  INV_X1 NOT_10667( .ZN(g26846), .A(II34997) );
  INV_X1 NOT_10668( .ZN(II35000), .A(g26336) );
  INV_X1 NOT_10669( .ZN(g26849), .A(II35000) );
  INV_X1 NOT_10670( .ZN(II35003), .A(g26592) );
  INV_X1 NOT_10671( .ZN(g26850), .A(II35003) );
  INV_X1 NOT_10672( .ZN(II35007), .A(g26596) );
  INV_X1 NOT_10673( .ZN(g26852), .A(II35007) );
  INV_X1 NOT_10674( .ZN(II35011), .A(g26304) );
  INV_X1 NOT_10675( .ZN(g26854), .A(II35011) );
  INV_X1 NOT_10676( .ZN(II35014), .A(g26498) );
  INV_X1 NOT_10677( .ZN(g26855), .A(II35014) );
  INV_X1 NOT_10678( .ZN(II35017), .A(g26616) );
  INV_X1 NOT_10679( .ZN(g26858), .A(II35017) );
  INV_X1 NOT_10680( .ZN(II35028), .A(g26513) );
  INV_X1 NOT_10681( .ZN(g26861), .A(II35028) );
  INV_X1 NOT_10682( .ZN(II35031), .A(g26529) );
  INV_X1 NOT_10683( .ZN(g26864), .A(II35031) );
  INV_X1 NOT_10684( .ZN(II35049), .A(g26530) );
  INV_X1 NOT_10685( .ZN(g26868), .A(II35049) );
  INV_X1 NOT_10686( .ZN(II35053), .A(g26655) );
  INV_X1 NOT_10687( .ZN(g26872), .A(II35053) );
  INV_X1 NOT_10688( .ZN(II35064), .A(g26531) );
  INV_X1 NOT_10689( .ZN(g26875), .A(II35064) );
  INV_X1 NOT_10690( .ZN(II35067), .A(g26659) );
  INV_X1 NOT_10691( .ZN(g26876), .A(II35067) );
  INV_X1 NOT_10692( .ZN(II35072), .A(g26661) );
  INV_X1 NOT_10693( .ZN(g26881), .A(II35072) );
  INV_X1 NOT_10694( .ZN(II35076), .A(g26532) );
  INV_X1 NOT_10695( .ZN(g26883), .A(II35076) );
  INV_X1 NOT_10696( .ZN(II35079), .A(g26664) );
  INV_X1 NOT_10697( .ZN(g26884), .A(II35079) );
  INV_X1 NOT_10698( .ZN(II35083), .A(g26665) );
  INV_X4 NOT_10699( .ZN(g26886), .A(II35083) );
  INV_X1 NOT_10700( .ZN(II35087), .A(g26667) );
  INV_X1 NOT_10701( .ZN(g26890), .A(II35087) );
  INV_X1 NOT_10702( .ZN(II35092), .A(g26669) );
  INV_X1 NOT_10703( .ZN(g26895), .A(II35092) );
  INV_X1 NOT_10704( .ZN(II35095), .A(g26670) );
  INV_X1 NOT_10705( .ZN(g26896), .A(II35095) );
  INV_X1 NOT_10706( .ZN(II35099), .A(g26672) );
  INV_X1 NOT_10707( .ZN(g26900), .A(II35099) );
  INV_X1 NOT_10708( .ZN(II35106), .A(g26675) );
  INV_X1 NOT_10709( .ZN(g26909), .A(II35106) );
  INV_X1 NOT_10710( .ZN(II35109), .A(g26676) );
  INV_X1 NOT_10711( .ZN(g26910), .A(II35109) );
  INV_X1 NOT_10712( .ZN(II35116), .A(g26025) );
  INV_X1 NOT_10713( .ZN(g26921), .A(II35116) );
  INV_X1 NOT_10714( .ZN(g26922), .A(g26283) );
  INV_X1 NOT_10715( .ZN(g26935), .A(g26327) );
  INV_X1 NOT_10716( .ZN(g26944), .A(g26374) );
  INV_X1 NOT_10717( .ZN(g26950), .A(g26417) );
  INV_X1 NOT_10718( .ZN(II35136), .A(g26660) );
  INV_X1 NOT_10719( .ZN(g26953), .A(II35136) );
  INV_X1 NOT_10720( .ZN(g26954), .A(g26549) );
  INV_X1 NOT_10721( .ZN(II35141), .A(g26666) );
  INV_X1 NOT_10722( .ZN(g26956), .A(II35141) );
  INV_X1 NOT_10723( .ZN(g26957), .A(g26577) );
  INV_X1 NOT_10724( .ZN(II35146), .A(g26671) );
  INV_X1 NOT_10725( .ZN(g26959), .A(II35146) );
  INV_X1 NOT_10726( .ZN(g26960), .A(g26597) );
  INV_X1 NOT_10727( .ZN(II35153), .A(g26677) );
  INV_X1 NOT_10728( .ZN(g26964), .A(II35153) );
  INV_X1 NOT_10729( .ZN(II35172), .A(g26272) );
  INV_X1 NOT_10730( .ZN(g26983), .A(II35172) );
  INV_X1 NOT_10731( .ZN(g26987), .A(g26056) );
  INV_X1 NOT_10732( .ZN(g27010), .A(g26063) );
  INV_X1 NOT_10733( .ZN(g27036), .A(g26070) );
  INV_X1 NOT_10734( .ZN(g27064), .A(g26076) );
  INV_X1 NOT_10735( .ZN(II35254), .A(g26048) );
  INV_X1 NOT_10736( .ZN(g27075), .A(II35254) );
  INV_X1 NOT_10737( .ZN(II35283), .A(g26031) );
  INV_X1 NOT_10738( .ZN(g27102), .A(II35283) );
  INV_X1 NOT_10739( .ZN(II35297), .A(g26199) );
  INV_X1 NOT_10740( .ZN(g27114), .A(II35297) );
  INV_X1 NOT_10741( .ZN(II35301), .A(g26037) );
  INV_X1 NOT_10742( .ZN(g27116), .A(II35301) );
  INV_X1 NOT_10743( .ZN(II35313), .A(g26534) );
  INV_X1 NOT_10744( .ZN(g27126), .A(II35313) );
  INV_X1 NOT_10745( .ZN(II35319), .A(g26183) );
  INV_X1 NOT_10746( .ZN(g27132), .A(II35319) );
  INV_X1 NOT_10747( .ZN(g27133), .A(g26105) );
  INV_X1 NOT_10748( .ZN(g27134), .A(g26175) );
  INV_X1 NOT_10749( .ZN(g27135), .A(g26178) );
  INV_X1 NOT_10750( .ZN(g27136), .A(g26196) );
  INV_X1 NOT_10751( .ZN(g27137), .A(g26202) );
  INV_X1 NOT_10752( .ZN(g27138), .A(g26223) );
  INV_X1 NOT_10753( .ZN(g27139), .A(g26226) );
  INV_X1 NOT_10754( .ZN(g27140), .A(g26136) );
  INV_X1 NOT_10755( .ZN(g27141), .A(g26251) );
  INV_X1 NOT_10756( .ZN(g27142), .A(g26254) );
  INV_X1 NOT_10757( .ZN(g27143), .A(g26150) );
  INV_X4 NOT_10758( .ZN(II35334), .A(g26106) );
  INV_X1 NOT_10759( .ZN(g27145), .A(II35334) );
  INV_X1 NOT_10760( .ZN(g27146), .A(g26358) );
  INV_X1 NOT_10761( .ZN(g27148), .A(g26393) );
  INV_X1 NOT_10762( .ZN(II35341), .A(g26120) );
  INV_X1 NOT_10763( .ZN(g27150), .A(II35341) );
  INV_X1 NOT_10764( .ZN(g27151), .A(g26401) );
  INV_X1 NOT_10765( .ZN(g27153), .A(g26429) );
  INV_X1 NOT_10766( .ZN(II35347), .A(g26265) );
  INV_X1 NOT_10767( .ZN(g27154), .A(II35347) );
  INV_X1 NOT_10768( .ZN(g27155), .A(g26434) );
  INV_X1 NOT_10769( .ZN(II35351), .A(g26272) );
  INV_X1 NOT_10770( .ZN(g27156), .A(II35351) );
  INV_X1 NOT_10771( .ZN(II35355), .A(g26130) );
  INV_X1 NOT_10772( .ZN(g27158), .A(II35355) );
  INV_X1 NOT_10773( .ZN(g27159), .A(g26442) );
  INV_X1 NOT_10774( .ZN(II35360), .A(g26295) );
  INV_X1 NOT_10775( .ZN(g27161), .A(II35360) );
  INV_X1 NOT_10776( .ZN(g27162), .A(g26461) );
  INV_X1 NOT_10777( .ZN(II35364), .A(g26304) );
  INV_X1 NOT_10778( .ZN(g27163), .A(II35364) );
  INV_X1 NOT_10779( .ZN(g27164), .A(g26466) );
  INV_X1 NOT_10780( .ZN(II35369), .A(g26144) );
  INV_X1 NOT_10781( .ZN(g27166), .A(II35369) );
  INV_X1 NOT_10782( .ZN(g27167), .A(g26474) );
  INV_X1 NOT_10783( .ZN(II35373), .A(g26189) );
  INV_X1 NOT_10784( .ZN(g27168), .A(II35373) );
  INV_X1 NOT_10785( .ZN(II35376), .A(g26336) );
  INV_X1 NOT_10786( .ZN(g27171), .A(II35376) );
  INV_X1 NOT_10787( .ZN(g27172), .A(g26485) );
  INV_X1 NOT_10788( .ZN(g27173), .A(g26490) );
  INV_X1 NOT_10789( .ZN(II35383), .A(g26160) );
  INV_X1 NOT_10790( .ZN(g27176), .A(II35383) );
  INV_X1 NOT_10791( .ZN(g27177), .A(g26501) );
  INV_X1 NOT_10792( .ZN(II35389), .A(g26168) );
  INV_X1 NOT_10793( .ZN(g27180), .A(II35389) );
  INV_X1 NOT_10794( .ZN(II35394), .A(g26183) );
  INV_X1 NOT_10795( .ZN(g27183), .A(II35394) );
  INV_X1 NOT_10796( .ZN(II35399), .A(g26199) );
  INV_X1 NOT_10797( .ZN(g27186), .A(II35399) );
  INV_X1 NOT_10798( .ZN(II35404), .A(g26864) );
  INV_X1 NOT_10799( .ZN(g27189), .A(II35404) );
  INV_X1 NOT_10800( .ZN(II35407), .A(g27145) );
  INV_X1 NOT_10801( .ZN(g27190), .A(II35407) );
  INV_X1 NOT_10802( .ZN(II35410), .A(g26872) );
  INV_X1 NOT_10803( .ZN(g27191), .A(II35410) );
  INV_X1 NOT_10804( .ZN(II35413), .A(g26876) );
  INV_X1 NOT_10805( .ZN(g27192), .A(II35413) );
  INV_X1 NOT_10806( .ZN(II35416), .A(g26884) );
  INV_X1 NOT_10807( .ZN(g27193), .A(II35416) );
  INV_X1 NOT_10808( .ZN(II35419), .A(g26828) );
  INV_X1 NOT_10809( .ZN(g27194), .A(II35419) );
  INV_X1 NOT_10810( .ZN(II35422), .A(g26830) );
  INV_X4 NOT_10811( .ZN(g27195), .A(II35422) );
  INV_X1 NOT_10812( .ZN(II35425), .A(g26832) );
  INV_X1 NOT_10813( .ZN(g27196), .A(II35425) );
  INV_X1 NOT_10814( .ZN(II35428), .A(g26953) );
  INV_X1 NOT_10815( .ZN(g27197), .A(II35428) );
  INV_X1 NOT_10816( .ZN(II35431), .A(g26868) );
  INV_X1 NOT_10817( .ZN(g27198), .A(II35431) );
  INV_X1 NOT_10818( .ZN(II35434), .A(g27150) );
  INV_X1 NOT_10819( .ZN(g27199), .A(II35434) );
  INV_X1 NOT_10820( .ZN(II35437), .A(g27183) );
  INV_X1 NOT_10821( .ZN(g27200), .A(II35437) );
  INV_X1 NOT_10822( .ZN(II35440), .A(g27186) );
  INV_X1 NOT_10823( .ZN(g27201), .A(II35440) );
  INV_X1 NOT_10824( .ZN(II35443), .A(g26757) );
  INV_X1 NOT_10825( .ZN(g27202), .A(II35443) );
  INV_X1 NOT_10826( .ZN(II35446), .A(g26762) );
  INV_X1 NOT_10827( .ZN(g27203), .A(II35446) );
  INV_X1 NOT_10828( .ZN(II35449), .A(g27154) );
  INV_X1 NOT_10829( .ZN(g27204), .A(II35449) );
  INV_X1 NOT_10830( .ZN(II35452), .A(g27161) );
  INV_X1 NOT_10831( .ZN(g27205), .A(II35452) );
  INV_X1 NOT_10832( .ZN(II35455), .A(g26881) );
  INV_X1 NOT_10833( .ZN(g27206), .A(II35455) );
  INV_X1 NOT_10834( .ZN(II35458), .A(g26886) );
  INV_X1 NOT_10835( .ZN(g27207), .A(II35458) );
  INV_X1 NOT_10836( .ZN(II35461), .A(g26895) );
  INV_X1 NOT_10837( .ZN(g27208), .A(II35461) );
  INV_X1 NOT_10838( .ZN(II35464), .A(g26831) );
  INV_X1 NOT_10839( .ZN(g27209), .A(II35464) );
  INV_X1 NOT_10840( .ZN(II35467), .A(g26834) );
  INV_X1 NOT_10841( .ZN(g27210), .A(II35467) );
  INV_X1 NOT_10842( .ZN(II35470), .A(g26840) );
  INV_X1 NOT_10843( .ZN(g27211), .A(II35470) );
  INV_X1 NOT_10844( .ZN(II35473), .A(g27156) );
  INV_X1 NOT_10845( .ZN(g27212), .A(II35473) );
  INV_X1 NOT_10846( .ZN(II35476), .A(g27163) );
  INV_X1 NOT_10847( .ZN(g27213), .A(II35476) );
  INV_X1 NOT_10848( .ZN(II35479), .A(g27171) );
  INV_X1 NOT_10849( .ZN(g27214), .A(II35479) );
  INV_X1 NOT_10850( .ZN(II35482), .A(g27176) );
  INV_X1 NOT_10851( .ZN(g27215), .A(II35482) );
  INV_X1 NOT_10852( .ZN(II35485), .A(g27180) );
  INV_X1 NOT_10853( .ZN(g27216), .A(II35485) );
  INV_X1 NOT_10854( .ZN(II35488), .A(g26819) );
  INV_X1 NOT_10855( .ZN(g27217), .A(II35488) );
  INV_X1 NOT_10856( .ZN(II35491), .A(g26956) );
  INV_X1 NOT_10857( .ZN(g27218), .A(II35491) );
  INV_X1 NOT_10858( .ZN(II35494), .A(g26875) );
  INV_X1 NOT_10859( .ZN(g27219), .A(II35494) );
  INV_X1 NOT_10860( .ZN(II35497), .A(g27158) );
  INV_X1 NOT_10861( .ZN(g27220), .A(II35497) );
  INV_X1 NOT_10862( .ZN(II35500), .A(g26890) );
  INV_X1 NOT_10863( .ZN(g27221), .A(II35500) );
  INV_X1 NOT_10864( .ZN(II35503), .A(g26896) );
  INV_X1 NOT_10865( .ZN(g27222), .A(II35503) );
  INV_X1 NOT_10866( .ZN(II35506), .A(g26909) );
  INV_X1 NOT_10867( .ZN(g27223), .A(II35506) );
  INV_X1 NOT_10868( .ZN(II35509), .A(g26836) );
  INV_X1 NOT_10869( .ZN(g27224), .A(II35509) );
  INV_X1 NOT_10870( .ZN(II35512), .A(g26843) );
  INV_X1 NOT_10871( .ZN(g27225), .A(II35512) );
  INV_X4 NOT_10872( .ZN(II35515), .A(g26850) );
  INV_X1 NOT_10873( .ZN(g27226), .A(II35515) );
  INV_X1 NOT_10874( .ZN(II35518), .A(g26959) );
  INV_X1 NOT_10875( .ZN(g27227), .A(II35518) );
  INV_X1 NOT_10876( .ZN(II35521), .A(g26883) );
  INV_X1 NOT_10877( .ZN(g27228), .A(II35521) );
  INV_X1 NOT_10878( .ZN(II35524), .A(g27166) );
  INV_X1 NOT_10879( .ZN(g27229), .A(II35524) );
  INV_X1 NOT_10880( .ZN(II35527), .A(g26900) );
  INV_X1 NOT_10881( .ZN(g27230), .A(II35527) );
  INV_X1 NOT_10882( .ZN(II35530), .A(g26910) );
  INV_X1 NOT_10883( .ZN(g27231), .A(II35530) );
  INV_X1 NOT_10884( .ZN(II35533), .A(g26921) );
  INV_X1 NOT_10885( .ZN(g27232), .A(II35533) );
  INV_X1 NOT_10886( .ZN(II35536), .A(g26844) );
  INV_X1 NOT_10887( .ZN(g27233), .A(II35536) );
  INV_X1 NOT_10888( .ZN(II35539), .A(g26852) );
  INV_X1 NOT_10889( .ZN(g27234), .A(II35539) );
  INV_X1 NOT_10890( .ZN(II35542), .A(g26858) );
  INV_X1 NOT_10891( .ZN(g27235), .A(II35542) );
  INV_X1 NOT_10892( .ZN(II35545), .A(g26964) );
  INV_X1 NOT_10893( .ZN(g27236), .A(II35545) );
  INV_X1 NOT_10894( .ZN(II35548), .A(g27116) );
  INV_X1 NOT_10895( .ZN(g27237), .A(II35548) );
  INV_X1 NOT_10896( .ZN(II35551), .A(g27075) );
  INV_X1 NOT_10897( .ZN(g27238), .A(II35551) );
  INV_X1 NOT_10898( .ZN(II35554), .A(g27102) );
  INV_X1 NOT_10899( .ZN(g27239), .A(II35554) );
  INV_X1 NOT_10900( .ZN(g27349), .A(g27126) );
  INV_X4 NOT_10901( .ZN(II35667), .A(g27120) );
  INV_X1 NOT_10902( .ZN(g27353), .A(II35667) );
  INV_X1 NOT_10903( .ZN(II35673), .A(g27123) );
  INV_X1 NOT_10904( .ZN(g27357), .A(II35673) );
  INV_X1 NOT_10905( .ZN(II35678), .A(g27129) );
  INV_X1 NOT_10906( .ZN(g27360), .A(II35678) );
  INV_X1 NOT_10907( .ZN(II35681), .A(g26869) );
  INV_X1 NOT_10908( .ZN(g27361), .A(II35681) );
  INV_X1 NOT_10909( .ZN(II35686), .A(g27131) );
  INV_X1 NOT_10910( .ZN(g27366), .A(II35686) );
  INV_X1 NOT_10911( .ZN(II35689), .A(g26878) );
  INV_X1 NOT_10912( .ZN(g27367), .A(II35689) );
  INV_X1 NOT_10913( .ZN(II35695), .A(g26887) );
  INV_X1 NOT_10914( .ZN(g27373), .A(II35695) );
  INV_X1 NOT_10915( .ZN(II35698), .A(g26897) );
  INV_X1 NOT_10916( .ZN(g27376), .A(II35698) );
  INV_X1 NOT_10917( .ZN(II35708), .A(g26974) );
  INV_X1 NOT_10918( .ZN(g27380), .A(II35708) );
  INV_X1 NOT_10919( .ZN(II35711), .A(g26974) );
  INV_X1 NOT_10920( .ZN(g27381), .A(II35711) );
  INV_X1 NOT_10921( .ZN(g27383), .A(g27133) );
  INV_X1 NOT_10922( .ZN(g27384), .A(g27140) );
  INV_X1 NOT_10923( .ZN(II35723), .A(g27168) );
  INV_X1 NOT_10924( .ZN(g27385), .A(II35723) );
  INV_X1 NOT_10925( .ZN(g27386), .A(g27143) );
  INV_X1 NOT_10926( .ZN(II35727), .A(g26902) );
  INV_X1 NOT_10927( .ZN(g27387), .A(II35727) );
  INV_X1 NOT_10928( .ZN(II35731), .A(g26892) );
  INV_X1 NOT_10929( .ZN(g27391), .A(II35731) );
  INV_X1 NOT_10930( .ZN(II35737), .A(g26915) );
  INV_X1 NOT_10931( .ZN(g27397), .A(II35737) );
  INV_X1 NOT_10932( .ZN(II35741), .A(g27118) );
  INV_X1 NOT_10933( .ZN(g27401), .A(II35741) );
  INV_X1 NOT_10934( .ZN(II35744), .A(g26906) );
  INV_X1 NOT_10935( .ZN(g27404), .A(II35744) );
  INV_X1 NOT_10936( .ZN(II35750), .A(g26928) );
  INV_X1 NOT_10937( .ZN(g27410), .A(II35750) );
  INV_X1 NOT_10938( .ZN(II35756), .A(g27117) );
  INV_X1 NOT_10939( .ZN(g27416), .A(II35756) );
  INV_X1 NOT_10940( .ZN(II35759), .A(g27121) );
  INV_X1 NOT_10941( .ZN(g27419), .A(II35759) );
  INV_X1 NOT_10942( .ZN(II35762), .A(g26918) );
  INV_X1 NOT_10943( .ZN(g27422), .A(II35762) );
  INV_X1 NOT_10944( .ZN(II35768), .A(g26941) );
  INV_X1 NOT_10945( .ZN(g27428), .A(II35768) );
  INV_X1 NOT_10946( .ZN(II35772), .A(g26772) );
  INV_X1 NOT_10947( .ZN(g27432), .A(II35772) );
  INV_X1 NOT_10948( .ZN(II35777), .A(g27119) );
  INV_X1 NOT_10949( .ZN(g27437), .A(II35777) );
  INV_X1 NOT_10950( .ZN(II35780), .A(g27124) );
  INV_X1 NOT_10951( .ZN(g27440), .A(II35780) );
  INV_X1 NOT_10952( .ZN(II35783), .A(g26931) );
  INV_X1 NOT_10953( .ZN(g27443), .A(II35783) );
  INV_X1 NOT_10954( .ZN(g27449), .A(g26837) );
  INV_X1 NOT_10955( .ZN(II35791), .A(g26779) );
  INV_X1 NOT_10956( .ZN(g27451), .A(II35791) );
  INV_X1 NOT_10957( .ZN(II35796), .A(g27122) );
  INV_X1 NOT_10958( .ZN(g27456), .A(II35796) );
  INV_X1 NOT_10959( .ZN(II35799), .A(g27130) );
  INV_X1 NOT_10960( .ZN(g27459), .A(II35799) );
  INV_X1 NOT_10961( .ZN(II35803), .A(g26803) );
  INV_X1 NOT_10962( .ZN(g27463), .A(II35803) );
  INV_X1 NOT_10963( .ZN(g27465), .A(g26846) );
  INV_X1 NOT_10964( .ZN(II35809), .A(g26785) );
  INV_X1 NOT_10965( .ZN(g27467), .A(II35809) );
  INV_X1 NOT_10966( .ZN(II35814), .A(g27125) );
  INV_X1 NOT_10967( .ZN(g27472), .A(II35814) );
  INV_X1 NOT_10968( .ZN(II35817), .A(g26922) );
  INV_X1 NOT_10969( .ZN(g27475), .A(II35817) );
  INV_X1 NOT_10970( .ZN(II35821), .A(g26804) );
  INV_X1 NOT_10971( .ZN(g27479), .A(II35821) );
  INV_X1 NOT_10972( .ZN(II35824), .A(g26805) );
  INV_X1 NOT_10973( .ZN(g27480), .A(II35824) );
  INV_X1 NOT_10974( .ZN(II35829), .A(g26806) );
  INV_X1 NOT_10975( .ZN(g27483), .A(II35829) );
  INV_X1 NOT_10976( .ZN(g27484), .A(g26855) );
  INV_X1 NOT_10977( .ZN(II35834), .A(g26792) );
  INV_X1 NOT_10978( .ZN(g27486), .A(II35834) );
  INV_X1 NOT_10979( .ZN(II35837), .A(g26911) );
  INV_X1 NOT_10980( .ZN(g27489), .A(II35837) );
  INV_X1 NOT_10981( .ZN(II35841), .A(g26807) );
  INV_X1 NOT_10982( .ZN(g27493), .A(II35841) );
  INV_X1 NOT_10983( .ZN(II35844), .A(g26808) );
  INV_X1 NOT_10984( .ZN(g27494), .A(II35844) );
  INV_X1 NOT_10985( .ZN(II35849), .A(g26776) );
  INV_X1 NOT_10986( .ZN(g27497), .A(II35849) );
  INV_X1 NOT_10987( .ZN(II35852), .A(g26935) );
  INV_X1 NOT_10988( .ZN(g27498), .A(II35852) );
  INV_X1 NOT_10989( .ZN(II35856), .A(g26809) );
  INV_X1 NOT_10990( .ZN(g27502), .A(II35856) );
  INV_X1 NOT_10991( .ZN(II35859), .A(g26810) );
  INV_X1 NOT_10992( .ZN(g27503), .A(II35859) );
  INV_X1 NOT_10993( .ZN(II35863), .A(g26811) );
  INV_X1 NOT_10994( .ZN(g27505), .A(II35863) );
  INV_X1 NOT_10995( .ZN(g27506), .A(g26861) );
  INV_X1 NOT_10996( .ZN(II35868), .A(g26812) );
  INV_X1 NOT_10997( .ZN(g27508), .A(II35868) );
  INV_X1 NOT_10998( .ZN(II35872), .A(g26925) );
  INV_X1 NOT_10999( .ZN(g27510), .A(II35872) );
  INV_X1 NOT_11000( .ZN(II35876), .A(g26813) );
  INV_X1 NOT_11001( .ZN(g27514), .A(II35876) );
  INV_X1 NOT_11002( .ZN(II35879), .A(g26814) );
  INV_X1 NOT_11003( .ZN(g27515), .A(II35879) );
  INV_X1 NOT_11004( .ZN(II35883), .A(g26781) );
  INV_X1 NOT_11005( .ZN(g27517), .A(II35883) );
  INV_X1 NOT_11006( .ZN(II35886), .A(g26944) );
  INV_X1 NOT_11007( .ZN(g27518), .A(II35886) );
  INV_X1 NOT_11008( .ZN(II35890), .A(g26815) );
  INV_X1 NOT_11009( .ZN(g27522), .A(II35890) );
  INV_X1 NOT_11010( .ZN(II35893), .A(g26816) );
  INV_X1 NOT_11011( .ZN(g27523), .A(II35893) );
  INV_X1 NOT_11012( .ZN(II35897), .A(g26817) );
  INV_X1 NOT_11013( .ZN(g27525), .A(II35897) );
  INV_X1 NOT_11014( .ZN(II35900), .A(g26786) );
  INV_X1 NOT_11015( .ZN(g27526), .A(II35900) );
  INV_X1 NOT_11016( .ZN(II35915), .A(g26818) );
  INV_X1 NOT_11017( .ZN(g27533), .A(II35915) );
  INV_X1 NOT_11018( .ZN(II35919), .A(g26938) );
  INV_X1 NOT_11019( .ZN(g27535), .A(II35919) );
  INV_X1 NOT_11020( .ZN(II35923), .A(g26820) );
  INV_X1 NOT_11021( .ZN(g27539), .A(II35923) );
  INV_X1 NOT_11022( .ZN(II35926), .A(g26821) );
  INV_X1 NOT_11023( .ZN(g27540), .A(II35926) );
  INV_X1 NOT_11024( .ZN(II35930), .A(g26789) );
  INV_X1 NOT_11025( .ZN(g27542), .A(II35930) );
  INV_X1 NOT_11026( .ZN(II35933), .A(g26950) );
  INV_X1 NOT_11027( .ZN(g27543), .A(II35933) );
  INV_X1 NOT_11028( .ZN(II35937), .A(g26822) );
  INV_X1 NOT_11029( .ZN(g27547), .A(II35937) );
  INV_X1 NOT_11030( .ZN(II35940), .A(g26823) );
  INV_X1 NOT_11031( .ZN(g27548), .A(II35940) );
  INV_X1 NOT_11032( .ZN(II35953), .A(g26824) );
  INV_X1 NOT_11033( .ZN(g27553), .A(II35953) );
  INV_X1 NOT_11034( .ZN(II35957), .A(g26947) );
  INV_X1 NOT_11035( .ZN(g27555), .A(II35957) );
  INV_X1 NOT_11036( .ZN(II35961), .A(g26825) );
  INV_X1 NOT_11037( .ZN(g27559), .A(II35961) );
  INV_X1 NOT_11038( .ZN(II35964), .A(g26826) );
  INV_X1 NOT_11039( .ZN(g27560), .A(II35964) );
  INV_X1 NOT_11040( .ZN(II35968), .A(g26795) );
  INV_X1 NOT_11041( .ZN(g27562), .A(II35968) );
  INV_X1 NOT_11042( .ZN(II35983), .A(g26827) );
  INV_X1 NOT_11043( .ZN(g27569), .A(II35983) );
  INV_X1 NOT_11044( .ZN(II36008), .A(g26798) );
  INV_X1 NOT_11045( .ZN(g27586), .A(II36008) );
  INV_X1 NOT_11046( .ZN(g27589), .A(g27168) );
  INV_X1 NOT_11047( .ZN(g27590), .A(g27144) );
  INV_X1 NOT_11048( .ZN(g27595), .A(g27149) );
  INV_X1 NOT_11049( .ZN(g27599), .A(g27147) );
  INV_X1 NOT_11050( .ZN(g27604), .A(g27157) );
  INV_X1 NOT_11051( .ZN(g27608), .A(g27152) );
  INV_X1 NOT_11052( .ZN(g27613), .A(g27165) );
  INV_X1 NOT_11053( .ZN(g27617), .A(g27160) );
  INV_X1 NOT_11054( .ZN(g27622), .A(g27174) );
  INV_X1 NOT_11055( .ZN(II36032), .A(g27113) );
  INV_X1 NOT_11056( .ZN(g27632), .A(II36032) );
  INV_X1 NOT_11057( .ZN(II36042), .A(g26960) );
  INV_X1 NOT_11058( .ZN(g27662), .A(II36042) );
  INV_X1 NOT_11059( .ZN(II36046), .A(g26957) );
  INV_X1 NOT_11060( .ZN(g27667), .A(II36046) );
  INV_X1 NOT_11061( .ZN(II36052), .A(g26954) );
  INV_X1 NOT_11062( .ZN(g27674), .A(II36052) );
  INV_X1 NOT_11063( .ZN(II36060), .A(g27353) );
  INV_X1 NOT_11064( .ZN(g27683), .A(II36060) );
  INV_X1 NOT_11065( .ZN(II36063), .A(g27463) );
  INV_X1 NOT_11066( .ZN(g27684), .A(II36063) );
  INV_X1 NOT_11067( .ZN(II36066), .A(g27479) );
  INV_X1 NOT_11068( .ZN(g27685), .A(II36066) );
  INV_X1 NOT_11069( .ZN(II36069), .A(g27493) );
  INV_X1 NOT_11070( .ZN(g27686), .A(II36069) );
  INV_X1 NOT_11071( .ZN(II36072), .A(g27480) );
  INV_X1 NOT_11072( .ZN(g27687), .A(II36072) );
  INV_X1 NOT_11073( .ZN(II36075), .A(g27494) );
  INV_X1 NOT_11074( .ZN(g27688), .A(II36075) );
  INV_X1 NOT_11075( .ZN(II36078), .A(g27508) );
  INV_X1 NOT_11076( .ZN(g27689), .A(II36078) );
  INV_X1 NOT_11077( .ZN(II36081), .A(g27497) );
  INV_X1 NOT_11078( .ZN(g27690), .A(II36081) );
  INV_X1 NOT_11079( .ZN(II36084), .A(g27357) );
  INV_X1 NOT_11080( .ZN(g27691), .A(II36084) );
  INV_X1 NOT_11081( .ZN(II36087), .A(g27483) );
  INV_X1 NOT_11082( .ZN(g27692), .A(II36087) );
  INV_X1 NOT_11083( .ZN(II36090), .A(g27502) );
  INV_X1 NOT_11084( .ZN(g27693), .A(II36090) );
  INV_X1 NOT_11085( .ZN(II36093), .A(g27514) );
  INV_X1 NOT_11086( .ZN(g27694), .A(II36093) );
  INV_X1 NOT_11087( .ZN(II36096), .A(g27503) );
  INV_X1 NOT_11088( .ZN(g27695), .A(II36096) );
  INV_X1 NOT_11089( .ZN(II36099), .A(g27515) );
  INV_X1 NOT_11090( .ZN(g27696), .A(II36099) );
  INV_X4 NOT_11091( .ZN(II36102), .A(g27533) );
  INV_X4 NOT_11092( .ZN(g27697), .A(II36102) );
  INV_X4 NOT_11093( .ZN(II36105), .A(g27517) );
  INV_X4 NOT_11094( .ZN(g27698), .A(II36105) );
  INV_X4 NOT_11095( .ZN(II36108), .A(g27360) );
  INV_X4 NOT_11096( .ZN(g27699), .A(II36108) );
  INV_X4 NOT_11097( .ZN(II36111), .A(g27505) );
  INV_X1 NOT_11098( .ZN(g27700), .A(II36111) );
  INV_X1 NOT_11099( .ZN(II36114), .A(g27522) );
  INV_X1 NOT_11100( .ZN(g27701), .A(II36114) );
  INV_X1 NOT_11101( .ZN(II36117), .A(g27539) );
  INV_X1 NOT_11102( .ZN(g27702), .A(II36117) );
  INV_X1 NOT_11103( .ZN(II36120), .A(g27523) );
  INV_X1 NOT_11104( .ZN(g27703), .A(II36120) );
  INV_X1 NOT_11105( .ZN(II36123), .A(g27540) );
  INV_X1 NOT_11106( .ZN(g27704), .A(II36123) );
  INV_X1 NOT_11107( .ZN(II36126), .A(g27553) );
  INV_X1 NOT_11108( .ZN(g27705), .A(II36126) );
  INV_X1 NOT_11109( .ZN(II36129), .A(g27542) );
  INV_X1 NOT_11110( .ZN(g27706), .A(II36129) );
  INV_X1 NOT_11111( .ZN(II36132), .A(g27366) );
  INV_X1 NOT_11112( .ZN(g27707), .A(II36132) );
  INV_X1 NOT_11113( .ZN(II36135), .A(g27525) );
  INV_X1 NOT_11114( .ZN(g27708), .A(II36135) );
  INV_X1 NOT_11115( .ZN(II36138), .A(g27547) );
  INV_X1 NOT_11116( .ZN(g27709), .A(II36138) );
  INV_X1 NOT_11117( .ZN(II36141), .A(g27559) );
  INV_X1 NOT_11118( .ZN(g27710), .A(II36141) );
  INV_X1 NOT_11119( .ZN(II36144), .A(g27548) );
  INV_X1 NOT_11120( .ZN(g27711), .A(II36144) );
  INV_X1 NOT_11121( .ZN(II36147), .A(g27560) );
  INV_X1 NOT_11122( .ZN(g27712), .A(II36147) );
  INV_X1 NOT_11123( .ZN(II36150), .A(g27569) );
  INV_X1 NOT_11124( .ZN(g27713), .A(II36150) );
  INV_X1 NOT_11125( .ZN(II36153), .A(g27562) );
  INV_X1 NOT_11126( .ZN(g27714), .A(II36153) );
  INV_X1 NOT_11127( .ZN(II36156), .A(g27586) );
  INV_X1 NOT_11128( .ZN(g27715), .A(II36156) );
  INV_X1 NOT_11129( .ZN(II36159), .A(g27526) );
  INV_X1 NOT_11130( .ZN(g27716), .A(II36159) );
  INV_X1 NOT_11131( .ZN(II36162), .A(g27385) );
  INV_X1 NOT_11132( .ZN(g27717), .A(II36162) );
  INV_X1 NOT_11133( .ZN(g27748), .A(g27632) );
  INV_X1 NOT_11134( .ZN(II36213), .A(g27571) );
  INV_X1 NOT_11135( .ZN(g27776), .A(II36213) );
  INV_X1 NOT_11136( .ZN(II36217), .A(g27580) );
  INV_X1 NOT_11137( .ZN(g27780), .A(II36217) );
  INV_X1 NOT_11138( .ZN(II36221), .A(g27662) );
  INV_X1 NOT_11139( .ZN(g27784), .A(II36221) );
  INV_X1 NOT_11140( .ZN(II36224), .A(g27589) );
  INV_X1 NOT_11141( .ZN(g27785), .A(II36224) );
  INV_X1 NOT_11142( .ZN(II36227), .A(g27594) );
  INV_X1 NOT_11143( .ZN(g27786), .A(II36227) );
  INV_X1 NOT_11144( .ZN(II36230), .A(g27583) );
  INV_X1 NOT_11145( .ZN(g27787), .A(II36230) );
  INV_X1 NOT_11146( .ZN(II36234), .A(g27667) );
  INV_X1 NOT_11147( .ZN(g27791), .A(II36234) );
  INV_X1 NOT_11148( .ZN(II36237), .A(g27662) );
  INV_X1 NOT_11149( .ZN(g27792), .A(II36237) );
  INV_X1 NOT_11150( .ZN(II36240), .A(g27603) );
  INV_X1 NOT_11151( .ZN(g27793), .A(II36240) );
  INV_X1 NOT_11152( .ZN(II36243), .A(g27587) );
  INV_X1 NOT_11153( .ZN(g27794), .A(II36243) );
  INV_X1 NOT_11154( .ZN(II36246), .A(g27674) );
  INV_X1 NOT_11155( .ZN(g27797), .A(II36246) );
  INV_X1 NOT_11156( .ZN(II36250), .A(g27612) );
  INV_X1 NOT_11157( .ZN(g27799), .A(II36250) );
  INV_X1 NOT_11158( .ZN(II36253), .A(g27674) );
  INV_X1 NOT_11159( .ZN(g27800), .A(II36253) );
  INV_X1 NOT_11160( .ZN(II36264), .A(g27621) );
  INV_X1 NOT_11161( .ZN(g27805), .A(II36264) );
  INV_X1 NOT_11162( .ZN(II36267), .A(g27395) );
  INV_X1 NOT_11163( .ZN(g27806), .A(II36267) );
  INV_X1 NOT_11164( .ZN(II36280), .A(g27390) );
  INV_X1 NOT_11165( .ZN(g27817), .A(II36280) );
  INV_X1 NOT_11166( .ZN(II36283), .A(g27408) );
  INV_X1 NOT_11167( .ZN(g27820), .A(II36283) );
  INV_X1 NOT_11168( .ZN(II36296), .A(g27626) );
  INV_X1 NOT_11169( .ZN(g27831), .A(II36296) );
  INV_X1 NOT_11170( .ZN(II36307), .A(g27400) );
  INV_X1 NOT_11171( .ZN(g27839), .A(II36307) );
  INV_X1 NOT_11172( .ZN(II36311), .A(g27426) );
  INV_X1 NOT_11173( .ZN(g27843), .A(II36311) );
  INV_X1 NOT_11174( .ZN(II36321), .A(g27627) );
  INV_X1 NOT_11175( .ZN(g27847), .A(II36321) );
  INV_X1 NOT_11176( .ZN(II36327), .A(g27413) );
  INV_X1 NOT_11177( .ZN(g27858), .A(II36327) );
  INV_X1 NOT_11178( .ZN(II36330), .A(g27447) );
  INV_X1 NOT_11179( .ZN(g27861), .A(II36330) );
  INV_X1 NOT_11180( .ZN(II36337), .A(g27628) );
  INV_X1 NOT_11181( .ZN(g27872), .A(II36337) );
  INV_X1 NOT_11182( .ZN(II36341), .A(g27431) );
  INV_X1 NOT_11183( .ZN(g27879), .A(II36341) );
  INV_X1 NOT_11184( .ZN(II36347), .A(g27630) );
  INV_X1 NOT_11185( .ZN(g27889), .A(II36347) );
  INV_X1 NOT_11186( .ZN(II36354), .A(g27662) );
  INV_X1 NOT_11187( .ZN(g27903), .A(II36354) );
  INV_X1 NOT_11188( .ZN(II36358), .A(g27672) );
  INV_X1 NOT_11189( .ZN(g27905), .A(II36358) );
  INV_X1 NOT_11190( .ZN(II36362), .A(g27667) );
  INV_X1 NOT_11191( .ZN(g27907), .A(II36362) );
  INV_X1 NOT_11192( .ZN(II36367), .A(g27678) );
  INV_X1 NOT_11193( .ZN(g27910), .A(II36367) );
  INV_X1 NOT_11194( .ZN(II36371), .A(g27674) );
  INV_X1 NOT_11195( .ZN(g27912), .A(II36371) );
  INV_X1 NOT_11196( .ZN(II36379), .A(g27682) );
  INV_X1 NOT_11197( .ZN(g27918), .A(II36379) );
  INV_X1 NOT_11198( .ZN(II36382), .A(g27563) );
  INV_X1 NOT_11199( .ZN(g27919), .A(II36382) );
  INV_X1 NOT_11200( .ZN(II36390), .A(g27243) );
  INV_X1 NOT_11201( .ZN(g27927), .A(II36390) );
  INV_X1 NOT_11202( .ZN(II36393), .A(g27572) );
  INV_X1 NOT_11203( .ZN(g27928), .A(II36393) );
  INV_X1 NOT_11204( .ZN(II36397), .A(g27574) );
  INV_X1 NOT_11205( .ZN(g27932), .A(II36397) );
  INV_X1 NOT_11206( .ZN(II36404), .A(g27450) );
  INV_X1 NOT_11207( .ZN(g27939), .A(II36404) );
  INV_X1 NOT_11208( .ZN(II36407), .A(g27581) );
  INV_X1 NOT_11209( .ZN(g27942), .A(II36407) );
  INV_X1 NOT_11210( .ZN(II36411), .A(g27582) );
  INV_X1 NOT_11211( .ZN(g27946), .A(II36411) );
  INV_X1 NOT_11212( .ZN(II36417), .A(g27462) );
  INV_X1 NOT_11213( .ZN(g27952), .A(II36417) );
  INV_X1 NOT_11214( .ZN(II36420), .A(g27253) );
  INV_X1 NOT_11215( .ZN(g27955), .A(II36420) );
  INV_X1 NOT_11216( .ZN(II36423), .A(g27466) );
  INV_X1 NOT_11217( .ZN(g27956), .A(II36423) );
  INV_X1 NOT_11218( .ZN(II36426), .A(g27584) );
  INV_X1 NOT_11219( .ZN(g27959), .A(II36426) );
  INV_X1 NOT_11220( .ZN(II36432), .A(g27585) );
  INV_X1 NOT_11221( .ZN(g27965), .A(II36432) );
  INV_X1 NOT_11222( .ZN(g27969), .A(g27361) );
  INV_X1 NOT_11223( .ZN(II36438), .A(g27255) );
  INV_X1 NOT_11224( .ZN(g27971), .A(II36438) );
  INV_X1 NOT_11225( .ZN(II36441), .A(g27256) );
  INV_X1 NOT_11226( .ZN(g27972), .A(II36441) );
  INV_X1 NOT_11227( .ZN(II36444), .A(g27482) );
  INV_X1 NOT_11228( .ZN(g27973), .A(II36444) );
  INV_X1 NOT_11229( .ZN(II36447), .A(g27257) );
  INV_X1 NOT_11230( .ZN(g27976), .A(II36447) );
  INV_X1 NOT_11231( .ZN(II36450), .A(g27485) );
  INV_X1 NOT_11232( .ZN(g27977), .A(II36450) );
  INV_X1 NOT_11233( .ZN(II36454), .A(g27588) );
  INV_X1 NOT_11234( .ZN(g27981), .A(II36454) );
  INV_X1 NOT_11235( .ZN(II36459), .A(g27258) );
  INV_X1 NOT_11236( .ZN(g27986), .A(II36459) );
  INV_X1 NOT_11237( .ZN(II36462), .A(g27259) );
  INV_X1 NOT_11238( .ZN(g27987), .A(II36462) );
  INV_X1 NOT_11239( .ZN(II36465), .A(g27260) );
  INV_X1 NOT_11240( .ZN(g27988), .A(II36465) );
  INV_X1 NOT_11241( .ZN(II36468), .A(g27261) );
  INV_X1 NOT_11242( .ZN(g27989), .A(II36468) );
  INV_X1 NOT_11243( .ZN(g27990), .A(g27367) );
  INV_X1 NOT_11244( .ZN(II36473), .A(g27262) );
  INV_X1 NOT_11245( .ZN(g27992), .A(II36473) );
  INV_X1 NOT_11246( .ZN(II36476), .A(g27263) );
  INV_X1 NOT_11247( .ZN(g27993), .A(II36476) );
  INV_X1 NOT_11248( .ZN(II36479), .A(g27504) );
  INV_X1 NOT_11249( .ZN(g27994), .A(II36479) );
  INV_X1 NOT_11250( .ZN(II36483), .A(g27264) );
  INV_X1 NOT_11251( .ZN(g27998), .A(II36483) );
  INV_X1 NOT_11252( .ZN(II36486), .A(g27507) );
  INV_X1 NOT_11253( .ZN(g27999), .A(II36486) );
  INV_X1 NOT_11254( .ZN(II36490), .A(g27265) );
  INV_X1 NOT_11255( .ZN(g28003), .A(II36490) );
  INV_X1 NOT_11256( .ZN(II36493), .A(g27266) );
  INV_X1 NOT_11257( .ZN(g28004), .A(II36493) );
  INV_X1 NOT_11258( .ZN(II36496), .A(g27267) );
  INV_X1 NOT_11259( .ZN(g28005), .A(II36496) );
  INV_X1 NOT_11260( .ZN(II36499), .A(g27268) );
  INV_X1 NOT_11261( .ZN(g28006), .A(II36499) );
  INV_X1 NOT_11262( .ZN(II36502), .A(g27269) );
  INV_X1 NOT_11263( .ZN(g28007), .A(II36502) );
  INV_X1 NOT_11264( .ZN(II36507), .A(g27270) );
  INV_X1 NOT_11265( .ZN(g28010), .A(II36507) );
  INV_X1 NOT_11266( .ZN(II36510), .A(g27271) );
  INV_X1 NOT_11267( .ZN(g28011), .A(II36510) );
  INV_X1 NOT_11268( .ZN(II36513), .A(g27272) );
  INV_X1 NOT_11269( .ZN(g28012), .A(II36513) );
  INV_X1 NOT_11270( .ZN(II36516), .A(g27273) );
  INV_X1 NOT_11271( .ZN(g28013), .A(II36516) );
  INV_X1 NOT_11272( .ZN(g28014), .A(g27373) );
  INV_X1 NOT_11273( .ZN(II36521), .A(g27274) );
  INV_X1 NOT_11274( .ZN(g28016), .A(II36521) );
  INV_X1 NOT_11275( .ZN(II36524), .A(g27275) );
  INV_X1 NOT_11276( .ZN(g28017), .A(II36524) );
  INV_X1 NOT_11277( .ZN(II36527), .A(g27524) );
  INV_X1 NOT_11278( .ZN(g28018), .A(II36527) );
  INV_X1 NOT_11279( .ZN(II36530), .A(g27276) );
  INV_X1 NOT_11280( .ZN(g28021), .A(II36530) );
  INV_X1 NOT_11281( .ZN(II36533), .A(g27277) );
  INV_X1 NOT_11282( .ZN(g28022), .A(II36533) );
  INV_X1 NOT_11283( .ZN(II36536), .A(g27278) );
  INV_X1 NOT_11284( .ZN(g28023), .A(II36536) );
  INV_X1 NOT_11285( .ZN(II36539), .A(g27279) );
  INV_X1 NOT_11286( .ZN(g28024), .A(II36539) );
  INV_X1 NOT_11287( .ZN(II36542), .A(g27280) );
  INV_X1 NOT_11288( .ZN(g28025), .A(II36542) );
  INV_X1 NOT_11289( .ZN(II36545), .A(g27281) );
  INV_X1 NOT_11290( .ZN(g28026), .A(II36545) );
  INV_X1 NOT_11291( .ZN(II36551), .A(g27282) );
  INV_X1 NOT_11292( .ZN(g28030), .A(II36551) );
  INV_X1 NOT_11293( .ZN(II36554), .A(g27283) );
  INV_X1 NOT_11294( .ZN(g28031), .A(II36554) );
  INV_X1 NOT_11295( .ZN(II36557), .A(g27284) );
  INV_X1 NOT_11296( .ZN(g28032), .A(II36557) );
  INV_X1 NOT_11297( .ZN(II36560), .A(g27285) );
  INV_X1 NOT_11298( .ZN(g28033), .A(II36560) );
  INV_X1 NOT_11299( .ZN(II36563), .A(g27286) );
  INV_X1 NOT_11300( .ZN(g28034), .A(II36563) );
  INV_X1 NOT_11301( .ZN(II36568), .A(g27287) );
  INV_X1 NOT_11302( .ZN(g28037), .A(II36568) );
  INV_X1 NOT_11303( .ZN(II36571), .A(g27288) );
  INV_X1 NOT_11304( .ZN(g28038), .A(II36571) );
  INV_X1 NOT_11305( .ZN(II36574), .A(g27289) );
  INV_X1 NOT_11306( .ZN(g28039), .A(II36574) );
  INV_X1 NOT_11307( .ZN(II36577), .A(g27290) );
  INV_X1 NOT_11308( .ZN(g28040), .A(II36577) );
  INV_X1 NOT_11309( .ZN(g28041), .A(g27376) );
  INV_X1 NOT_11310( .ZN(II36582), .A(g27291) );
  INV_X1 NOT_11311( .ZN(g28043), .A(II36582) );
  INV_X1 NOT_11312( .ZN(II36585), .A(g27292) );
  INV_X1 NOT_11313( .ZN(g28044), .A(II36585) );
  INV_X1 NOT_11314( .ZN(II36588), .A(g27293) );
  INV_X1 NOT_11315( .ZN(g28045), .A(II36588) );
  INV_X1 NOT_11316( .ZN(II36598), .A(g27294) );
  INV_X1 NOT_11317( .ZN(g28047), .A(II36598) );
  INV_X1 NOT_11318( .ZN(II36601), .A(g27295) );
  INV_X1 NOT_11319( .ZN(g28048), .A(II36601) );
  INV_X1 NOT_11320( .ZN(II36604), .A(g27296) );
  INV_X1 NOT_11321( .ZN(g28049), .A(II36604) );
  INV_X1 NOT_11322( .ZN(II36609), .A(g27297) );
  INV_X1 NOT_11323( .ZN(g28052), .A(II36609) );
  INV_X1 NOT_11324( .ZN(II36612), .A(g27298) );
  INV_X1 NOT_11325( .ZN(g28053), .A(II36612) );
  INV_X1 NOT_11326( .ZN(II36615), .A(g27299) );
  INV_X4 NOT_11327( .ZN(g28054), .A(II36615) );
  INV_X4 NOT_11328( .ZN(II36618), .A(g27300) );
  INV_X1 NOT_11329( .ZN(g28055), .A(II36618) );
  INV_X1 NOT_11330( .ZN(II36621), .A(g27301) );
  INV_X1 NOT_11331( .ZN(g28056), .A(II36621) );
  INV_X1 NOT_11332( .ZN(II36627), .A(g27302) );
  INV_X1 NOT_11333( .ZN(g28060), .A(II36627) );
  INV_X1 NOT_11334( .ZN(II36630), .A(g27303) );
  INV_X1 NOT_11335( .ZN(g28061), .A(II36630) );
  INV_X1 NOT_11336( .ZN(II36633), .A(g27304) );
  INV_X1 NOT_11337( .ZN(g28062), .A(II36633) );
  INV_X1 NOT_11338( .ZN(II36636), .A(g27305) );
  INV_X1 NOT_11339( .ZN(g28063), .A(II36636) );
  INV_X1 NOT_11340( .ZN(II36639), .A(g27306) );
  INV_X1 NOT_11341( .ZN(g28064), .A(II36639) );
  INV_X1 NOT_11342( .ZN(II36644), .A(g27307) );
  INV_X1 NOT_11343( .ZN(g28067), .A(II36644) );
  INV_X1 NOT_11344( .ZN(II36647), .A(g27308) );
  INV_X1 NOT_11345( .ZN(g28068), .A(II36647) );
  INV_X1 NOT_11346( .ZN(II36650), .A(g27309) );
  INV_X1 NOT_11347( .ZN(g28069), .A(II36650) );
  INV_X1 NOT_11348( .ZN(II36653), .A(g27310) );
  INV_X1 NOT_11349( .ZN(g28070), .A(II36653) );
  INV_X1 NOT_11350( .ZN(II36656), .A(g27311) );
  INV_X1 NOT_11351( .ZN(g28071), .A(II36656) );
  INV_X1 NOT_11352( .ZN(II36659), .A(g27312) );
  INV_X1 NOT_11353( .ZN(g28072), .A(II36659) );
  INV_X1 NOT_11354( .ZN(II36663), .A(g27313) );
  INV_X1 NOT_11355( .ZN(g28074), .A(II36663) );
  INV_X1 NOT_11356( .ZN(II36673), .A(g27314) );
  INV_X1 NOT_11357( .ZN(g28076), .A(II36673) );
  INV_X1 NOT_11358( .ZN(II36676), .A(g27315) );
  INV_X1 NOT_11359( .ZN(g28077), .A(II36676) );
  INV_X1 NOT_11360( .ZN(II36679), .A(g27316) );
  INV_X1 NOT_11361( .ZN(g28078), .A(II36679) );
  INV_X1 NOT_11362( .ZN(II36684), .A(g27317) );
  INV_X1 NOT_11363( .ZN(g28081), .A(II36684) );
  INV_X1 NOT_11364( .ZN(II36687), .A(g27318) );
  INV_X1 NOT_11365( .ZN(g28082), .A(II36687) );
  INV_X1 NOT_11366( .ZN(II36690), .A(g27319) );
  INV_X1 NOT_11367( .ZN(g28083), .A(II36690) );
  INV_X1 NOT_11368( .ZN(II36693), .A(g27320) );
  INV_X1 NOT_11369( .ZN(g28084), .A(II36693) );
  INV_X1 NOT_11370( .ZN(II36696), .A(g27321) );
  INV_X1 NOT_11371( .ZN(g28085), .A(II36696) );
  INV_X1 NOT_11372( .ZN(II36702), .A(g27322) );
  INV_X1 NOT_11373( .ZN(g28089), .A(II36702) );
  INV_X1 NOT_11374( .ZN(II36705), .A(g27323) );
  INV_X1 NOT_11375( .ZN(g28090), .A(II36705) );
  INV_X1 NOT_11376( .ZN(II36708), .A(g27324) );
  INV_X1 NOT_11377( .ZN(g28091), .A(II36708) );
  INV_X1 NOT_11378( .ZN(II36711), .A(g27325) );
  INV_X1 NOT_11379( .ZN(g28092), .A(II36711) );
  INV_X1 NOT_11380( .ZN(II36714), .A(g27326) );
  INV_X1 NOT_11381( .ZN(g28093), .A(II36714) );
  INV_X1 NOT_11382( .ZN(II36718), .A(g27327) );
  INV_X1 NOT_11383( .ZN(g28095), .A(II36718) );
  INV_X1 NOT_11384( .ZN(II36721), .A(g27328) );
  INV_X1 NOT_11385( .ZN(g28096), .A(II36721) );
  INV_X1 NOT_11386( .ZN(II36724), .A(g27329) );
  INV_X1 NOT_11387( .ZN(g28097), .A(II36724) );
  INV_X1 NOT_11388( .ZN(II36728), .A(g27330) );
  INV_X1 NOT_11389( .ZN(g28099), .A(II36728) );
  INV_X1 NOT_11390( .ZN(II36738), .A(g27331) );
  INV_X1 NOT_11391( .ZN(g28101), .A(II36738) );
  INV_X1 NOT_11392( .ZN(II36741), .A(g27332) );
  INV_X1 NOT_11393( .ZN(g28102), .A(II36741) );
  INV_X1 NOT_11394( .ZN(II36744), .A(g27333) );
  INV_X1 NOT_11395( .ZN(g28103), .A(II36744) );
  INV_X1 NOT_11396( .ZN(II36749), .A(g27334) );
  INV_X1 NOT_11397( .ZN(g28106), .A(II36749) );
  INV_X1 NOT_11398( .ZN(II36752), .A(g27335) );
  INV_X1 NOT_11399( .ZN(g28107), .A(II36752) );
  INV_X1 NOT_11400( .ZN(II36755), .A(g27336) );
  INV_X1 NOT_11401( .ZN(g28108), .A(II36755) );
  INV_X1 NOT_11402( .ZN(II36758), .A(g27337) );
  INV_X1 NOT_11403( .ZN(g28109), .A(II36758) );
  INV_X1 NOT_11404( .ZN(II36761), .A(g27338) );
  INV_X1 NOT_11405( .ZN(g28110), .A(II36761) );
  INV_X1 NOT_11406( .ZN(II36766), .A(g27339) );
  INV_X1 NOT_11407( .ZN(g28113), .A(II36766) );
  INV_X1 NOT_11408( .ZN(II36769), .A(g27340) );
  INV_X1 NOT_11409( .ZN(g28114), .A(II36769) );
  INV_X1 NOT_11410( .ZN(II36772), .A(g27341) );
  INV_X1 NOT_11411( .ZN(g28115), .A(II36772) );
  INV_X1 NOT_11412( .ZN(II36776), .A(g27342) );
  INV_X1 NOT_11413( .ZN(g28117), .A(II36776) );
  INV_X1 NOT_11414( .ZN(II36786), .A(g27343) );
  INV_X1 NOT_11415( .ZN(g28119), .A(II36786) );
  INV_X1 NOT_11416( .ZN(II36789), .A(g27344) );
  INV_X1 NOT_11417( .ZN(g28120), .A(II36789) );
  INV_X1 NOT_11418( .ZN(II36792), .A(g27345) );
  INV_X1 NOT_11419( .ZN(g28121), .A(II36792) );
  INV_X1 NOT_11420( .ZN(II36797), .A(g27346) );
  INV_X1 NOT_11421( .ZN(g28124), .A(II36797) );
  INV_X1 NOT_11422( .ZN(II36800), .A(g27347) );
  INV_X1 NOT_11423( .ZN(g28125), .A(II36800) );
  INV_X1 NOT_11424( .ZN(II36803), .A(g27348) );
  INV_X1 NOT_11425( .ZN(g28126), .A(II36803) );
  INV_X1 NOT_11426( .ZN(g28128), .A(g27528) );
  INV_X1 NOT_11427( .ZN(II36808), .A(g27354) );
  INV_X1 NOT_11428( .ZN(g28132), .A(II36808) );
  INV_X1 NOT_11429( .ZN(g28133), .A(g27550) );
  INV_X1 NOT_11430( .ZN(g28137), .A(g27566) );
  INV_X1 NOT_11431( .ZN(g28141), .A(g27576) );
  INV_X1 NOT_11432( .ZN(g28149), .A(g27667) );
  INV_X1 NOT_11433( .ZN(g28150), .A(g27387) );
  INV_X1 NOT_11434( .ZN(g28151), .A(g27381) );
  INV_X1 NOT_11435( .ZN(g28152), .A(g27391) );
  INV_X1 NOT_11436( .ZN(g28153), .A(g27397) );
  INV_X1 NOT_11437( .ZN(g28154), .A(g27401) );
  INV_X1 NOT_11438( .ZN(g28155), .A(g27404) );
  INV_X1 NOT_11439( .ZN(g28156), .A(g27410) );
  INV_X1 NOT_11440( .ZN(g28158), .A(g27416) );
  INV_X1 NOT_11441( .ZN(g28159), .A(g27419) );
  INV_X1 NOT_11442( .ZN(g28160), .A(g27422) );
  INV_X1 NOT_11443( .ZN(g28161), .A(g27428) );
  INV_X1 NOT_11444( .ZN(g28162), .A(g27432) );
  INV_X1 NOT_11445( .ZN(g28163), .A(g27437) );
  INV_X1 NOT_11446( .ZN(g28164), .A(g27440) );
  INV_X1 NOT_11447( .ZN(g28165), .A(g27443) );
  INV_X1 NOT_11448( .ZN(g28166), .A(g27451) );
  INV_X1 NOT_11449( .ZN(g28167), .A(g27456) );
  INV_X1 NOT_11450( .ZN(g28168), .A(g27459) );
  INV_X1 NOT_11451( .ZN(g28169), .A(g27467) );
  INV_X1 NOT_11452( .ZN(g28170), .A(g27472) );
  INV_X1 NOT_11453( .ZN(g28172), .A(g27475) );
  INV_X1 NOT_11454( .ZN(g28173), .A(g27486) );
  INV_X1 NOT_11455( .ZN(g28174), .A(g27489) );
  INV_X1 NOT_11456( .ZN(g28175), .A(g27498) );
  INV_X1 NOT_11457( .ZN(g28177), .A(g27510) );
  INV_X1 NOT_11458( .ZN(g28178), .A(g27518) );
  INV_X1 NOT_11459( .ZN(II36848), .A(g27383) );
  INV_X1 NOT_11460( .ZN(g28179), .A(II36848) );
  INV_X1 NOT_11461( .ZN(g28186), .A(g27535) );
  INV_X1 NOT_11462( .ZN(g28187), .A(g27543) );
  INV_X1 NOT_11463( .ZN(g28190), .A(g27555) );
  INV_X1 NOT_11464( .ZN(II36860), .A(g27386) );
  INV_X1 NOT_11465( .ZN(g28194), .A(II36860) );
  INV_X1 NOT_11466( .ZN(II36864), .A(g27384) );
  INV_X1 NOT_11467( .ZN(g28200), .A(II36864) );
  INV_X1 NOT_11468( .ZN(II36867), .A(g27786) );
  INV_X1 NOT_11469( .ZN(g28206), .A(II36867) );
  INV_X1 NOT_11470( .ZN(II36870), .A(g27955) );
  INV_X1 NOT_11471( .ZN(g28207), .A(II36870) );
  INV_X1 NOT_11472( .ZN(II36873), .A(g27971) );
  INV_X1 NOT_11473( .ZN(g28208), .A(II36873) );
  INV_X1 NOT_11474( .ZN(II36876), .A(g27986) );
  INV_X1 NOT_11475( .ZN(g28209), .A(II36876) );
  INV_X1 NOT_11476( .ZN(II36879), .A(g27972) );
  INV_X1 NOT_11477( .ZN(g28210), .A(II36879) );
  INV_X1 NOT_11478( .ZN(II36882), .A(g27987) );
  INV_X1 NOT_11479( .ZN(g28211), .A(II36882) );
  INV_X1 NOT_11480( .ZN(II36885), .A(g28003) );
  INV_X1 NOT_11481( .ZN(g28212), .A(II36885) );
  INV_X1 NOT_11482( .ZN(II36888), .A(g27988) );
  INV_X1 NOT_11483( .ZN(g28213), .A(II36888) );
  INV_X1 NOT_11484( .ZN(II36891), .A(g28004) );
  INV_X1 NOT_11485( .ZN(g28214), .A(II36891) );
  INV_X1 NOT_11486( .ZN(II36894), .A(g28022) );
  INV_X1 NOT_11487( .ZN(g28215), .A(II36894) );
  INV_X1 NOT_11488( .ZN(II36897), .A(g28005) );
  INV_X1 NOT_11489( .ZN(g28216), .A(II36897) );
  INV_X1 NOT_11490( .ZN(II36900), .A(g28023) );
  INV_X1 NOT_11491( .ZN(g28217), .A(II36900) );
  INV_X1 NOT_11492( .ZN(II36903), .A(g28045) );
  INV_X1 NOT_11493( .ZN(g28218), .A(II36903) );
  INV_X1 NOT_11494( .ZN(II36906), .A(g27989) );
  INV_X1 NOT_11495( .ZN(g28219), .A(II36906) );
  INV_X1 NOT_11496( .ZN(II36909), .A(g28006) );
  INV_X1 NOT_11497( .ZN(g28220), .A(II36909) );
  INV_X1 NOT_11498( .ZN(II36912), .A(g28024) );
  INV_X1 NOT_11499( .ZN(g28221), .A(II36912) );
  INV_X1 NOT_11500( .ZN(II36915), .A(g28007) );
  INV_X1 NOT_11501( .ZN(g28222), .A(II36915) );
  INV_X1 NOT_11502( .ZN(II36918), .A(g28025) );
  INV_X1 NOT_11503( .ZN(g28223), .A(II36918) );
  INV_X1 NOT_11504( .ZN(II36921), .A(g28047) );
  INV_X1 NOT_11505( .ZN(g28224), .A(II36921) );
  INV_X1 NOT_11506( .ZN(II36924), .A(g28026) );
  INV_X1 NOT_11507( .ZN(g28225), .A(II36924) );
  INV_X1 NOT_11508( .ZN(II36927), .A(g28048) );
  INV_X1 NOT_11509( .ZN(g28226), .A(II36927) );
  INV_X1 NOT_11510( .ZN(II36930), .A(g28071) );
  INV_X4 NOT_11511( .ZN(g28227), .A(II36930) );
  INV_X1 NOT_11512( .ZN(II36933), .A(g28049) );
  INV_X1 NOT_11513( .ZN(g28228), .A(II36933) );
  INV_X1 NOT_11514( .ZN(II36936), .A(g28072) );
  INV_X1 NOT_11515( .ZN(g28229), .A(II36936) );
  INV_X1 NOT_11516( .ZN(II36939), .A(g28095) );
  INV_X1 NOT_11517( .ZN(g28230), .A(II36939) );
  INV_X1 NOT_11518( .ZN(II36942), .A(g27905) );
  INV_X1 NOT_11519( .ZN(g28231), .A(II36942) );
  INV_X1 NOT_11520( .ZN(II36945), .A(g27793) );
  INV_X1 NOT_11521( .ZN(g28232), .A(II36945) );
  INV_X1 NOT_11522( .ZN(II36948), .A(g27976) );
  INV_X1 NOT_11523( .ZN(g28233), .A(II36948) );
  INV_X1 NOT_11524( .ZN(II36951), .A(g27992) );
  INV_X1 NOT_11525( .ZN(g28234), .A(II36951) );
  INV_X1 NOT_11526( .ZN(II36954), .A(g28010) );
  INV_X1 NOT_11527( .ZN(g28235), .A(II36954) );
  INV_X1 NOT_11528( .ZN(II36957), .A(g27993) );
  INV_X1 NOT_11529( .ZN(g28236), .A(II36957) );
  INV_X1 NOT_11530( .ZN(II36960), .A(g28011) );
  INV_X1 NOT_11531( .ZN(g28237), .A(II36960) );
  INV_X1 NOT_11532( .ZN(II36963), .A(g28030) );
  INV_X1 NOT_11533( .ZN(g28238), .A(II36963) );
  INV_X1 NOT_11534( .ZN(II36966), .A(g28012) );
  INV_X1 NOT_11535( .ZN(g28239), .A(II36966) );
  INV_X1 NOT_11536( .ZN(II36969), .A(g28031) );
  INV_X1 NOT_11537( .ZN(g28240), .A(II36969) );
  INV_X1 NOT_11538( .ZN(II36972), .A(g28052) );
  INV_X1 NOT_11539( .ZN(g28241), .A(II36972) );
  INV_X1 NOT_11540( .ZN(II36975), .A(g28032) );
  INV_X1 NOT_11541( .ZN(g28242), .A(II36975) );
  INV_X1 NOT_11542( .ZN(II36978), .A(g28053) );
  INV_X1 NOT_11543( .ZN(g28243), .A(II36978) );
  INV_X1 NOT_11544( .ZN(II36981), .A(g28074) );
  INV_X1 NOT_11545( .ZN(g28244), .A(II36981) );
  INV_X1 NOT_11546( .ZN(II36984), .A(g28013) );
  INV_X1 NOT_11547( .ZN(g28245), .A(II36984) );
  INV_X1 NOT_11548( .ZN(II36987), .A(g28033) );
  INV_X1 NOT_11549( .ZN(g28246), .A(II36987) );
  INV_X1 NOT_11550( .ZN(II36990), .A(g28054) );
  INV_X1 NOT_11551( .ZN(g28247), .A(II36990) );
  INV_X1 NOT_11552( .ZN(II36993), .A(g28034) );
  INV_X1 NOT_11553( .ZN(g28248), .A(II36993) );
  INV_X1 NOT_11554( .ZN(II36996), .A(g28055) );
  INV_X1 NOT_11555( .ZN(g28249), .A(II36996) );
  INV_X1 NOT_11556( .ZN(II36999), .A(g28076) );
  INV_X1 NOT_11557( .ZN(g28250), .A(II36999) );
  INV_X1 NOT_11558( .ZN(II37002), .A(g28056) );
  INV_X1 NOT_11559( .ZN(g28251), .A(II37002) );
  INV_X1 NOT_11560( .ZN(II37005), .A(g28077) );
  INV_X1 NOT_11561( .ZN(g28252), .A(II37005) );
  INV_X1 NOT_11562( .ZN(II37008), .A(g28096) );
  INV_X1 NOT_11563( .ZN(g28253), .A(II37008) );
  INV_X1 NOT_11564( .ZN(II37011), .A(g28078) );
  INV_X1 NOT_11565( .ZN(g28254), .A(II37011) );
  INV_X1 NOT_11566( .ZN(II37014), .A(g28097) );
  INV_X1 NOT_11567( .ZN(g28255), .A(II37014) );
  INV_X1 NOT_11568( .ZN(II37017), .A(g28113) );
  INV_X1 NOT_11569( .ZN(g28256), .A(II37017) );
  INV_X1 NOT_11570( .ZN(II37020), .A(g27910) );
  INV_X1 NOT_11571( .ZN(g28257), .A(II37020) );
  INV_X1 NOT_11572( .ZN(II37023), .A(g27799) );
  INV_X1 NOT_11573( .ZN(g28258), .A(II37023) );
  INV_X1 NOT_11574( .ZN(II37026), .A(g27998) );
  INV_X1 NOT_11575( .ZN(g28259), .A(II37026) );
  INV_X1 NOT_11576( .ZN(II37029), .A(g28016) );
  INV_X1 NOT_11577( .ZN(g28260), .A(II37029) );
  INV_X1 NOT_11578( .ZN(II37032), .A(g28037) );
  INV_X1 NOT_11579( .ZN(g28261), .A(II37032) );
  INV_X1 NOT_11580( .ZN(II37035), .A(g28017) );
  INV_X1 NOT_11581( .ZN(g28262), .A(II37035) );
  INV_X1 NOT_11582( .ZN(II37038), .A(g28038) );
  INV_X1 NOT_11583( .ZN(g28263), .A(II37038) );
  INV_X1 NOT_11584( .ZN(II37041), .A(g28060) );
  INV_X1 NOT_11585( .ZN(g28264), .A(II37041) );
  INV_X1 NOT_11586( .ZN(II37044), .A(g28039) );
  INV_X1 NOT_11587( .ZN(g28265), .A(II37044) );
  INV_X1 NOT_11588( .ZN(II37047), .A(g28061) );
  INV_X1 NOT_11589( .ZN(g28266), .A(II37047) );
  INV_X1 NOT_11590( .ZN(II37050), .A(g28081) );
  INV_X1 NOT_11591( .ZN(g28267), .A(II37050) );
  INV_X1 NOT_11592( .ZN(II37053), .A(g28062) );
  INV_X1 NOT_11593( .ZN(g28268), .A(II37053) );
  INV_X1 NOT_11594( .ZN(II37056), .A(g28082) );
  INV_X1 NOT_11595( .ZN(g28269), .A(II37056) );
  INV_X1 NOT_11596( .ZN(II37059), .A(g28099) );
  INV_X1 NOT_11597( .ZN(g28270), .A(II37059) );
  INV_X1 NOT_11598( .ZN(II37062), .A(g28040) );
  INV_X1 NOT_11599( .ZN(g28271), .A(II37062) );
  INV_X1 NOT_11600( .ZN(II37065), .A(g28063) );
  INV_X1 NOT_11601( .ZN(g28272), .A(II37065) );
  INV_X1 NOT_11602( .ZN(II37068), .A(g28083) );
  INV_X1 NOT_11603( .ZN(g28273), .A(II37068) );
  INV_X1 NOT_11604( .ZN(II37071), .A(g28064) );
  INV_X1 NOT_11605( .ZN(g28274), .A(II37071) );
  INV_X1 NOT_11606( .ZN(II37074), .A(g28084) );
  INV_X1 NOT_11607( .ZN(g28275), .A(II37074) );
  INV_X1 NOT_11608( .ZN(II37077), .A(g28101) );
  INV_X1 NOT_11609( .ZN(g28276), .A(II37077) );
  INV_X1 NOT_11610( .ZN(II37080), .A(g28085) );
  INV_X1 NOT_11611( .ZN(g28277), .A(II37080) );
  INV_X1 NOT_11612( .ZN(II37083), .A(g28102) );
  INV_X1 NOT_11613( .ZN(g28278), .A(II37083) );
  INV_X1 NOT_11614( .ZN(II37086), .A(g28114) );
  INV_X16 NOT_11615( .ZN(g28279), .A(II37086) );
  INV_X1 NOT_11616( .ZN(II37089), .A(g28103) );
  INV_X1 NOT_11617( .ZN(g28280), .A(II37089) );
  INV_X1 NOT_11618( .ZN(II37092), .A(g28115) );
  INV_X1 NOT_11619( .ZN(g28281), .A(II37092) );
  INV_X1 NOT_11620( .ZN(II37095), .A(g28124) );
  INV_X1 NOT_11621( .ZN(g28282), .A(II37095) );
  INV_X1 NOT_11622( .ZN(II37098), .A(g27918) );
  INV_X1 NOT_11623( .ZN(g28283), .A(II37098) );
  INV_X1 NOT_11624( .ZN(II37101), .A(g27805) );
  INV_X1 NOT_11625( .ZN(g28284), .A(II37101) );
  INV_X1 NOT_11626( .ZN(II37104), .A(g28021) );
  INV_X1 NOT_11627( .ZN(g28285), .A(II37104) );
  INV_X1 NOT_11628( .ZN(II37107), .A(g28043) );
  INV_X1 NOT_11629( .ZN(g28286), .A(II37107) );
  INV_X1 NOT_11630( .ZN(II37110), .A(g28067) );
  INV_X1 NOT_11631( .ZN(g28287), .A(II37110) );
  INV_X1 NOT_11632( .ZN(II37113), .A(g28044) );
  INV_X1 NOT_11633( .ZN(g28288), .A(II37113) );
  INV_X1 NOT_11634( .ZN(II37116), .A(g28068) );
  INV_X1 NOT_11635( .ZN(g28289), .A(II37116) );
  INV_X1 NOT_11636( .ZN(II37119), .A(g28089) );
  INV_X1 NOT_11637( .ZN(g28290), .A(II37119) );
  INV_X1 NOT_11638( .ZN(II37122), .A(g28069) );
  INV_X1 NOT_11639( .ZN(g28291), .A(II37122) );
  INV_X16 NOT_11640( .ZN(II37125), .A(g28090) );
  INV_X1 NOT_11641( .ZN(g28292), .A(II37125) );
  INV_X1 NOT_11642( .ZN(II37128), .A(g28106) );
  INV_X1 NOT_11643( .ZN(g28293), .A(II37128) );
  INV_X1 NOT_11644( .ZN(II37131), .A(g28091) );
  INV_X1 NOT_11645( .ZN(g28294), .A(II37131) );
  INV_X1 NOT_11646( .ZN(II37134), .A(g28107) );
  INV_X1 NOT_11647( .ZN(g28295), .A(II37134) );
  INV_X1 NOT_11648( .ZN(II37137), .A(g28117) );
  INV_X1 NOT_11649( .ZN(g28296), .A(II37137) );
  INV_X1 NOT_11650( .ZN(II37140), .A(g28070) );
  INV_X1 NOT_11651( .ZN(g28297), .A(II37140) );
  INV_X1 NOT_11652( .ZN(II37143), .A(g28092) );
  INV_X1 NOT_11653( .ZN(g28298), .A(II37143) );
  INV_X1 NOT_11654( .ZN(II37146), .A(g28108) );
  INV_X1 NOT_11655( .ZN(g28299), .A(II37146) );
  INV_X1 NOT_11656( .ZN(II37149), .A(g28093) );
  INV_X1 NOT_11657( .ZN(g28300), .A(II37149) );
  INV_X1 NOT_11658( .ZN(II37152), .A(g28109) );
  INV_X1 NOT_11659( .ZN(g28301), .A(II37152) );
  INV_X1 NOT_11660( .ZN(II37155), .A(g28119) );
  INV_X1 NOT_11661( .ZN(g28302), .A(II37155) );
  INV_X1 NOT_11662( .ZN(II37158), .A(g28110) );
  INV_X1 NOT_11663( .ZN(g28303), .A(II37158) );
  INV_X1 NOT_11664( .ZN(II37161), .A(g28120) );
  INV_X1 NOT_11665( .ZN(g28304), .A(II37161) );
  INV_X1 NOT_11666( .ZN(II37164), .A(g28125) );
  INV_X1 NOT_11667( .ZN(g28305), .A(II37164) );
  INV_X1 NOT_11668( .ZN(II37167), .A(g28121) );
  INV_X1 NOT_11669( .ZN(g28306), .A(II37167) );
  INV_X1 NOT_11670( .ZN(II37170), .A(g28126) );
  INV_X1 NOT_11671( .ZN(g28307), .A(II37170) );
  INV_X1 NOT_11672( .ZN(II37173), .A(g28132) );
  INV_X1 NOT_11673( .ZN(g28308), .A(II37173) );
  INV_X1 NOT_11674( .ZN(II37176), .A(g27927) );
  INV_X1 NOT_11675( .ZN(g28309), .A(II37176) );
  INV_X1 NOT_11676( .ZN(II37179), .A(g27784) );
  INV_X1 NOT_11677( .ZN(g28310), .A(II37179) );
  INV_X1 NOT_11678( .ZN(II37182), .A(g27791) );
  INV_X1 NOT_11679( .ZN(g28311), .A(II37182) );
  INV_X1 NOT_11680( .ZN(II37185), .A(g27797) );
  INV_X1 NOT_11681( .ZN(g28312), .A(II37185) );
  INV_X1 NOT_11682( .ZN(II37188), .A(g27785) );
  INV_X1 NOT_11683( .ZN(g28313), .A(II37188) );
  INV_X1 NOT_11684( .ZN(II37191), .A(g27792) );
  INV_X1 NOT_11685( .ZN(g28314), .A(II37191) );
  INV_X1 NOT_11686( .ZN(II37194), .A(g27800) );
  INV_X1 NOT_11687( .ZN(g28315), .A(II37194) );
  INV_X1 NOT_11688( .ZN(II37197), .A(g27903) );
  INV_X1 NOT_11689( .ZN(g28316), .A(II37197) );
  INV_X1 NOT_11690( .ZN(II37200), .A(g27907) );
  INV_X1 NOT_11691( .ZN(g28317), .A(II37200) );
  INV_X1 NOT_11692( .ZN(II37203), .A(g27912) );
  INV_X1 NOT_11693( .ZN(g28318), .A(II37203) );
  INV_X1 NOT_11694( .ZN(II37228), .A(g28194) );
  INV_X1 NOT_11695( .ZN(g28341), .A(II37228) );
  INV_X1 NOT_11696( .ZN(II37232), .A(g28200) );
  INV_X1 NOT_11697( .ZN(g28343), .A(II37232) );
  INV_X1 NOT_11698( .ZN(II37238), .A(g28179) );
  INV_X1 NOT_11699( .ZN(g28347), .A(II37238) );
  INV_X1 NOT_11700( .ZN(II37252), .A(g28200) );
  INV_X1 NOT_11701( .ZN(g28359), .A(II37252) );
  INV_X1 NOT_11702( .ZN(II37260), .A(g28179) );
  INV_X1 NOT_11703( .ZN(g28365), .A(II37260) );
  INV_X1 NOT_11704( .ZN(II37266), .A(g28200) );
  INV_X1 NOT_11705( .ZN(g28369), .A(II37266) );
  INV_X1 NOT_11706( .ZN(II37269), .A(g28145) );
  INV_X1 NOT_11707( .ZN(g28370), .A(II37269) );
  INV_X1 NOT_11708( .ZN(II37273), .A(g28179) );
  INV_X1 NOT_11709( .ZN(g28372), .A(II37273) );
  INV_X1 NOT_11710( .ZN(II37277), .A(g28146) );
  INV_X1 NOT_11711( .ZN(g28374), .A(II37277) );
  INV_X1 NOT_11712( .ZN(II37280), .A(g28179) );
  INV_X1 NOT_11713( .ZN(g28375), .A(II37280) );
  INV_X1 NOT_11714( .ZN(II37284), .A(g28147) );
  INV_X1 NOT_11715( .ZN(g28377), .A(II37284) );
  INV_X1 NOT_11716( .ZN(II37291), .A(g28148) );
  INV_X1 NOT_11717( .ZN(g28382), .A(II37291) );
  INV_X1 NOT_11718( .ZN(II37319), .A(g28149) );
  INV_X1 NOT_11719( .ZN(g28390), .A(II37319) );
  INV_X1 NOT_11720( .ZN(II37330), .A(g28194) );
  INV_X1 NOT_11721( .ZN(g28393), .A(II37330) );
  INV_X1 NOT_11722( .ZN(II37334), .A(g28194) );
  INV_X1 NOT_11723( .ZN(g28395), .A(II37334) );
  INV_X1 NOT_11724( .ZN(g28419), .A(g28151) );
  INV_X1 NOT_11725( .ZN(II37379), .A(g28199) );
  INV_X1 NOT_11726( .ZN(g28432), .A(II37379) );
  INV_X1 NOT_11727( .ZN(II37386), .A(g28194) );
  INV_X1 NOT_11728( .ZN(g28437), .A(II37386) );
  INV_X1 NOT_11729( .ZN(II37394), .A(g27718) );
  INV_X1 NOT_11730( .ZN(g28443), .A(II37394) );
  INV_X1 NOT_11731( .ZN(II37400), .A(g28200) );
  INV_X1 NOT_11732( .ZN(g28447), .A(II37400) );
  INV_X1 NOT_11733( .ZN(II37410), .A(g27722) );
  INV_X1 NOT_11734( .ZN(g28455), .A(II37410) );
  INV_X1 NOT_11735( .ZN(II37415), .A(g28179) );
  INV_X1 NOT_11736( .ZN(g28458), .A(II37415) );
  INV_X1 NOT_11737( .ZN(II37426), .A(g27724) );
  INV_X1 NOT_11738( .ZN(g28467), .A(II37426) );
  INV_X1 NOT_11739( .ZN(g28483), .A(g27776) );
  INV_X1 NOT_11740( .ZN(g28491), .A(g27780) );
  INV_X1 NOT_11741( .ZN(g28496), .A(g27787) );
  INV_X1 NOT_11742( .ZN(II37459), .A(g27759) );
  INV_X1 NOT_11743( .ZN(g28498), .A(II37459) );
  INV_X1 NOT_11744( .ZN(g28500), .A(g27794) );
  INV_X1 NOT_11745( .ZN(II37467), .A(g27760) );
  INV_X1 NOT_11746( .ZN(g28524), .A(II37467) );
  INV_X1 NOT_11747( .ZN(II37471), .A(g27761) );
  INV_X1 NOT_11748( .ZN(g28526), .A(II37471) );
  INV_X1 NOT_11749( .ZN(II37474), .A(g27762) );
  INV_X1 NOT_11750( .ZN(g28527), .A(II37474) );
  INV_X1 NOT_11751( .ZN(II37481), .A(g27763) );
  INV_X1 NOT_11752( .ZN(g28552), .A(II37481) );
  INV_X1 NOT_11753( .ZN(II37484), .A(g27764) );
  INV_X1 NOT_11754( .ZN(g28553), .A(II37484) );
  INV_X1 NOT_11755( .ZN(g28554), .A(g27806) );
  INV_X1 NOT_11756( .ZN(II37488), .A(g27765) );
  INV_X1 NOT_11757( .ZN(g28555), .A(II37488) );
  INV_X1 NOT_11758( .ZN(II37494), .A(g27766) );
  INV_X1 NOT_11759( .ZN(g28579), .A(II37494) );
  INV_X1 NOT_11760( .ZN(II37497), .A(g27767) );
  INV_X1 NOT_11761( .ZN(g28580), .A(II37497) );
  INV_X1 NOT_11762( .ZN(g28581), .A(g27817) );
  INV_X1 NOT_11763( .ZN(g28582), .A(g27820) );
  INV_X1 NOT_11764( .ZN(II37502), .A(g27768) );
  INV_X1 NOT_11765( .ZN(g28583), .A(II37502) );
  INV_X1 NOT_11766( .ZN(II37508), .A(g27769) );
  INV_X1 NOT_11767( .ZN(g28607), .A(II37508) );
  INV_X1 NOT_11768( .ZN(g28608), .A(g27831) );
  INV_X1 NOT_11769( .ZN(g28609), .A(g27839) );
  INV_X1 NOT_11770( .ZN(g28610), .A(g27843) );
  INV_X1 NOT_11771( .ZN(II37514), .A(g27771) );
  INV_X1 NOT_11772( .ZN(g28611), .A(II37514) );
  INV_X1 NOT_11773( .ZN(g28612), .A(g28046) );
  INV_X1 NOT_11774( .ZN(g28616), .A(g27847) );
  INV_X1 NOT_11775( .ZN(g28617), .A(g27858) );
  INV_X1 NOT_11776( .ZN(g28618), .A(g27861) );
  INV_X1 NOT_11777( .ZN(g28619), .A(g28075) );
  INV_X1 NOT_11778( .ZN(g28623), .A(g27872) );
  INV_X1 NOT_11779( .ZN(g28624), .A(g27879) );
  INV_X1 NOT_11780( .ZN(g28625), .A(g28100) );
  INV_X1 NOT_11781( .ZN(g28629), .A(g27889) );
  INV_X1 NOT_11782( .ZN(g28630), .A(g28118) );
  INV_X1 NOT_11783( .ZN(g28638), .A(g28200) );
  INV_X1 NOT_11784( .ZN(g28639), .A(g27919) );
  INV_X1 NOT_11785( .ZN(g28640), .A(g27928) );
  INV_X1 NOT_11786( .ZN(g28641), .A(g27932) );
  INV_X1 NOT_11787( .ZN(g28642), .A(g27939) );
  INV_X1 NOT_11788( .ZN(g28643), .A(g27942) );
  INV_X1 NOT_11789( .ZN(g28644), .A(g27946) );
  INV_X1 NOT_11790( .ZN(g28645), .A(g27952) );
  INV_X1 NOT_11791( .ZN(g28646), .A(g27956) );
  INV_X1 NOT_11792( .ZN(g28647), .A(g27959) );
  INV_X1 NOT_11793( .ZN(g28648), .A(g27965) );
  INV_X1 NOT_11794( .ZN(g28649), .A(g27973) );
  INV_X1 NOT_11795( .ZN(g28650), .A(g27977) );
  INV_X1 NOT_11796( .ZN(g28651), .A(g27981) );
  INV_X1 NOT_11797( .ZN(g28652), .A(g27994) );
  INV_X1 NOT_11798( .ZN(g28653), .A(g27999) );
  INV_X1 NOT_11799( .ZN(g28655), .A(g28018) );
  INV_X1 NOT_11800( .ZN(II37566), .A(g28370) );
  INV_X1 NOT_11801( .ZN(g28673), .A(II37566) );
  INV_X1 NOT_11802( .ZN(II37569), .A(g28498) );
  INV_X1 NOT_11803( .ZN(g28674), .A(II37569) );
  INV_X1 NOT_11804( .ZN(II37572), .A(g28524) );
  INV_X1 NOT_11805( .ZN(g28675), .A(II37572) );
  INV_X1 NOT_11806( .ZN(II37575), .A(g28527) );
  INV_X1 NOT_11807( .ZN(g28676), .A(II37575) );
  INV_X16 NOT_11808( .ZN(II37578), .A(g28432) );
  INV_X16 NOT_11809( .ZN(g28677), .A(II37578) );
  INV_X1 NOT_11810( .ZN(II37581), .A(g28374) );
  INV_X1 NOT_11811( .ZN(g28678), .A(II37581) );
  INV_X1 NOT_11812( .ZN(II37584), .A(g28526) );
  INV_X1 NOT_11813( .ZN(g28679), .A(II37584) );
  INV_X1 NOT_11814( .ZN(II37587), .A(g28552) );
  INV_X1 NOT_11815( .ZN(g28680), .A(II37587) );
  INV_X1 NOT_11816( .ZN(II37590), .A(g28555) );
  INV_X1 NOT_11817( .ZN(g28681), .A(II37590) );
  INV_X1 NOT_11818( .ZN(II37593), .A(g28443) );
  INV_X1 NOT_11819( .ZN(g28682), .A(II37593) );
  INV_X1 NOT_11820( .ZN(II37596), .A(g28377) );
  INV_X1 NOT_11821( .ZN(g28683), .A(II37596) );
  INV_X1 NOT_11822( .ZN(II37599), .A(g28553) );
  INV_X1 NOT_11823( .ZN(g28684), .A(II37599) );
  INV_X1 NOT_11824( .ZN(II37602), .A(g28579) );
  INV_X1 NOT_11825( .ZN(g28685), .A(II37602) );
  INV_X1 NOT_11826( .ZN(II37605), .A(g28583) );
  INV_X1 NOT_11827( .ZN(g28686), .A(II37605) );
  INV_X1 NOT_11828( .ZN(II37608), .A(g28455) );
  INV_X1 NOT_11829( .ZN(g28687), .A(II37608) );
  INV_X1 NOT_11830( .ZN(II37611), .A(g28382) );
  INV_X1 NOT_11831( .ZN(g28688), .A(II37611) );
  INV_X1 NOT_11832( .ZN(II37614), .A(g28580) );
  INV_X1 NOT_11833( .ZN(g28689), .A(II37614) );
  INV_X1 NOT_11834( .ZN(II37617), .A(g28607) );
  INV_X1 NOT_11835( .ZN(g28690), .A(II37617) );
  INV_X1 NOT_11836( .ZN(II37620), .A(g28611) );
  INV_X1 NOT_11837( .ZN(g28691), .A(II37620) );
  INV_X1 NOT_11838( .ZN(II37623), .A(g28467) );
  INV_X1 NOT_11839( .ZN(g28692), .A(II37623) );
  INV_X1 NOT_11840( .ZN(II37626), .A(g28393) );
  INV_X1 NOT_11841( .ZN(g28693), .A(II37626) );
  INV_X1 NOT_11842( .ZN(II37629), .A(g28369) );
  INV_X1 NOT_11843( .ZN(g28694), .A(II37629) );
  INV_X1 NOT_11844( .ZN(II37632), .A(g28372) );
  INV_X1 NOT_11845( .ZN(g28695), .A(II37632) );
  INV_X1 NOT_11846( .ZN(II37635), .A(g28390) );
  INV_X1 NOT_11847( .ZN(g28696), .A(II37635) );
  INV_X1 NOT_11848( .ZN(II37638), .A(g28395) );
  INV_X1 NOT_11849( .ZN(g28697), .A(II37638) );
  INV_X1 NOT_11850( .ZN(II37641), .A(g28375) );
  INV_X1 NOT_11851( .ZN(g28698), .A(II37641) );
  INV_X1 NOT_11852( .ZN(II37644), .A(g28341) );
  INV_X1 NOT_11853( .ZN(g28699), .A(II37644) );
  INV_X1 NOT_11854( .ZN(II37647), .A(g28343) );
  INV_X1 NOT_11855( .ZN(g28700), .A(II37647) );
  INV_X1 NOT_11856( .ZN(II37650), .A(g28347) );
  INV_X1 NOT_11857( .ZN(g28701), .A(II37650) );
  INV_X1 NOT_11858( .ZN(II37653), .A(g28359) );
  INV_X1 NOT_11859( .ZN(g28702), .A(II37653) );
  INV_X1 NOT_11860( .ZN(II37656), .A(g28365) );
  INV_X1 NOT_11861( .ZN(g28703), .A(II37656) );
  INV_X1 NOT_11862( .ZN(II37659), .A(g28437) );
  INV_X1 NOT_11863( .ZN(g28704), .A(II37659) );
  INV_X1 NOT_11864( .ZN(II37662), .A(g28447) );
  INV_X1 NOT_11865( .ZN(g28705), .A(II37662) );
  INV_X1 NOT_11866( .ZN(II37665), .A(g28458) );
  INV_X1 NOT_11867( .ZN(g28706), .A(II37665) );
  INV_X1 NOT_11868( .ZN(g28720), .A(g28495) );
  INV_X1 NOT_11869( .ZN(g28721), .A(g28490) );
  INV_X1 NOT_11870( .ZN(g28723), .A(g28528) );
  INV_X1 NOT_11871( .ZN(g28725), .A(g28499) );
  INV_X1 NOT_11872( .ZN(g28727), .A(g28489) );
  INV_X1 NOT_11873( .ZN(g28730), .A(g28470) );
  INV_X1 NOT_11874( .ZN(g28734), .A(g28525) );
  INV_X1 NOT_11875( .ZN(g28740), .A(g28488) );
  INV_X1 NOT_11876( .ZN(II37702), .A(g28512) );
  INV_X1 NOT_11877( .ZN(g28741), .A(II37702) );
  INV_X1 NOT_11878( .ZN(II37712), .A(g28512) );
  INV_X1 NOT_11879( .ZN(g28751), .A(II37712) );
  INV_X1 NOT_11880( .ZN(II37716), .A(g28540) );
  INV_X1 NOT_11881( .ZN(g28755), .A(II37716) );
  INV_X1 NOT_11882( .ZN(II37725), .A(g28540) );
  INV_X1 NOT_11883( .ZN(g28764), .A(II37725) );
  INV_X1 NOT_11884( .ZN(II37729), .A(g28567) );
  INV_X1 NOT_11885( .ZN(g28768), .A(II37729) );
  INV_X1 NOT_11886( .ZN(II37736), .A(g28567) );
  INV_X1 NOT_11887( .ZN(g28775), .A(II37736) );
  INV_X1 NOT_11888( .ZN(II37740), .A(g28595) );
  INV_X1 NOT_11889( .ZN(g28779), .A(II37740) );
  INV_X1 NOT_11890( .ZN(II37746), .A(g28595) );
  INV_X1 NOT_11891( .ZN(g28785), .A(II37746) );
  INV_X1 NOT_11892( .ZN(II37752), .A(g28512) );
  INV_X1 NOT_11893( .ZN(g28791), .A(II37752) );
  INV_X1 NOT_11894( .ZN(II37757), .A(g28512) );
  INV_X1 NOT_11895( .ZN(g28796), .A(II37757) );
  INV_X1 NOT_11896( .ZN(II37760), .A(g28540) );
  INV_X1 NOT_11897( .ZN(g28799), .A(II37760) );
  INV_X1 NOT_11898( .ZN(II37765), .A(g28512) );
  INV_X1 NOT_11899( .ZN(g28804), .A(II37765) );
  INV_X1 NOT_11900( .ZN(II37768), .A(g28540) );
  INV_X1 NOT_11901( .ZN(g28807), .A(II37768) );
  INV_X1 NOT_11902( .ZN(II37771), .A(g28567) );
  INV_X1 NOT_11903( .ZN(g28810), .A(II37771) );
  INV_X1 NOT_11904( .ZN(II37775), .A(g28540) );
  INV_X1 NOT_11905( .ZN(g28814), .A(II37775) );
  INV_X1 NOT_11906( .ZN(II37778), .A(g28567) );
  INV_X1 NOT_11907( .ZN(g28817), .A(II37778) );
  INV_X1 NOT_11908( .ZN(II37781), .A(g28595) );
  INV_X1 NOT_11909( .ZN(g28820), .A(II37781) );
  INV_X1 NOT_11910( .ZN(II37784), .A(g28567) );
  INV_X1 NOT_11911( .ZN(g28823), .A(II37784) );
  INV_X1 NOT_11912( .ZN(II37787), .A(g28595) );
  INV_X1 NOT_11913( .ZN(g28826), .A(II37787) );
  INV_X1 NOT_11914( .ZN(II37790), .A(g28595) );
  INV_X1 NOT_11915( .ZN(g28829), .A(II37790) );
  INV_X1 NOT_11916( .ZN(II37793), .A(g28638) );
  INV_X1 NOT_11917( .ZN(g28832), .A(II37793) );
  INV_X1 NOT_11918( .ZN(II37796), .A(g28634) );
  INV_X1 NOT_11919( .ZN(g28833), .A(II37796) );
  INV_X1 NOT_11920( .ZN(II37800), .A(g28635) );
  INV_X1 NOT_11921( .ZN(g28835), .A(II37800) );
  INV_X1 NOT_11922( .ZN(II37804), .A(g28636) );
  INV_X1 NOT_11923( .ZN(g28837), .A(II37804) );
  INV_X1 NOT_11924( .ZN(II37808), .A(g28637) );
  INV_X1 NOT_11925( .ZN(g28839), .A(II37808) );
  INV_X1 NOT_11926( .ZN(g28855), .A(g28409) );
  INV_X1 NOT_11927( .ZN(g28859), .A(g28413) );
  INV_X1 NOT_11928( .ZN(g28863), .A(g28417) );
  INV_X1 NOT_11929( .ZN(g28867), .A(g28418) );
  INV_X1 NOT_11930( .ZN(II37842), .A(g28501) );
  INV_X1 NOT_11931( .ZN(g28871), .A(II37842) );
  INV_X1 NOT_11932( .ZN(II37846), .A(g28501) );
  INV_X1 NOT_11933( .ZN(g28877), .A(II37846) );
  INV_X1 NOT_11934( .ZN(II37851), .A(g28668) );
  INV_X1 NOT_11935( .ZN(g28882), .A(II37851) );
  INV_X1 NOT_11936( .ZN(II37854), .A(g28529) );
  INV_X1 NOT_11937( .ZN(g28883), .A(II37854) );
  INV_X1 NOT_11938( .ZN(II37858), .A(g28501) );
  INV_X1 NOT_11939( .ZN(g28889), .A(II37858) );
  INV_X1 NOT_11940( .ZN(II37863), .A(g28529) );
  INV_X1 NOT_11941( .ZN(g28894), .A(II37863) );
  INV_X1 NOT_11942( .ZN(II37868), .A(g28321) );
  INV_X1 NOT_11943( .ZN(g28899), .A(II37868) );
  INV_X1 NOT_11944( .ZN(II37871), .A(g28556) );
  INV_X1 NOT_11945( .ZN(g28900), .A(II37871) );
  INV_X1 NOT_11946( .ZN(II37875), .A(g28501) );
  INV_X1 NOT_11947( .ZN(g28906), .A(II37875) );
  INV_X1 NOT_11948( .ZN(II37880), .A(g28529) );
  INV_X1 NOT_11949( .ZN(g28911), .A(II37880) );
  INV_X1 NOT_11950( .ZN(II37885), .A(g28556) );
  INV_X1 NOT_11951( .ZN(g28916), .A(II37885) );
  INV_X1 NOT_11952( .ZN(II37891), .A(g28325) );
  INV_X1 NOT_11953( .ZN(g28924), .A(II37891) );
  INV_X1 NOT_11954( .ZN(II37894), .A(g28584) );
  INV_X1 NOT_11955( .ZN(g28925), .A(II37894) );
  INV_X1 NOT_11956( .ZN(II37897), .A(g28501) );
  INV_X1 NOT_11957( .ZN(g28928), .A(II37897) );
  INV_X1 NOT_11958( .ZN(II37901), .A(g28529) );
  INV_X1 NOT_11959( .ZN(g28932), .A(II37901) );
  INV_X1 NOT_11960( .ZN(II37906), .A(g28556) );
  INV_X1 NOT_11961( .ZN(g28937), .A(II37906) );
  INV_X1 NOT_11962( .ZN(II37912), .A(g28584) );
  INV_X1 NOT_11963( .ZN(g28945), .A(II37912) );
  INV_X1 NOT_11964( .ZN(II37917), .A(g28328) );
  INV_X1 NOT_11965( .ZN(g28950), .A(II37917) );
  INV_X1 NOT_11966( .ZN(II37920), .A(g28501) );
  INV_X1 NOT_11967( .ZN(g28951), .A(II37920) );
  INV_X1 NOT_11968( .ZN(II37924), .A(g28529) );
  INV_X1 NOT_11969( .ZN(g28955), .A(II37924) );
  INV_X1 NOT_11970( .ZN(II37928), .A(g28556) );
  INV_X1 NOT_11971( .ZN(g28959), .A(II37928) );
  INV_X1 NOT_11972( .ZN(II37934), .A(g28584) );
  INV_X1 NOT_11973( .ZN(g28967), .A(II37934) );
  INV_X1 NOT_11974( .ZN(II37939), .A(g28501) );
  INV_X1 NOT_11975( .ZN(g28972), .A(II37939) );
  INV_X1 NOT_11976( .ZN(II37942), .A(g28501) );
  INV_X1 NOT_11977( .ZN(g28975), .A(II37942) );
  INV_X1 NOT_11978( .ZN(II37946), .A(g28529) );
  INV_X1 NOT_11979( .ZN(g28979), .A(II37946) );
  INV_X1 NOT_11980( .ZN(II37950), .A(g28556) );
  INV_X1 NOT_11981( .ZN(g28983), .A(II37950) );
  INV_X16 NOT_11982( .ZN(II37956), .A(g28584) );
  INV_X16 NOT_11983( .ZN(g28993), .A(II37956) );
  INV_X16 NOT_11984( .ZN(II37961), .A(g28501) );
  INV_X1 NOT_11985( .ZN(g28998), .A(II37961) );
  INV_X1 NOT_11986( .ZN(II37965), .A(g28529) );
  INV_X1 NOT_11987( .ZN(g29002), .A(II37965) );
  INV_X1 NOT_11988( .ZN(II37968), .A(g28529) );
  INV_X1 NOT_11989( .ZN(g29005), .A(II37968) );
  INV_X1 NOT_11990( .ZN(II37973), .A(g28556) );
  INV_X1 NOT_11991( .ZN(g29010), .A(II37973) );
  INV_X1 NOT_11992( .ZN(II37978), .A(g28584) );
  INV_X1 NOT_11993( .ZN(g29019), .A(II37978) );
  INV_X1 NOT_11994( .ZN(II37982), .A(g28501) );
  INV_X1 NOT_11995( .ZN(g29023), .A(II37982) );
  INV_X1 NOT_11996( .ZN(II37986), .A(g28529) );
  INV_X1 NOT_11997( .ZN(g29027), .A(II37986) );
  INV_X1 NOT_11998( .ZN(II37991), .A(g28556) );
  INV_X1 NOT_11999( .ZN(g29032), .A(II37991) );
  INV_X1 NOT_12000( .ZN(II37994), .A(g28556) );
  INV_X1 NOT_12001( .ZN(g29035), .A(II37994) );
  INV_X1 NOT_12002( .ZN(II37999), .A(g28584) );
  INV_X1 NOT_12003( .ZN(g29042), .A(II37999) );
  INV_X1 NOT_12004( .ZN(II38003), .A(g28529) );
  INV_X1 NOT_12005( .ZN(g29046), .A(II38003) );
  INV_X1 NOT_12006( .ZN(II38007), .A(g28556) );
  INV_X1 NOT_12007( .ZN(g29050), .A(II38007) );
  INV_X1 NOT_12008( .ZN(II38011), .A(g28584) );
  INV_X1 NOT_12009( .ZN(g29054), .A(II38011) );
  INV_X1 NOT_12010( .ZN(II38014), .A(g28584) );
  INV_X1 NOT_12011( .ZN(g29057), .A(II38014) );
  INV_X1 NOT_12012( .ZN(II38018), .A(g28342) );
  INV_X1 NOT_12013( .ZN(g29061), .A(II38018) );
  INV_X1 NOT_12014( .ZN(II38024), .A(g28556) );
  INV_X1 NOT_12015( .ZN(g29065), .A(II38024) );
  INV_X1 NOT_12016( .ZN(II38028), .A(g28584) );
  INV_X1 NOT_12017( .ZN(g29069), .A(II38028) );
  INV_X1 NOT_12018( .ZN(II38032), .A(g28344) );
  INV_X1 NOT_12019( .ZN(g29073), .A(II38032) );
  INV_X1 NOT_12020( .ZN(II38035), .A(g28345) );
  INV_X1 NOT_12021( .ZN(g29074), .A(II38035) );
  INV_X1 NOT_12022( .ZN(II38038), .A(g28346) );
  INV_X1 NOT_12023( .ZN(g29075), .A(II38038) );
  INV_X1 NOT_12024( .ZN(II38042), .A(g28584) );
  INV_X1 NOT_12025( .ZN(g29077), .A(II38042) );
  INV_X1 NOT_12026( .ZN(II38046), .A(g28348) );
  INV_X1 NOT_12027( .ZN(g29081), .A(II38046) );
  INV_X1 NOT_12028( .ZN(II38049), .A(g28349) );
  INV_X1 NOT_12029( .ZN(g29082), .A(II38049) );
  INV_X1 NOT_12030( .ZN(II38053), .A(g28350) );
  INV_X1 NOT_12031( .ZN(g29084), .A(II38053) );
  INV_X1 NOT_12032( .ZN(II38056), .A(g28351) );
  INV_X1 NOT_12033( .ZN(g29085), .A(II38056) );
  INV_X1 NOT_12034( .ZN(II38059), .A(g28352) );
  INV_X1 NOT_12035( .ZN(g29086), .A(II38059) );
  INV_X1 NOT_12036( .ZN(II38064), .A(g28353) );
  INV_X1 NOT_12037( .ZN(g29089), .A(II38064) );
  INV_X1 NOT_12038( .ZN(II38068), .A(g28354) );
  INV_X1 NOT_12039( .ZN(g29091), .A(II38068) );
  INV_X1 NOT_12040( .ZN(II38071), .A(g28355) );
  INV_X1 NOT_12041( .ZN(g29092), .A(II38071) );
  INV_X1 NOT_12042( .ZN(II38074), .A(g28356) );
  INV_X1 NOT_12043( .ZN(g29093), .A(II38074) );
  INV_X1 NOT_12044( .ZN(II38077), .A(g28357) );
  INV_X1 NOT_12045( .ZN(g29094), .A(II38077) );
  INV_X1 NOT_12046( .ZN(II38080), .A(g28358) );
  INV_X1 NOT_12047( .ZN(g29095), .A(II38080) );
  INV_X1 NOT_12048( .ZN(II38085), .A(g28360) );
  INV_X1 NOT_12049( .ZN(g29098), .A(II38085) );
  INV_X1 NOT_12050( .ZN(II38088), .A(g28361) );
  INV_X1 NOT_12051( .ZN(g29099), .A(II38088) );
  INV_X1 NOT_12052( .ZN(II38091), .A(g28362) );
  INV_X1 NOT_12053( .ZN(g29100), .A(II38091) );
  INV_X1 NOT_12054( .ZN(II38094), .A(g28363) );
  INV_X1 NOT_12055( .ZN(g29101), .A(II38094) );
  INV_X1 NOT_12056( .ZN(II38097), .A(g28364) );
  INV_X1 NOT_12057( .ZN(g29102), .A(II38097) );
  INV_X1 NOT_12058( .ZN(II38101), .A(g28366) );
  INV_X1 NOT_12059( .ZN(g29104), .A(II38101) );
  INV_X1 NOT_12060( .ZN(II38104), .A(g28367) );
  INV_X1 NOT_12061( .ZN(g29105), .A(II38104) );
  INV_X1 NOT_12062( .ZN(II38107), .A(g28368) );
  INV_X1 NOT_12063( .ZN(g29106), .A(II38107) );
  INV_X1 NOT_12064( .ZN(II38111), .A(g28371) );
  INV_X1 NOT_12065( .ZN(g29108), .A(II38111) );
  INV_X1 NOT_12066( .ZN(II38119), .A(g28420) );
  INV_X1 NOT_12067( .ZN(g29117), .A(II38119) );
  INV_X1 NOT_12068( .ZN(II38122), .A(g28421) );
  INV_X1 NOT_12069( .ZN(g29118), .A(II38122) );
  INV_X1 NOT_12070( .ZN(II38125), .A(g28425) );
  INV_X1 NOT_12071( .ZN(g29119), .A(II38125) );
  INV_X1 NOT_12072( .ZN(II38128), .A(g28419) );
  INV_X1 NOT_12073( .ZN(g29120), .A(II38128) );
  INV_X1 NOT_12074( .ZN(II38136), .A(g28833) );
  INV_X1 NOT_12075( .ZN(g29131), .A(II38136) );
  INV_X1 NOT_12076( .ZN(II38139), .A(g29061) );
  INV_X1 NOT_12077( .ZN(g29132), .A(II38139) );
  INV_X1 NOT_12078( .ZN(II38142), .A(g29073) );
  INV_X1 NOT_12079( .ZN(g29133), .A(II38142) );
  INV_X1 NOT_12080( .ZN(II38145), .A(g29081) );
  INV_X1 NOT_12081( .ZN(g29134), .A(II38145) );
  INV_X1 NOT_12082( .ZN(II38148), .A(g29074) );
  INV_X1 NOT_12083( .ZN(g29135), .A(II38148) );
  INV_X1 NOT_12084( .ZN(II38151), .A(g29082) );
  INV_X1 NOT_12085( .ZN(g29136), .A(II38151) );
  INV_X1 NOT_12086( .ZN(II38154), .A(g29089) );
  INV_X1 NOT_12087( .ZN(g29137), .A(II38154) );
  INV_X1 NOT_12088( .ZN(II38157), .A(g28882) );
  INV_X1 NOT_12089( .ZN(g29138), .A(II38157) );
  INV_X1 NOT_12090( .ZN(II38160), .A(g28835) );
  INV_X1 NOT_12091( .ZN(g29139), .A(II38160) );
  INV_X1 NOT_12092( .ZN(II38163), .A(g29075) );
  INV_X1 NOT_12093( .ZN(g29140), .A(II38163) );
  INV_X1 NOT_12094( .ZN(II38166), .A(g29084) );
  INV_X1 NOT_12095( .ZN(g29141), .A(II38166) );
  INV_X1 NOT_12096( .ZN(II38169), .A(g29091) );
  INV_X1 NOT_12097( .ZN(g29142), .A(II38169) );
  INV_X1 NOT_12098( .ZN(II38172), .A(g29085) );
  INV_X1 NOT_12099( .ZN(g29143), .A(II38172) );
  INV_X1 NOT_12100( .ZN(II38175), .A(g29092) );
  INV_X1 NOT_12101( .ZN(g29144), .A(II38175) );
  INV_X1 NOT_12102( .ZN(II38178), .A(g29098) );
  INV_X1 NOT_12103( .ZN(g29145), .A(II38178) );
  INV_X1 NOT_12104( .ZN(II38181), .A(g28899) );
  INV_X1 NOT_12105( .ZN(g29146), .A(II38181) );
  INV_X1 NOT_12106( .ZN(II38184), .A(g28837) );
  INV_X1 NOT_12107( .ZN(g29147), .A(II38184) );
  INV_X1 NOT_12108( .ZN(II38187), .A(g29086) );
  INV_X1 NOT_12109( .ZN(g29148), .A(II38187) );
  INV_X1 NOT_12110( .ZN(II38190), .A(g29093) );
  INV_X1 NOT_12111( .ZN(g29149), .A(II38190) );
  INV_X1 NOT_12112( .ZN(II38193), .A(g29099) );
  INV_X1 NOT_12113( .ZN(g29150), .A(II38193) );
  INV_X1 NOT_12114( .ZN(II38196), .A(g29094) );
  INV_X1 NOT_12115( .ZN(g29151), .A(II38196) );
  INV_X1 NOT_12116( .ZN(II38199), .A(g29100) );
  INV_X1 NOT_12117( .ZN(g29152), .A(II38199) );
  INV_X1 NOT_12118( .ZN(II38202), .A(g29104) );
  INV_X1 NOT_12119( .ZN(g29153), .A(II38202) );
  INV_X1 NOT_12120( .ZN(II38205), .A(g28924) );
  INV_X1 NOT_12121( .ZN(g29154), .A(II38205) );
  INV_X1 NOT_12122( .ZN(II38208), .A(g28839) );
  INV_X1 NOT_12123( .ZN(g29155), .A(II38208) );
  INV_X1 NOT_12124( .ZN(II38211), .A(g29095) );
  INV_X1 NOT_12125( .ZN(g29156), .A(II38211) );
  INV_X1 NOT_12126( .ZN(II38214), .A(g29101) );
  INV_X1 NOT_12127( .ZN(g29157), .A(II38214) );
  INV_X1 NOT_12128( .ZN(II38217), .A(g29105) );
  INV_X1 NOT_12129( .ZN(g29158), .A(II38217) );
  INV_X1 NOT_12130( .ZN(II38220), .A(g29102) );
  INV_X1 NOT_12131( .ZN(g29159), .A(II38220) );
  INV_X1 NOT_12132( .ZN(II38223), .A(g29106) );
  INV_X1 NOT_12133( .ZN(g29160), .A(II38223) );
  INV_X1 NOT_12134( .ZN(II38226), .A(g29108) );
  INV_X1 NOT_12135( .ZN(g29161), .A(II38226) );
  INV_X1 NOT_12136( .ZN(II38229), .A(g28950) );
  INV_X1 NOT_12137( .ZN(g29162), .A(II38229) );
  INV_X1 NOT_12138( .ZN(II38232), .A(g29117) );
  INV_X1 NOT_12139( .ZN(g29163), .A(II38232) );
  INV_X1 NOT_12140( .ZN(II38235), .A(g29118) );
  INV_X1 NOT_12141( .ZN(g29164), .A(II38235) );
  INV_X1 NOT_12142( .ZN(II38238), .A(g29119) );
  INV_X1 NOT_12143( .ZN(g29165), .A(II38238) );
  INV_X1 NOT_12144( .ZN(II38241), .A(g28832) );
  INV_X1 NOT_12145( .ZN(g29166), .A(II38241) );
  INV_X1 NOT_12146( .ZN(II38245), .A(g28920) );
  INV_X1 NOT_12147( .ZN(g29168), .A(II38245) );
  INV_X1 NOT_12148( .ZN(II38250), .A(g28941) );
  INV_X1 NOT_12149( .ZN(g29171), .A(II38250) );
  INV_X1 NOT_12150( .ZN(II38258), .A(g28963) );
  INV_X1 NOT_12151( .ZN(g29177), .A(II38258) );
  INV_X1 NOT_12152( .ZN(II38272), .A(g29013) );
  INV_X1 NOT_12153( .ZN(g29189), .A(II38272) );
  INV_X1 NOT_12154( .ZN(II38275), .A(g28987) );
  INV_X1 NOT_12155( .ZN(g29190), .A(II38275) );
  INV_X1 NOT_12156( .ZN(II38278), .A(g28963) );
  INV_X1 NOT_12157( .ZN(g29191), .A(II38278) );
  INV_X1 NOT_12158( .ZN(g29192), .A(g28954) );
  INV_X1 NOT_12159( .ZN(II38282), .A(g28941) );
  INV_X1 NOT_12160( .ZN(g29193), .A(II38282) );
  INV_X1 NOT_12161( .ZN(II38321), .A(g29113) );
  INV_X1 NOT_12162( .ZN(g29230), .A(II38321) );
  INV_X1 NOT_12163( .ZN(II38330), .A(g29120) );
  INV_X1 NOT_12164( .ZN(g29237), .A(II38330) );
  INV_X1 NOT_12165( .ZN(II38339), .A(g29120) );
  INV_X1 NOT_12166( .ZN(g29244), .A(II38339) );
  INV_X1 NOT_12167( .ZN(II38342), .A(g28886) );
  INV_X16 NOT_12168( .ZN(g29245), .A(II38342) );
  INV_X16 NOT_12169( .ZN(II38345), .A(g29109) );
  INV_X1 NOT_12170( .ZN(g29246), .A(II38345) );
  INV_X1 NOT_12171( .ZN(II38348), .A(g28874) );
  INV_X1 NOT_12172( .ZN(g29247), .A(II38348) );
  INV_X1 NOT_12173( .ZN(II38352), .A(g29110) );
  INV_X1 NOT_12174( .ZN(g29249), .A(II38352) );
  INV_X1 NOT_12175( .ZN(II38355), .A(g29039) );
  INV_X1 NOT_12176( .ZN(g29250), .A(II38355) );
  INV_X1 NOT_12177( .ZN(II38360), .A(g29111) );
  INV_X1 NOT_12178( .ZN(g29253), .A(II38360) );
  INV_X1 NOT_12179( .ZN(II38363), .A(g29016) );
  INV_X1 NOT_12180( .ZN(g29254), .A(II38363) );
  INV_X1 NOT_12181( .ZN(II38369), .A(g29112) );
  INV_X1 NOT_12182( .ZN(g29258), .A(II38369) );
  INV_X1 NOT_12183( .ZN(g29266), .A(g28741) );
  INV_X1 NOT_12184( .ZN(II38386), .A(g28734) );
  INV_X1 NOT_12185( .ZN(g29267), .A(II38386) );
  INV_X1 NOT_12186( .ZN(g29268), .A(g28751) );
  INV_X1 NOT_12187( .ZN(g29269), .A(g28755) );
  INV_X1 NOT_12188( .ZN(II38391), .A(g28730) );
  INV_X1 NOT_12189( .ZN(g29270), .A(II38391) );
  INV_X1 NOT_12190( .ZN(g29271), .A(g28764) );
  INV_X1 NOT_12191( .ZN(g29272), .A(g28768) );
  INV_X1 NOT_12192( .ZN(II38396), .A(g28727) );
  INV_X1 NOT_12193( .ZN(g29273), .A(II38396) );
  INV_X1 NOT_12194( .ZN(g29274), .A(g28775) );
  INV_X1 NOT_12195( .ZN(g29275), .A(g28779) );
  INV_X1 NOT_12196( .ZN(II38401), .A(g28725) );
  INV_X1 NOT_12197( .ZN(g29276), .A(II38401) );
  INV_X1 NOT_12198( .ZN(g29277), .A(g28785) );
  INV_X1 NOT_12199( .ZN(II38405), .A(g28723) );
  INV_X1 NOT_12200( .ZN(g29278), .A(II38405) );
  INV_X1 NOT_12201( .ZN(II38408), .A(g28721) );
  INV_X1 NOT_12202( .ZN(g29279), .A(II38408) );
  INV_X1 NOT_12203( .ZN(g29280), .A(g28791) );
  INV_X1 NOT_12204( .ZN(II38412), .A(g28720) );
  INV_X1 NOT_12205( .ZN(g29281), .A(II38412) );
  INV_X1 NOT_12206( .ZN(g29282), .A(g28796) );
  INV_X1 NOT_12207( .ZN(g29283), .A(g28799) );
  INV_X1 NOT_12208( .ZN(g29285), .A(g28804) );
  INV_X1 NOT_12209( .ZN(g29286), .A(g28807) );
  INV_X1 NOT_12210( .ZN(g29287), .A(g28810) );
  INV_X1 NOT_12211( .ZN(II38421), .A(g28740) );
  INV_X1 NOT_12212( .ZN(g29288), .A(II38421) );
  INV_X1 NOT_12213( .ZN(g29290), .A(g28814) );
  INV_X1 NOT_12214( .ZN(g29291), .A(g28817) );
  INV_X1 NOT_12215( .ZN(g29292), .A(g28820) );
  INV_X1 NOT_12216( .ZN(II38428), .A(g28732) );
  INV_X1 NOT_12217( .ZN(g29293), .A(II38428) );
  INV_X1 NOT_12218( .ZN(g29295), .A(g28823) );
  INV_X1 NOT_12219( .ZN(g29296), .A(g28826) );
  INV_X1 NOT_12220( .ZN(II38434), .A(g28735) );
  INV_X1 NOT_12221( .ZN(g29297), .A(II38434) );
  INV_X1 NOT_12222( .ZN(II38437), .A(g28736) );
  INV_X1 NOT_12223( .ZN(g29298), .A(II38437) );
  INV_X1 NOT_12224( .ZN(II38440), .A(g28738) );
  INV_X1 NOT_12225( .ZN(g29299), .A(II38440) );
  INV_X1 NOT_12226( .ZN(g29301), .A(g28829) );
  INV_X1 NOT_12227( .ZN(II38447), .A(g28744) );
  INV_X1 NOT_12228( .ZN(g29304), .A(II38447) );
  INV_X1 NOT_12229( .ZN(II38450), .A(g28745) );
  INV_X1 NOT_12230( .ZN(g29305), .A(II38450) );
  INV_X1 NOT_12231( .ZN(II38453), .A(g28746) );
  INV_X1 NOT_12232( .ZN(g29306), .A(II38453) );
  INV_X1 NOT_12233( .ZN(II38456), .A(g28747) );
  INV_X1 NOT_12234( .ZN(g29307), .A(II38456) );
  INV_X1 NOT_12235( .ZN(II38459), .A(g28749) );
  INV_X1 NOT_12236( .ZN(g29308), .A(II38459) );
  INV_X1 NOT_12237( .ZN(II38462), .A(g29120) );
  INV_X1 NOT_12238( .ZN(g29309), .A(II38462) );
  INV_X1 NOT_12239( .ZN(II38466), .A(g28754) );
  INV_X1 NOT_12240( .ZN(g29311), .A(II38466) );
  INV_X1 NOT_12241( .ZN(II38471), .A(g28758) );
  INV_X1 NOT_12242( .ZN(g29314), .A(II38471) );
  INV_X1 NOT_12243( .ZN(II38474), .A(g28759) );
  INV_X1 NOT_12244( .ZN(g29315), .A(II38474) );
  INV_X1 NOT_12245( .ZN(II38477), .A(g28760) );
  INV_X1 NOT_12246( .ZN(g29316), .A(II38477) );
  INV_X1 NOT_12247( .ZN(II38480), .A(g28761) );
  INV_X1 NOT_12248( .ZN(g29317), .A(II38480) );
  INV_X1 NOT_12249( .ZN(II38483), .A(g28990) );
  INV_X1 NOT_12250( .ZN(g29318), .A(II38483) );
  INV_X1 NOT_12251( .ZN(II38486), .A(g28763) );
  INV_X1 NOT_12252( .ZN(g29319), .A(II38486) );
  INV_X1 NOT_12253( .ZN(II38491), .A(g28767) );
  INV_X1 NOT_12254( .ZN(g29322), .A(II38491) );
  INV_X1 NOT_12255( .ZN(II38496), .A(g28771) );
  INV_X1 NOT_12256( .ZN(g29325), .A(II38496) );
  INV_X1 NOT_12257( .ZN(II38499), .A(g28772) );
  INV_X1 NOT_12258( .ZN(g29326), .A(II38499) );
  INV_X1 NOT_12259( .ZN(II38502), .A(g28773) );
  INV_X1 NOT_12260( .ZN(g29327), .A(II38502) );
  INV_X1 NOT_12261( .ZN(II38505), .A(g28774) );
  INV_X1 NOT_12262( .ZN(g29328), .A(II38505) );
  INV_X1 NOT_12263( .ZN(II38510), .A(g28778) );
  INV_X1 NOT_12264( .ZN(g29331), .A(II38510) );
  INV_X1 NOT_12265( .ZN(II38515), .A(g28782) );
  INV_X1 NOT_12266( .ZN(g29334), .A(II38515) );
  INV_X1 NOT_12267( .ZN(II38518), .A(g28783) );
  INV_X1 NOT_12268( .ZN(g29335), .A(II38518) );
  INV_X1 NOT_12269( .ZN(II38524), .A(g28788) );
  INV_X16 NOT_12270( .ZN(g29339), .A(II38524) );
  INV_X16 NOT_12271( .ZN(II38536), .A(g28920) );
  INV_X1 NOT_12272( .ZN(g29349), .A(II38536) );
  INV_X1 NOT_12273( .ZN(II38539), .A(g29113) );
  INV_X1 NOT_12274( .ZN(g29350), .A(II38539) );
  INV_X1 NOT_12275( .ZN(g29356), .A(g29120) );
  INV_X1 NOT_12276( .ZN(g29358), .A(g29120) );
  INV_X1 NOT_12277( .ZN(II38548), .A(g28903) );
  INV_X1 NOT_12278( .ZN(g29359), .A(II38548) );
  INV_X1 NOT_12279( .ZN(g29360), .A(g28871) );
  INV_X1 NOT_12280( .ZN(g29361), .A(g28877) );
  INV_X1 NOT_12281( .ZN(g29362), .A(g28883) );
  INV_X1 NOT_12282( .ZN(g29363), .A(g28889) );
  INV_X1 NOT_12283( .ZN(g29364), .A(g28894) );
  INV_X1 NOT_12284( .ZN(g29365), .A(g28900) );
  INV_X1 NOT_12285( .ZN(g29366), .A(g28906) );
  INV_X1 NOT_12286( .ZN(g29367), .A(g28911) );
  INV_X1 NOT_12287( .ZN(g29368), .A(g28916) );
  INV_X1 NOT_12288( .ZN(g29369), .A(g28925) );
  INV_X1 NOT_12289( .ZN(g29370), .A(g28928) );
  INV_X1 NOT_12290( .ZN(g29371), .A(g28932) );
  INV_X1 NOT_12291( .ZN(g29372), .A(g28937) );
  INV_X1 NOT_12292( .ZN(g29373), .A(g28945) );
  INV_X1 NOT_12293( .ZN(g29374), .A(g28951) );
  INV_X1 NOT_12294( .ZN(g29375), .A(g28955) );
  INV_X1 NOT_12295( .ZN(g29376), .A(g28959) );
  INV_X1 NOT_12296( .ZN(g29377), .A(g28967) );
  INV_X1 NOT_12297( .ZN(g29378), .A(g28972) );
  INV_X1 NOT_12298( .ZN(g29379), .A(g28975) );
  INV_X1 NOT_12299( .ZN(g29380), .A(g28979) );
  INV_X1 NOT_12300( .ZN(g29381), .A(g28983) );
  INV_X1 NOT_12301( .ZN(g29382), .A(g28993) );
  INV_X1 NOT_12302( .ZN(g29383), .A(g28998) );
  INV_X1 NOT_12303( .ZN(g29384), .A(g29002) );
  INV_X1 NOT_12304( .ZN(g29385), .A(g29005) );
  INV_X1 NOT_12305( .ZN(g29386), .A(g29010) );
  INV_X1 NOT_12306( .ZN(g29387), .A(g29019) );
  INV_X1 NOT_12307( .ZN(g29388), .A(g29023) );
  INV_X1 NOT_12308( .ZN(g29389), .A(g29027) );
  INV_X1 NOT_12309( .ZN(g29390), .A(g29032) );
  INV_X1 NOT_12310( .ZN(g29391), .A(g29035) );
  INV_X1 NOT_12311( .ZN(g29392), .A(g29042) );
  INV_X1 NOT_12312( .ZN(g29393), .A(g29046) );
  INV_X1 NOT_12313( .ZN(g29394), .A(g29050) );
  INV_X1 NOT_12314( .ZN(g29395), .A(g29054) );
  INV_X1 NOT_12315( .ZN(g29396), .A(g29057) );
  INV_X1 NOT_12316( .ZN(g29397), .A(g29065) );
  INV_X1 NOT_12317( .ZN(g29398), .A(g29069) );
  INV_X1 NOT_12318( .ZN(II38591), .A(g28987) );
  INV_X1 NOT_12319( .ZN(g29400), .A(II38591) );
  INV_X1 NOT_12320( .ZN(II38594), .A(g28990) );
  INV_X1 NOT_12321( .ZN(g29401), .A(II38594) );
  INV_X1 NOT_12322( .ZN(g29402), .A(g29077) );
  INV_X1 NOT_12323( .ZN(II38599), .A(g29013) );
  INV_X1 NOT_12324( .ZN(g29404), .A(II38599) );
  INV_X1 NOT_12325( .ZN(II38602), .A(g29016) );
  INV_X1 NOT_12326( .ZN(g29405), .A(II38602) );
  INV_X1 NOT_12327( .ZN(II38606), .A(g29039) );
  INV_X1 NOT_12328( .ZN(g29407), .A(II38606) );
  INV_X1 NOT_12329( .ZN(II38609), .A(g28874) );
  INV_X1 NOT_12330( .ZN(g29408), .A(II38609) );
  INV_X1 NOT_12331( .ZN(II38613), .A(g28886) );
  INV_X1 NOT_12332( .ZN(g29410), .A(II38613) );
  INV_X16 NOT_12333( .ZN(II38617), .A(g28903) );
  INV_X1 NOT_12334( .ZN(g29412), .A(II38617) );
  INV_X1 NOT_12335( .ZN(II38620), .A(g29246) );
  INV_X1 NOT_12336( .ZN(g29413), .A(II38620) );
  INV_X1 NOT_12337( .ZN(II38623), .A(g29293) );
  INV_X1 NOT_12338( .ZN(g29414), .A(II38623) );
  INV_X1 NOT_12339( .ZN(II38626), .A(g29297) );
  INV_X1 NOT_12340( .ZN(g29415), .A(II38626) );
  INV_X1 NOT_12341( .ZN(II38629), .A(g29304) );
  INV_X1 NOT_12342( .ZN(g29416), .A(II38629) );
  INV_X1 NOT_12343( .ZN(II38632), .A(g29298) );
  INV_X1 NOT_12344( .ZN(g29417), .A(II38632) );
  INV_X1 NOT_12345( .ZN(II38635), .A(g29305) );
  INV_X1 NOT_12346( .ZN(g29418), .A(II38635) );
  INV_X1 NOT_12347( .ZN(II38638), .A(g29311) );
  INV_X1 NOT_12348( .ZN(g29419), .A(II38638) );
  INV_X1 NOT_12349( .ZN(II38641), .A(g29249) );
  INV_X1 NOT_12350( .ZN(g29420), .A(II38641) );
  INV_X1 NOT_12351( .ZN(II38644), .A(g29299) );
  INV_X1 NOT_12352( .ZN(g29421), .A(II38644) );
  INV_X1 NOT_12353( .ZN(II38647), .A(g29306) );
  INV_X1 NOT_12354( .ZN(g29422), .A(II38647) );
  INV_X1 NOT_12355( .ZN(II38650), .A(g29314) );
  INV_X1 NOT_12356( .ZN(g29423), .A(II38650) );
  INV_X1 NOT_12357( .ZN(II38653), .A(g29307) );
  INV_X1 NOT_12358( .ZN(g29424), .A(II38653) );
  INV_X1 NOT_12359( .ZN(II38656), .A(g29315) );
  INV_X1 NOT_12360( .ZN(g29425), .A(II38656) );
  INV_X1 NOT_12361( .ZN(II38659), .A(g29322) );
  INV_X1 NOT_12362( .ZN(g29426), .A(II38659) );
  INV_X1 NOT_12363( .ZN(II38662), .A(g29253) );
  INV_X1 NOT_12364( .ZN(g29427), .A(II38662) );
  INV_X1 NOT_12365( .ZN(II38665), .A(g29412) );
  INV_X1 NOT_12366( .ZN(g29428), .A(II38665) );
  INV_X1 NOT_12367( .ZN(II38668), .A(g29168) );
  INV_X1 NOT_12368( .ZN(g29429), .A(II38668) );
  INV_X1 NOT_12369( .ZN(II38671), .A(g29171) );
  INV_X1 NOT_12370( .ZN(g29430), .A(II38671) );
  INV_X1 NOT_12371( .ZN(II38674), .A(g29177) );
  INV_X1 NOT_12372( .ZN(g29431), .A(II38674) );
  INV_X1 NOT_12373( .ZN(II38677), .A(g29400) );
  INV_X1 NOT_12374( .ZN(g29432), .A(II38677) );
  INV_X1 NOT_12375( .ZN(II38680), .A(g29404) );
  INV_X1 NOT_12376( .ZN(g29433), .A(II38680) );
  INV_X1 NOT_12377( .ZN(II38683), .A(g29308) );
  INV_X1 NOT_12378( .ZN(g29434), .A(II38683) );
  INV_X1 NOT_12379( .ZN(II38686), .A(g29316) );
  INV_X1 NOT_12380( .ZN(g29435), .A(II38686) );
  INV_X1 NOT_12381( .ZN(II38689), .A(g29325) );
  INV_X1 NOT_12382( .ZN(g29436), .A(II38689) );
  INV_X1 NOT_12383( .ZN(II38692), .A(g29317) );
  INV_X1 NOT_12384( .ZN(g29437), .A(II38692) );
  INV_X1 NOT_12385( .ZN(II38695), .A(g29326) );
  INV_X1 NOT_12386( .ZN(g29438), .A(II38695) );
  INV_X1 NOT_12387( .ZN(II38698), .A(g29331) );
  INV_X1 NOT_12388( .ZN(g29439), .A(II38698) );
  INV_X1 NOT_12389( .ZN(II38701), .A(g29401) );
  INV_X1 NOT_12390( .ZN(g29440), .A(II38701) );
  INV_X1 NOT_12391( .ZN(II38704), .A(g29405) );
  INV_X1 NOT_12392( .ZN(g29441), .A(II38704) );
  INV_X1 NOT_12393( .ZN(II38707), .A(g29407) );
  INV_X1 NOT_12394( .ZN(g29442), .A(II38707) );
  INV_X1 NOT_12395( .ZN(II38710), .A(g29408) );
  INV_X1 NOT_12396( .ZN(g29443), .A(II38710) );
  INV_X1 NOT_12397( .ZN(II38713), .A(g29410) );
  INV_X16 NOT_12398( .ZN(g29444), .A(II38713) );
  INV_X1 NOT_12399( .ZN(II38716), .A(g29230) );
  INV_X1 NOT_12400( .ZN(g29445), .A(II38716) );
  INV_X1 NOT_12401( .ZN(II38719), .A(g29258) );
  INV_X1 NOT_12402( .ZN(g29446), .A(II38719) );
  INV_X1 NOT_12403( .ZN(II38722), .A(g29319) );
  INV_X1 NOT_12404( .ZN(g29447), .A(II38722) );
  INV_X1 NOT_12405( .ZN(II38725), .A(g29327) );
  INV_X1 NOT_12406( .ZN(g29448), .A(II38725) );
  INV_X1 NOT_12407( .ZN(II38728), .A(g29334) );
  INV_X1 NOT_12408( .ZN(g29449), .A(II38728) );
  INV_X1 NOT_12409( .ZN(II38731), .A(g29328) );
  INV_X1 NOT_12410( .ZN(g29450), .A(II38731) );
  INV_X1 NOT_12411( .ZN(II38734), .A(g29335) );
  INV_X1 NOT_12412( .ZN(g29451), .A(II38734) );
  INV_X1 NOT_12413( .ZN(II38737), .A(g29339) );
  INV_X1 NOT_12414( .ZN(g29452), .A(II38737) );
  INV_X1 NOT_12415( .ZN(II38740), .A(g29288) );
  INV_X1 NOT_12416( .ZN(g29453), .A(II38740) );
  INV_X1 NOT_12417( .ZN(II38743), .A(g29267) );
  INV_X1 NOT_12418( .ZN(g29454), .A(II38743) );
  INV_X1 NOT_12419( .ZN(II38746), .A(g29270) );
  INV_X1 NOT_12420( .ZN(g29455), .A(II38746) );
  INV_X1 NOT_12421( .ZN(II38749), .A(g29273) );
  INV_X1 NOT_12422( .ZN(g29456), .A(II38749) );
  INV_X1 NOT_12423( .ZN(II38752), .A(g29276) );
  INV_X1 NOT_12424( .ZN(g29457), .A(II38752) );
  INV_X1 NOT_12425( .ZN(II38755), .A(g29278) );
  INV_X1 NOT_12426( .ZN(g29458), .A(II38755) );
  INV_X1 NOT_12427( .ZN(II38758), .A(g29279) );
  INV_X1 NOT_12428( .ZN(g29459), .A(II38758) );
  INV_X1 NOT_12429( .ZN(II38761), .A(g29281) );
  INV_X1 NOT_12430( .ZN(g29460), .A(II38761) );
  INV_X1 NOT_12431( .ZN(II38764), .A(g29237) );
  INV_X1 NOT_12432( .ZN(g29461), .A(II38764) );
  INV_X1 NOT_12433( .ZN(II38767), .A(g29244) );
  INV_X1 NOT_12434( .ZN(g29462), .A(II38767) );
  INV_X1 NOT_12435( .ZN(II38770), .A(g29309) );
  INV_X1 NOT_12436( .ZN(g29463), .A(II38770) );
  INV_X1 NOT_12437( .ZN(g29491), .A(g29350) );
  INV_X1 NOT_12438( .ZN(II38801), .A(g29358) );
  INV_X1 NOT_12439( .ZN(g29495), .A(II38801) );
  INV_X1 NOT_12440( .ZN(II38804), .A(g29353) );
  INV_X1 NOT_12441( .ZN(g29496), .A(II38804) );
  INV_X1 NOT_12442( .ZN(II38807), .A(g29356) );
  INV_X1 NOT_12443( .ZN(g29497), .A(II38807) );
  INV_X1 NOT_12444( .ZN(II38817), .A(g29354) );
  INV_X1 NOT_12445( .ZN(g29499), .A(II38817) );
  INV_X1 NOT_12446( .ZN(II38827), .A(g29355) );
  INV_X1 NOT_12447( .ZN(g29501), .A(II38827) );
  INV_X1 NOT_12448( .ZN(II38838), .A(g29357) );
  INV_X1 NOT_12449( .ZN(g29504), .A(II38838) );
  INV_X1 NOT_12450( .ZN(II38848), .A(g29167) );
  INV_X1 NOT_12451( .ZN(g29506), .A(II38848) );
  INV_X1 NOT_12452( .ZN(II38851), .A(g29169) );
  INV_X1 NOT_12453( .ZN(g29507), .A(II38851) );
  INV_X1 NOT_12454( .ZN(II38854), .A(g29170) );
  INV_X1 NOT_12455( .ZN(g29508), .A(II38854) );
  INV_X16 NOT_12456( .ZN(II38857), .A(g29172) );
  INV_X16 NOT_12457( .ZN(g29509), .A(II38857) );
  INV_X1 NOT_12458( .ZN(II38860), .A(g29173) );
  INV_X1 NOT_12459( .ZN(g29510), .A(II38860) );
  INV_X1 NOT_12460( .ZN(II38863), .A(g29178) );
  INV_X1 NOT_12461( .ZN(g29511), .A(II38863) );
  INV_X1 NOT_12462( .ZN(II38866), .A(g29179) );
  INV_X1 NOT_12463( .ZN(g29512), .A(II38866) );
  INV_X1 NOT_12464( .ZN(II38869), .A(g29181) );
  INV_X1 NOT_12465( .ZN(g29513), .A(II38869) );
  INV_X1 NOT_12466( .ZN(II38872), .A(g29182) );
  INV_X1 NOT_12467( .ZN(g29514), .A(II38872) );
  INV_X1 NOT_12468( .ZN(II38875), .A(g29184) );
  INV_X1 NOT_12469( .ZN(g29515), .A(II38875) );
  INV_X1 NOT_12470( .ZN(II38878), .A(g29185) );
  INV_X1 NOT_12471( .ZN(g29516), .A(II38878) );
  INV_X1 NOT_12472( .ZN(II38881), .A(g29187) );
  INV_X1 NOT_12473( .ZN(g29517), .A(II38881) );
  INV_X1 NOT_12474( .ZN(II38885), .A(g29192) );
  INV_X1 NOT_12475( .ZN(g29519), .A(II38885) );
  INV_X1 NOT_12476( .ZN(II38898), .A(g29194) );
  INV_X1 NOT_12477( .ZN(g29530), .A(II38898) );
  INV_X1 NOT_12478( .ZN(II38905), .A(g29197) );
  INV_X1 NOT_12479( .ZN(g29535), .A(II38905) );
  INV_X1 NOT_12480( .ZN(II38909), .A(g29198) );
  INV_X1 NOT_12481( .ZN(g29537), .A(II38909) );
  INV_X1 NOT_12482( .ZN(II38916), .A(g29201) );
  INV_X1 NOT_12483( .ZN(g29542), .A(II38916) );
  INV_X1 NOT_12484( .ZN(II38920), .A(g29204) );
  INV_X1 NOT_12485( .ZN(g29544), .A(II38920) );
  INV_X1 NOT_12486( .ZN(II38924), .A(g29205) );
  INV_X1 NOT_12487( .ZN(g29546), .A(II38924) );
  INV_X1 NOT_12488( .ZN(II38931), .A(g29209) );
  INV_X1 NOT_12489( .ZN(g29551), .A(II38931) );
  INV_X1 NOT_12490( .ZN(II38936), .A(g29212) );
  INV_X1 NOT_12491( .ZN(g29554), .A(II38936) );
  INV_X1 NOT_12492( .ZN(II38940), .A(g29213) );
  INV_X1 NOT_12493( .ZN(g29556), .A(II38940) );
  INV_X1 NOT_12494( .ZN(II38947), .A(g29218) );
  INV_X1 NOT_12495( .ZN(g29561), .A(II38947) );
  INV_X1 NOT_12496( .ZN(II38951), .A(g29221) );
  INV_X1 NOT_12497( .ZN(g29563), .A(II38951) );
  INV_X1 NOT_12498( .ZN(II38958), .A(g29226) );
  INV_X1 NOT_12499( .ZN(g29568), .A(II38958) );
  INV_X1 NOT_12500( .ZN(II38975), .A(g29348) );
  INV_X1 NOT_12501( .ZN(g29583), .A(II38975) );
  INV_X1 NOT_12502( .ZN(II38999), .A(g29496) );
  INV_X1 NOT_12503( .ZN(g29627), .A(II38999) );
  INV_X1 NOT_12504( .ZN(II39002), .A(g29506) );
  INV_X1 NOT_12505( .ZN(g29628), .A(II39002) );
  INV_X1 NOT_12506( .ZN(II39005), .A(g29507) );
  INV_X1 NOT_12507( .ZN(g29629), .A(II39005) );
  INV_X1 NOT_12508( .ZN(II39008), .A(g29509) );
  INV_X1 NOT_12509( .ZN(g29630), .A(II39008) );
  INV_X1 NOT_12510( .ZN(II39011), .A(g29530) );
  INV_X1 NOT_12511( .ZN(g29631), .A(II39011) );
  INV_X1 NOT_12512( .ZN(II39014), .A(g29535) );
  INV_X1 NOT_12513( .ZN(g29632), .A(II39014) );
  INV_X1 NOT_12514( .ZN(II39017), .A(g29542) );
  INV_X1 NOT_12515( .ZN(g29633), .A(II39017) );
  INV_X1 NOT_12516( .ZN(II39020), .A(g29499) );
  INV_X1 NOT_12517( .ZN(g29634), .A(II39020) );
  INV_X1 NOT_12518( .ZN(II39023), .A(g29508) );
  INV_X1 NOT_12519( .ZN(g29635), .A(II39023) );
  INV_X1 NOT_12520( .ZN(II39026), .A(g29510) );
  INV_X1 NOT_12521( .ZN(g29636), .A(II39026) );
  INV_X1 NOT_12522( .ZN(II39029), .A(g29512) );
  INV_X1 NOT_12523( .ZN(g29637), .A(II39029) );
  INV_X1 NOT_12524( .ZN(II39032), .A(g29537) );
  INV_X1 NOT_12525( .ZN(g29638), .A(II39032) );
  INV_X1 NOT_12526( .ZN(II39035), .A(g29544) );
  INV_X1 NOT_12527( .ZN(g29639), .A(II39035) );
  INV_X1 NOT_12528( .ZN(II39038), .A(g29551) );
  INV_X1 NOT_12529( .ZN(g29640), .A(II39038) );
  INV_X1 NOT_12530( .ZN(II39041), .A(g29501) );
  INV_X1 NOT_12531( .ZN(g29641), .A(II39041) );
  INV_X1 NOT_12532( .ZN(II39044), .A(g29511) );
  INV_X1 NOT_12533( .ZN(g29642), .A(II39044) );
  INV_X1 NOT_12534( .ZN(II39047), .A(g29513) );
  INV_X1 NOT_12535( .ZN(g29643), .A(II39047) );
  INV_X1 NOT_12536( .ZN(II39050), .A(g29515) );
  INV_X1 NOT_12537( .ZN(g29644), .A(II39050) );
  INV_X1 NOT_12538( .ZN(II39053), .A(g29546) );
  INV_X1 NOT_12539( .ZN(g29645), .A(II39053) );
  INV_X1 NOT_12540( .ZN(II39056), .A(g29554) );
  INV_X1 NOT_12541( .ZN(g29646), .A(II39056) );
  INV_X1 NOT_12542( .ZN(II39059), .A(g29561) );
  INV_X1 NOT_12543( .ZN(g29647), .A(II39059) );
  INV_X1 NOT_12544( .ZN(II39062), .A(g29504) );
  INV_X1 NOT_12545( .ZN(g29648), .A(II39062) );
  INV_X1 NOT_12546( .ZN(II39065), .A(g29514) );
  INV_X1 NOT_12547( .ZN(g29649), .A(II39065) );
  INV_X1 NOT_12548( .ZN(II39068), .A(g29516) );
  INV_X1 NOT_12549( .ZN(g29650), .A(II39068) );
  INV_X1 NOT_12550( .ZN(II39071), .A(g29517) );
  INV_X1 NOT_12551( .ZN(g29651), .A(II39071) );
  INV_X1 NOT_12552( .ZN(II39074), .A(g29556) );
  INV_X1 NOT_12553( .ZN(g29652), .A(II39074) );
  INV_X1 NOT_12554( .ZN(II39077), .A(g29563) );
  INV_X1 NOT_12555( .ZN(g29653), .A(II39077) );
  INV_X1 NOT_12556( .ZN(II39080), .A(g29568) );
  INV_X1 NOT_12557( .ZN(g29654), .A(II39080) );
  INV_X1 NOT_12558( .ZN(II39083), .A(g29519) );
  INV_X1 NOT_12559( .ZN(g29655), .A(II39083) );
  INV_X1 NOT_12560( .ZN(II39086), .A(g29497) );
  INV_X1 NOT_12561( .ZN(g29656), .A(II39086) );
  INV_X1 NOT_12562( .ZN(II39089), .A(g29495) );
  INV_X1 NOT_12563( .ZN(g29657), .A(II39089) );
  INV_X1 NOT_12564( .ZN(g29658), .A(g29574) );
  INV_X1 NOT_12565( .ZN(g29659), .A(g29571) );
  INV_X1 NOT_12566( .ZN(g29660), .A(g29578) );
  INV_X1 NOT_12567( .ZN(g29661), .A(g29576) );
  INV_X1 NOT_12568( .ZN(g29662), .A(g29570) );
  INV_X1 NOT_12569( .ZN(g29664), .A(g29552) );
  INV_X1 NOT_12570( .ZN(g29666), .A(g29577) );
  INV_X1 NOT_12571( .ZN(g29668), .A(g29569) );
  INV_X1 NOT_12572( .ZN(g29673), .A(g29583) );
  INV_X1 NOT_12573( .ZN(II39121), .A(g29579) );
  INV_X1 NOT_12574( .ZN(g29689), .A(II39121) );
  INV_X1 NOT_12575( .ZN(II39124), .A(g29606) );
  INV_X1 NOT_12576( .ZN(g29690), .A(II39124) );
  INV_X1 NOT_12577( .ZN(II39127), .A(g29608) );
  INV_X1 NOT_12578( .ZN(g29691), .A(II39127) );
  INV_X1 NOT_12579( .ZN(II39130), .A(g29580) );
  INV_X1 NOT_12580( .ZN(g29692), .A(II39130) );
  INV_X1 NOT_12581( .ZN(II39133), .A(g29609) );
  INV_X1 NOT_12582( .ZN(g29693), .A(II39133) );
  INV_X1 NOT_12583( .ZN(II39136), .A(g29611) );
  INV_X1 NOT_12584( .ZN(g29694), .A(II39136) );
  INV_X1 NOT_12585( .ZN(II39139), .A(g29612) );
  INV_X1 NOT_12586( .ZN(g29695), .A(II39139) );
  INV_X1 NOT_12587( .ZN(II39142), .A(g29581) );
  INV_X1 NOT_12588( .ZN(g29696), .A(II39142) );
  INV_X1 NOT_12589( .ZN(II39145), .A(g29613) );
  INV_X1 NOT_12590( .ZN(g29697), .A(II39145) );
  INV_X1 NOT_12591( .ZN(II39148), .A(g29616) );
  INV_X1 NOT_12592( .ZN(g29698), .A(II39148) );
  INV_X1 NOT_12593( .ZN(II39151), .A(g29617) );
  INV_X1 NOT_12594( .ZN(g29699), .A(II39151) );
  INV_X1 NOT_12595( .ZN(II39154), .A(g29582) );
  INV_X1 NOT_12596( .ZN(g29700), .A(II39154) );
  INV_X1 NOT_12597( .ZN(II39157), .A(g29618) );
  INV_X1 NOT_12598( .ZN(g29701), .A(II39157) );
  INV_X1 NOT_12599( .ZN(II39160), .A(g29620) );
  INV_X1 NOT_12600( .ZN(g29702), .A(II39160) );
  INV_X1 NOT_12601( .ZN(II39164), .A(g29621) );
  INV_X1 NOT_12602( .ZN(g29704), .A(II39164) );
  INV_X1 NOT_12603( .ZN(II39168), .A(g29623) );
  INV_X1 NOT_12604( .ZN(g29708), .A(II39168) );
  INV_X1 NOT_12605( .ZN(g29716), .A(g29498) );
  INV_X1 NOT_12606( .ZN(g29724), .A(g29500) );
  INV_X1 NOT_12607( .ZN(g29726), .A(g29503) );
  INV_X1 NOT_12608( .ZN(g29739), .A(g29505) );
  INV_X1 NOT_12609( .ZN(II39234), .A(g29689) );
  INV_X1 NOT_12610( .ZN(g29794), .A(II39234) );
  INV_X1 NOT_12611( .ZN(II39237), .A(g29690) );
  INV_X1 NOT_12612( .ZN(g29795), .A(II39237) );
  INV_X1 NOT_12613( .ZN(II39240), .A(g29691) );
  INV_X1 NOT_12614( .ZN(g29796), .A(II39240) );
  INV_X1 NOT_12615( .ZN(II39243), .A(g29694) );
  INV_X1 NOT_12616( .ZN(g29797), .A(II39243) );
  INV_X1 NOT_12617( .ZN(II39246), .A(g29692) );
  INV_X1 NOT_12618( .ZN(g29798), .A(II39246) );
  INV_X1 NOT_12619( .ZN(II39249), .A(g29693) );
  INV_X1 NOT_12620( .ZN(g29799), .A(II39249) );
  INV_X1 NOT_12621( .ZN(II39252), .A(g29695) );
  INV_X1 NOT_12622( .ZN(g29800), .A(II39252) );
  INV_X1 NOT_12623( .ZN(II39255), .A(g29698) );
  INV_X1 NOT_12624( .ZN(g29801), .A(II39255) );
  INV_X1 NOT_12625( .ZN(II39258), .A(g29696) );
  INV_X1 NOT_12626( .ZN(g29802), .A(II39258) );
  INV_X1 NOT_12627( .ZN(II39261), .A(g29697) );
  INV_X1 NOT_12628( .ZN(g29803), .A(II39261) );
  INV_X1 NOT_12629( .ZN(II39264), .A(g29699) );
  INV_X1 NOT_12630( .ZN(g29804), .A(II39264) );
  INV_X1 NOT_12631( .ZN(II39267), .A(g29702) );
  INV_X16 NOT_12632( .ZN(g29805), .A(II39267) );
  INV_X16 NOT_12633( .ZN(II39270), .A(g29700) );
  INV_X16 NOT_12634( .ZN(g29806), .A(II39270) );
  INV_X16 NOT_12635( .ZN(II39273), .A(g29701) );
  INV_X1 NOT_12636( .ZN(g29807), .A(II39273) );
  INV_X1 NOT_12637( .ZN(II39276), .A(g29704) );
  INV_X1 NOT_12638( .ZN(g29808), .A(II39276) );
  INV_X1 NOT_12639( .ZN(II39279), .A(g29708) );
  INV_X1 NOT_12640( .ZN(g29809), .A(II39279) );
  INV_X1 NOT_12641( .ZN(g29823), .A(g29663) );
  INV_X1 NOT_12642( .ZN(g29829), .A(g29665) );
  INV_X1 NOT_12643( .ZN(g29835), .A(g29667) );
  INV_X1 NOT_12644( .ZN(g29840), .A(g29669) );
  INV_X1 NOT_12645( .ZN(g29844), .A(g29670) );
  INV_X1 NOT_12646( .ZN(g29848), .A(g29761) );
  INV_X1 NOT_12647( .ZN(g29849), .A(g29671) );
  INV_X1 NOT_12648( .ZN(g29853), .A(g29672) );
  INV_X1 NOT_12649( .ZN(g29857), .A(g29676) );
  INV_X1 NOT_12650( .ZN(g29861), .A(g29677) );
  INV_X1 NOT_12651( .ZN(g29865), .A(g29678) );
  INV_X1 NOT_12652( .ZN(g29869), .A(g29679) );
  INV_X1 NOT_12653( .ZN(g29873), .A(g29680) );
  INV_X1 NOT_12654( .ZN(g29877), .A(g29681) );
  INV_X1 NOT_12655( .ZN(g29881), .A(g29682) );
  INV_X1 NOT_12656( .ZN(g29885), .A(g29683) );
  INV_X1 NOT_12657( .ZN(g29889), .A(g29684) );
  INV_X1 NOT_12658( .ZN(g29893), .A(g29685) );
  INV_X1 NOT_12659( .ZN(g29897), .A(g29686) );
  INV_X1 NOT_12660( .ZN(g29901), .A(g29687) );
  INV_X1 NOT_12661( .ZN(g29905), .A(g29688) );
  INV_X1 NOT_12662( .ZN(II39398), .A(g29664) );
  INV_X1 NOT_12663( .ZN(g29932), .A(II39398) );
  INV_X1 NOT_12664( .ZN(II39401), .A(g29662) );
  INV_X1 NOT_12665( .ZN(g29933), .A(II39401) );
  INV_X1 NOT_12666( .ZN(II39404), .A(g29661) );
  INV_X1 NOT_12667( .ZN(g29934), .A(II39404) );
  INV_X1 NOT_12668( .ZN(II39407), .A(g29660) );
  INV_X1 NOT_12669( .ZN(g29935), .A(II39407) );
  INV_X1 NOT_12670( .ZN(II39411), .A(g29659) );
  INV_X1 NOT_12671( .ZN(g29937), .A(II39411) );
  INV_X1 NOT_12672( .ZN(II39414), .A(g29658) );
  INV_X1 NOT_12673( .ZN(g29938), .A(II39414) );
  INV_X1 NOT_12674( .ZN(II39418), .A(g29668) );
  INV_X1 NOT_12675( .ZN(g29940), .A(II39418) );
  INV_X1 NOT_12676( .ZN(II39423), .A(g29666) );
  INV_X1 NOT_12677( .ZN(g29943), .A(II39423) );
  INV_X1 NOT_12678( .ZN(II39454), .A(g29940) );
  INV_X1 NOT_12679( .ZN(g29972), .A(II39454) );
  INV_X1 NOT_12680( .ZN(II39457), .A(g29943) );
  INV_X1 NOT_12681( .ZN(g29973), .A(II39457) );
  INV_X1 NOT_12682( .ZN(II39460), .A(g29932) );
  INV_X1 NOT_12683( .ZN(g29974), .A(II39460) );
  INV_X1 NOT_12684( .ZN(II39463), .A(g29933) );
  INV_X1 NOT_12685( .ZN(g29975), .A(II39463) );
  INV_X1 NOT_12686( .ZN(II39466), .A(g29934) );
  INV_X1 NOT_12687( .ZN(g29976), .A(II39466) );
  INV_X1 NOT_12688( .ZN(II39469), .A(g29935) );
  INV_X1 NOT_12689( .ZN(g29977), .A(II39469) );
  INV_X1 NOT_12690( .ZN(II39472), .A(g29937) );
  INV_X1 NOT_12691( .ZN(g29978), .A(II39472) );
  INV_X1 NOT_12692( .ZN(II39475), .A(g29938) );
  INV_X1 NOT_12693( .ZN(g29979), .A(II39475) );
  INV_X1 NOT_12694( .ZN(g30036), .A(g29912) );
  INV_X1 NOT_12695( .ZN(g30040), .A(g29914) );
  INV_X1 NOT_12696( .ZN(g30044), .A(g29916) );
  INV_X1 NOT_12697( .ZN(g30048), .A(g29920) );
  INV_X1 NOT_12698( .ZN(II39550), .A(g29848) );
  INV_X1 NOT_12699( .ZN(g30052), .A(II39550) );
  INV_X1 NOT_12700( .ZN(II39573), .A(g29936) );
  INV_X1 NOT_12701( .ZN(g30076), .A(II39573) );
  INV_X1 NOT_12702( .ZN(II39577), .A(g29939) );
  INV_X1 NOT_12703( .ZN(g30078), .A(II39577) );
  INV_X1 NOT_12704( .ZN(II39585), .A(g29941) );
  INV_X1 NOT_12705( .ZN(g30084), .A(II39585) );
  INV_X1 NOT_12706( .ZN(II39622), .A(g30052) );
  INV_X1 NOT_12707( .ZN(g30119), .A(II39622) );
  INV_X1 NOT_12708( .ZN(II39625), .A(g30076) );
  INV_X1 NOT_12709( .ZN(g30120), .A(II39625) );
  INV_X1 NOT_12710( .ZN(II39628), .A(g30078) );
  INV_X1 NOT_12711( .ZN(g30121), .A(II39628) );
  INV_X1 NOT_12712( .ZN(II39631), .A(g30084) );
  INV_X1 NOT_12713( .ZN(g30122), .A(II39631) );
  INV_X1 NOT_12714( .ZN(II39635), .A(g30055) );
  INV_X1 NOT_12715( .ZN(g30124), .A(II39635) );
  INV_X1 NOT_12716( .ZN(II39638), .A(g30056) );
  INV_X1 NOT_12717( .ZN(g30125), .A(II39638) );
  INV_X1 NOT_12718( .ZN(II39641), .A(g30057) );
  INV_X1 NOT_12719( .ZN(g30126), .A(II39641) );
  INV_X1 NOT_12720( .ZN(II39647), .A(g30058) );
  INV_X1 NOT_12721( .ZN(g30130), .A(II39647) );
  INV_X1 NOT_12722( .ZN(g30134), .A(g30010) );
  INV_X1 NOT_12723( .ZN(g30139), .A(g30011) );
  INV_X1 NOT_12724( .ZN(g30143), .A(g30012) );
  INV_X1 NOT_12725( .ZN(g30147), .A(g30013) );
  INV_X1 NOT_12726( .ZN(g30151), .A(g30014) );
  INV_X1 NOT_12727( .ZN(g30155), .A(g30015) );
  INV_X1 NOT_12728( .ZN(g30159), .A(g30016) );
  INV_X1 NOT_12729( .ZN(g30163), .A(g30017) );
  INV_X1 NOT_12730( .ZN(g30167), .A(g30018) );
  INV_X1 NOT_12731( .ZN(g30171), .A(g30019) );
  INV_X1 NOT_12732( .ZN(g30175), .A(g30020) );
  INV_X1 NOT_12733( .ZN(g30179), .A(g30021) );
  INV_X1 NOT_12734( .ZN(g30183), .A(g30022) );
  INV_X1 NOT_12735( .ZN(g30187), .A(g30023) );
  INV_X1 NOT_12736( .ZN(g30191), .A(g30024) );
  INV_X1 NOT_12737( .ZN(g30195), .A(g30025) );
  INV_X1 NOT_12738( .ZN(g30199), .A(g30026) );
  INV_X1 NOT_12739( .ZN(g30203), .A(g30027) );
  INV_X1 NOT_12740( .ZN(g30207), .A(g30028) );
  INV_X1 NOT_12741( .ZN(g30211), .A(g30029) );
  INV_X1 NOT_12742( .ZN(II39674), .A(g30072) );
  INV_X1 NOT_12743( .ZN(g30215), .A(II39674) );
  INV_X1 NOT_12744( .ZN(g30229), .A(g30030) );
  INV_X1 NOT_12745( .ZN(g30233), .A(g30031) );
  INV_X1 NOT_12746( .ZN(g30237), .A(g30032) );
  INV_X1 NOT_12747( .ZN(g30241), .A(g30033) );
  INV_X1 NOT_12748( .ZN(II39761), .A(g30072) );
  INV_X1 NOT_12749( .ZN(g30306), .A(II39761) );
  INV_X1 NOT_12750( .ZN(II39764), .A(g30060) );
  INV_X1 NOT_12751( .ZN(g30307), .A(II39764) );
  INV_X1 NOT_12752( .ZN(II39767), .A(g30061) );
  INV_X1 NOT_12753( .ZN(g30308), .A(II39767) );
  INV_X1 NOT_12754( .ZN(II39770), .A(g30063) );
  INV_X1 NOT_12755( .ZN(g30309), .A(II39770) );
  INV_X1 NOT_12756( .ZN(II39773), .A(g30064) );
  INV_X1 NOT_12757( .ZN(g30310), .A(II39773) );
  INV_X1 NOT_12758( .ZN(II39776), .A(g30066) );
  INV_X1 NOT_12759( .ZN(g30311), .A(II39776) );
  INV_X1 NOT_12760( .ZN(II39779), .A(g30053) );
  INV_X1 NOT_12761( .ZN(g30312), .A(II39779) );
  INV_X1 NOT_12762( .ZN(II39782), .A(g30054) );
  INV_X1 NOT_12763( .ZN(g30313), .A(II39782) );
  INV_X1 NOT_12764( .ZN(II39785), .A(g30124) );
  INV_X1 NOT_12765( .ZN(g30314), .A(II39785) );
  INV_X1 NOT_12766( .ZN(II39788), .A(g30125) );
  INV_X1 NOT_12767( .ZN(g30315), .A(II39788) );
  INV_X1 NOT_12768( .ZN(II39791), .A(g30126) );
  INV_X1 NOT_12769( .ZN(g30316), .A(II39791) );
  INV_X1 NOT_12770( .ZN(II39794), .A(g30130) );
  INV_X1 NOT_12771( .ZN(g30317), .A(II39794) );
  INV_X1 NOT_12772( .ZN(II39797), .A(g30307) );
  INV_X1 NOT_12773( .ZN(g30318), .A(II39797) );
  INV_X1 NOT_12774( .ZN(II39800), .A(g30309) );
  INV_X1 NOT_12775( .ZN(g30319), .A(II39800) );
  INV_X1 NOT_12776( .ZN(II39803), .A(g30308) );
  INV_X1 NOT_12777( .ZN(g30320), .A(II39803) );
  INV_X1 NOT_12778( .ZN(II39806), .A(g30310) );
  INV_X1 NOT_12779( .ZN(g30321), .A(II39806) );
  INV_X1 NOT_12780( .ZN(II39809), .A(g30311) );
  INV_X1 NOT_12781( .ZN(g30322), .A(II39809) );
  INV_X1 NOT_12782( .ZN(II39812), .A(g30312) );
  INV_X1 NOT_12783( .ZN(g30323), .A(II39812) );
  INV_X1 NOT_12784( .ZN(II39815), .A(g30313) );
  INV_X1 NOT_12785( .ZN(g30324), .A(II39815) );
  INV_X1 NOT_12786( .ZN(II39818), .A(g30215) );
  INV_X1 NOT_12787( .ZN(g30325), .A(II39818) );
  INV_X1 NOT_12788( .ZN(II39821), .A(g30267) );
  INV_X1 NOT_12789( .ZN(g30326), .A(II39821) );
  INV_X1 NOT_12790( .ZN(II39825), .A(g30268) );
  INV_X1 NOT_12791( .ZN(g30328), .A(II39825) );
  INV_X1 NOT_12792( .ZN(II39828), .A(g30269) );
  INV_X1 NOT_12793( .ZN(g30329), .A(II39828) );
  INV_X1 NOT_12794( .ZN(II39832), .A(g30270) );
  INV_X1 NOT_12795( .ZN(g30331), .A(II39832) );
  INV_X1 NOT_12796( .ZN(II39835), .A(g30271) );
  INV_X1 NOT_12797( .ZN(g30332), .A(II39835) );
  INV_X1 NOT_12798( .ZN(II39840), .A(g30272) );
  INV_X1 NOT_12799( .ZN(g30335), .A(II39840) );
  INV_X1 NOT_12800( .ZN(II39843), .A(g30273) );
  INV_X1 NOT_12801( .ZN(g30336), .A(II39843) );
  INV_X1 NOT_12802( .ZN(II39848), .A(g30274) );
  INV_X1 NOT_12803( .ZN(g30339), .A(II39848) );
  INV_X1 NOT_12804( .ZN(II39853), .A(g30275) );
  INV_X1 NOT_12805( .ZN(g30342), .A(II39853) );
  INV_X1 NOT_12806( .ZN(II39856), .A(g30276) );
  INV_X1 NOT_12807( .ZN(g30343), .A(II39856) );
  INV_X1 NOT_12808( .ZN(II39859), .A(g30277) );
  INV_X1 NOT_12809( .ZN(g30344), .A(II39859) );
  INV_X1 NOT_12810( .ZN(II39863), .A(g30278) );
  INV_X1 NOT_12811( .ZN(g30346), .A(II39863) );
  INV_X1 NOT_12812( .ZN(II39866), .A(g30279) );
  INV_X1 NOT_12813( .ZN(g30347), .A(II39866) );
  INV_X1 NOT_12814( .ZN(II39870), .A(g30280) );
  INV_X1 NOT_12815( .ZN(g30349), .A(II39870) );
  INV_X1 NOT_12816( .ZN(II39873), .A(g30281) );
  INV_X1 NOT_12817( .ZN(g30350), .A(II39873) );
  INV_X1 NOT_12818( .ZN(II39878), .A(g30282) );
  INV_X1 NOT_12819( .ZN(g30353), .A(II39878) );
  INV_X1 NOT_12820( .ZN(II39881), .A(g30283) );
  INV_X1 NOT_12821( .ZN(g30354), .A(II39881) );
  INV_X1 NOT_12822( .ZN(II39886), .A(g30284) );
  INV_X1 NOT_12823( .ZN(g30357), .A(II39886) );
  INV_X1 NOT_12824( .ZN(II39889), .A(g30285) );
  INV_X1 NOT_12825( .ZN(g30358), .A(II39889) );
  INV_X1 NOT_12826( .ZN(II39892), .A(g30286) );
  INV_X1 NOT_12827( .ZN(g30359), .A(II39892) );
  INV_X1 NOT_12828( .ZN(II39895), .A(g30287) );
  INV_X1 NOT_12829( .ZN(g30360), .A(II39895) );
  INV_X1 NOT_12830( .ZN(II39899), .A(g30288) );
  INV_X1 NOT_12831( .ZN(g30362), .A(II39899) );
  INV_X1 NOT_12832( .ZN(II39902), .A(g30289) );
  INV_X1 NOT_12833( .ZN(g30363), .A(II39902) );
  INV_X1 NOT_12834( .ZN(II39906), .A(g30290) );
  INV_X1 NOT_12835( .ZN(g30365), .A(II39906) );
  INV_X1 NOT_12836( .ZN(II39909), .A(g30291) );
  INV_X32 NOT_12837( .ZN(g30366), .A(II39909) );
  INV_X32 NOT_12838( .ZN(II39913), .A(g30292) );
  INV_X32 NOT_12839( .ZN(g30368), .A(II39913) );
  INV_X32 NOT_12840( .ZN(II39916), .A(g30293) );
  INV_X32 NOT_12841( .ZN(g30369), .A(II39916) );
  INV_X32 NOT_12842( .ZN(II39919), .A(g30294) );
  INV_X1 NOT_12843( .ZN(g30370), .A(II39919) );
  INV_X1 NOT_12844( .ZN(II39922), .A(g30295) );
  INV_X1 NOT_12845( .ZN(g30371), .A(II39922) );
  INV_X1 NOT_12846( .ZN(II39926), .A(g30296) );
  INV_X1 NOT_12847( .ZN(g30373), .A(II39926) );
  INV_X1 NOT_12848( .ZN(II39930), .A(g30297) );
  INV_X1 NOT_12849( .ZN(g30375), .A(II39930) );
  INV_X1 NOT_12850( .ZN(II39933), .A(g30298) );
  INV_X1 NOT_12851( .ZN(g30376), .A(II39933) );
  INV_X1 NOT_12852( .ZN(II39936), .A(g30299) );
  INV_X1 NOT_12853( .ZN(g30377), .A(II39936) );
  INV_X1 NOT_12854( .ZN(II39939), .A(g30300) );
  INV_X1 NOT_12855( .ZN(g30378), .A(II39939) );
  INV_X1 NOT_12856( .ZN(II39942), .A(g30301) );
  INV_X1 NOT_12857( .ZN(g30379), .A(II39942) );
  INV_X1 NOT_12858( .ZN(II39945), .A(g30302) );
  INV_X1 NOT_12859( .ZN(g30380), .A(II39945) );
  INV_X1 NOT_12860( .ZN(II39948), .A(g30303) );
  INV_X1 NOT_12861( .ZN(g30381), .A(II39948) );
  INV_X1 NOT_12862( .ZN(II39951), .A(g30304) );
  INV_X1 NOT_12863( .ZN(g30382), .A(II39951) );
  INV_X1 NOT_12864( .ZN(g30383), .A(g30306) );
  INV_X1 NOT_12865( .ZN(II39976), .A(g30245) );
  INV_X1 NOT_12866( .ZN(g30408), .A(II39976) );
  INV_X1 NOT_12867( .ZN(II39982), .A(g30305) );
  INV_X1 NOT_12868( .ZN(g30412), .A(II39982) );
  INV_X1 NOT_12869( .ZN(II39985), .A(g30246) );
  INV_X1 NOT_12870( .ZN(g30435), .A(II39985) );
  INV_X1 NOT_12871( .ZN(II39991), .A(g30247) );
  INV_X1 NOT_12872( .ZN(g30439), .A(II39991) );
  INV_X1 NOT_12873( .ZN(II39997), .A(g30248) );
  INV_X1 NOT_12874( .ZN(g30443), .A(II39997) );
  INV_X1 NOT_12875( .ZN(II40002), .A(g30249) );
  INV_X1 NOT_12876( .ZN(g30446), .A(II40002) );
  INV_X1 NOT_12877( .ZN(II40008), .A(g30250) );
  INV_X1 NOT_12878( .ZN(g30450), .A(II40008) );
  INV_X1 NOT_12879( .ZN(II40016), .A(g30251) );
  INV_X1 NOT_12880( .ZN(g30456), .A(II40016) );
  INV_X1 NOT_12881( .ZN(II40021), .A(g30252) );
  INV_X1 NOT_12882( .ZN(g30459), .A(II40021) );
  INV_X1 NOT_12883( .ZN(II40027), .A(g30253) );
  INV_X1 NOT_12884( .ZN(g30463), .A(II40027) );
  INV_X1 NOT_12885( .ZN(II40032), .A(g30254) );
  INV_X1 NOT_12886( .ZN(g30466), .A(II40032) );
  INV_X1 NOT_12887( .ZN(II40039), .A(g30255) );
  INV_X1 NOT_12888( .ZN(g30471), .A(II40039) );
  INV_X1 NOT_12889( .ZN(II40044), .A(g30256) );
  INV_X1 NOT_12890( .ZN(g30474), .A(II40044) );
  INV_X1 NOT_12891( .ZN(II40051), .A(g30257) );
  INV_X1 NOT_12892( .ZN(g30479), .A(II40051) );
  INV_X1 NOT_12893( .ZN(II40054), .A(g30258) );
  INV_X1 NOT_12894( .ZN(g30480), .A(II40054) );
  INV_X1 NOT_12895( .ZN(II40059), .A(g30259) );
  INV_X1 NOT_12896( .ZN(g30483), .A(II40059) );
  INV_X1 NOT_12897( .ZN(II40066), .A(g30260) );
  INV_X1 NOT_12898( .ZN(g30488), .A(II40066) );
  INV_X1 NOT_12899( .ZN(II40071), .A(g30261) );
  INV_X1 NOT_12900( .ZN(g30491), .A(II40071) );
  INV_X1 NOT_12901( .ZN(II40075), .A(g30262) );
  INV_X1 NOT_12902( .ZN(g30493), .A(II40075) );
  INV_X1 NOT_12903( .ZN(II40078), .A(g30263) );
  INV_X1 NOT_12904( .ZN(g30494), .A(II40078) );
  INV_X1 NOT_12905( .ZN(II40083), .A(g30264) );
  INV_X1 NOT_12906( .ZN(g30497), .A(II40083) );
  INV_X1 NOT_12907( .ZN(II40086), .A(g30265) );
  INV_X1 NOT_12908( .ZN(g30498), .A(II40086) );
  INV_X1 NOT_12909( .ZN(II40091), .A(g30266) );
  INV_X1 NOT_12910( .ZN(g30501), .A(II40091) );
  INV_X1 NOT_12911( .ZN(II40098), .A(g30491) );
  INV_X1 NOT_12912( .ZN(g30506), .A(II40098) );
  INV_X1 NOT_12913( .ZN(II40101), .A(g30326) );
  INV_X1 NOT_12914( .ZN(g30507), .A(II40101) );
  INV_X1 NOT_12915( .ZN(II40104), .A(g30342) );
  INV_X1 NOT_12916( .ZN(g30508), .A(II40104) );
  INV_X1 NOT_12917( .ZN(II40107), .A(g30343) );
  INV_X1 NOT_12918( .ZN(g30509), .A(II40107) );
  INV_X1 NOT_12919( .ZN(II40110), .A(g30357) );
  INV_X1 NOT_12920( .ZN(g30510), .A(II40110) );
  INV_X1 NOT_12921( .ZN(II40113), .A(g30368) );
  INV_X1 NOT_12922( .ZN(g30511), .A(II40113) );
  INV_X1 NOT_12923( .ZN(II40116), .A(g30408) );
  INV_X1 NOT_12924( .ZN(g30512), .A(II40116) );
  INV_X1 NOT_12925( .ZN(II40119), .A(g30435) );
  INV_X1 NOT_12926( .ZN(g30513), .A(II40119) );
  INV_X1 NOT_12927( .ZN(II40122), .A(g30443) );
  INV_X1 NOT_12928( .ZN(g30514), .A(II40122) );
  INV_X1 NOT_12929( .ZN(II40125), .A(g30466) );
  INV_X1 NOT_12930( .ZN(g30515), .A(II40125) );
  INV_X1 NOT_12931( .ZN(II40128), .A(g30479) );
  INV_X1 NOT_12932( .ZN(g30516), .A(II40128) );
  INV_X1 NOT_12933( .ZN(II40131), .A(g30493) );
  INV_X1 NOT_12934( .ZN(g30517), .A(II40131) );
  INV_X1 NOT_12935( .ZN(II40134), .A(g30480) );
  INV_X1 NOT_12936( .ZN(g30518), .A(II40134) );
  INV_X1 NOT_12937( .ZN(II40137), .A(g30494) );
  INV_X1 NOT_12938( .ZN(g30519), .A(II40137) );
  INV_X1 NOT_12939( .ZN(II40140), .A(g30328) );
  INV_X1 NOT_12940( .ZN(g30520), .A(II40140) );
  INV_X1 NOT_12941( .ZN(II40143), .A(g30329) );
  INV_X1 NOT_12942( .ZN(g30521), .A(II40143) );
  INV_X1 NOT_12943( .ZN(II40146), .A(g30344) );
  INV_X1 NOT_12944( .ZN(g30522), .A(II40146) );
  INV_X1 NOT_12945( .ZN(II40149), .A(g30358) );
  INV_X1 NOT_12946( .ZN(g30523), .A(II40149) );
  INV_X1 NOT_12947( .ZN(II40152), .A(g30359) );
  INV_X1 NOT_12948( .ZN(g30524), .A(II40152) );
  INV_X1 NOT_12949( .ZN(II40155), .A(g30369) );
  INV_X1 NOT_12950( .ZN(g30525), .A(II40155) );
  INV_X1 NOT_12951( .ZN(II40158), .A(g30376) );
  INV_X1 NOT_12952( .ZN(g30526), .A(II40158) );
  INV_X1 NOT_12953( .ZN(II40161), .A(g30439) );
  INV_X1 NOT_12954( .ZN(g30527), .A(II40161) );
  INV_X1 NOT_12955( .ZN(II40164), .A(g30446) );
  INV_X1 NOT_12956( .ZN(g30528), .A(II40164) );
  INV_X1 NOT_12957( .ZN(II40167), .A(g30456) );
  INV_X1 NOT_12958( .ZN(g30529), .A(II40167) );
  INV_X1 NOT_12959( .ZN(II40170), .A(g30483) );
  INV_X1 NOT_12960( .ZN(g30530), .A(II40170) );
  INV_X1 NOT_12961( .ZN(II40173), .A(g30497) );
  INV_X1 NOT_12962( .ZN(g30531), .A(II40173) );
  INV_X1 NOT_12963( .ZN(II40176), .A(g30331) );
  INV_X1 NOT_12964( .ZN(g30532), .A(II40176) );
  INV_X1 NOT_12965( .ZN(II40179), .A(g30498) );
  INV_X1 NOT_12966( .ZN(g30533), .A(II40179) );
  INV_X1 NOT_12967( .ZN(II40182), .A(g30332) );
  INV_X1 NOT_12968( .ZN(g30534), .A(II40182) );
  INV_X1 NOT_12969( .ZN(II40185), .A(g30346) );
  INV_X1 NOT_12970( .ZN(g30535), .A(II40185) );
  INV_X1 NOT_12971( .ZN(II40188), .A(g30347) );
  INV_X1 NOT_12972( .ZN(g30536), .A(II40188) );
  INV_X1 NOT_12973( .ZN(II40191), .A(g30360) );
  INV_X1 NOT_12974( .ZN(g30537), .A(II40191) );
  INV_X1 NOT_12975( .ZN(II40194), .A(g30370) );
  INV_X1 NOT_12976( .ZN(g30538), .A(II40194) );
  INV_X1 NOT_12977( .ZN(II40197), .A(g30371) );
  INV_X1 NOT_12978( .ZN(g30539), .A(II40197) );
  INV_X1 NOT_12979( .ZN(II40200), .A(g30377) );
  INV_X1 NOT_12980( .ZN(g30540), .A(II40200) );
  INV_X1 NOT_12981( .ZN(II40203), .A(g30380) );
  INV_X1 NOT_12982( .ZN(g30541), .A(II40203) );
  INV_X1 NOT_12983( .ZN(II40206), .A(g30450) );
  INV_X1 NOT_12984( .ZN(g30542), .A(II40206) );
  INV_X1 NOT_12985( .ZN(II40209), .A(g30459) );
  INV_X1 NOT_12986( .ZN(g30543), .A(II40209) );
  INV_X1 NOT_12987( .ZN(II40212), .A(g30471) );
  INV_X1 NOT_12988( .ZN(g30544), .A(II40212) );
  INV_X1 NOT_12989( .ZN(II40215), .A(g30501) );
  INV_X1 NOT_12990( .ZN(g30545), .A(II40215) );
  INV_X1 NOT_12991( .ZN(II40218), .A(g30335) );
  INV_X1 NOT_12992( .ZN(g30546), .A(II40218) );
  INV_X1 NOT_12993( .ZN(II40221), .A(g30349) );
  INV_X1 NOT_12994( .ZN(g30547), .A(II40221) );
  INV_X1 NOT_12995( .ZN(II40224), .A(g30336) );
  INV_X1 NOT_12996( .ZN(g30548), .A(II40224) );
  INV_X1 NOT_12997( .ZN(II40227), .A(g30350) );
  INV_X1 NOT_12998( .ZN(g30549), .A(II40227) );
  INV_X1 NOT_12999( .ZN(II40230), .A(g30362) );
  INV_X1 NOT_13000( .ZN(g30550), .A(II40230) );
  INV_X1 NOT_13001( .ZN(II40233), .A(g30363) );
  INV_X1 NOT_13002( .ZN(g30551), .A(II40233) );
  INV_X1 NOT_13003( .ZN(II40236), .A(g30373) );
  INV_X1 NOT_13004( .ZN(g30552), .A(II40236) );
  INV_X1 NOT_13005( .ZN(II40239), .A(g30378) );
  INV_X1 NOT_13006( .ZN(g30553), .A(II40239) );
  INV_X1 NOT_13007( .ZN(II40242), .A(g30379) );
  INV_X1 NOT_13008( .ZN(g30554), .A(II40242) );
  INV_X1 NOT_13009( .ZN(II40245), .A(g30381) );
  INV_X1 NOT_13010( .ZN(g30555), .A(II40245) );
  INV_X1 NOT_13011( .ZN(II40248), .A(g30382) );
  INV_X1 NOT_13012( .ZN(g30556), .A(II40248) );
  INV_X1 NOT_13013( .ZN(II40251), .A(g30463) );
  INV_X1 NOT_13014( .ZN(g30557), .A(II40251) );
  INV_X1 NOT_13015( .ZN(II40254), .A(g30474) );
  INV_X1 NOT_13016( .ZN(g30558), .A(II40254) );
  INV_X1 NOT_13017( .ZN(II40257), .A(g30488) );
  INV_X1 NOT_13018( .ZN(g30559), .A(II40257) );
  INV_X1 NOT_13019( .ZN(II40260), .A(g30339) );
  INV_X1 NOT_13020( .ZN(g30560), .A(II40260) );
  INV_X1 NOT_13021( .ZN(II40263), .A(g30353) );
  INV_X1 NOT_13022( .ZN(g30561), .A(II40263) );
  INV_X1 NOT_13023( .ZN(II40266), .A(g30365) );
  INV_X1 NOT_13024( .ZN(g30562), .A(II40266) );
  INV_X1 NOT_13025( .ZN(II40269), .A(g30354) );
  INV_X1 NOT_13026( .ZN(g30563), .A(II40269) );
  INV_X1 NOT_13027( .ZN(II40272), .A(g30366) );
  INV_X1 NOT_13028( .ZN(g30564), .A(II40272) );
  INV_X1 NOT_13029( .ZN(II40275), .A(g30375) );
  INV_X1 NOT_13030( .ZN(g30565), .A(II40275) );
  INV_X1 NOT_13031( .ZN(g30567), .A(g30403) );
  INV_X1 NOT_13032( .ZN(g30568), .A(g30402) );
  INV_X1 NOT_13033( .ZN(g30569), .A(g30406) );
  INV_X1 NOT_13034( .ZN(g30570), .A(g30404) );
  INV_X1 NOT_13035( .ZN(g30571), .A(g30401) );
  INV_X1 NOT_13036( .ZN(g30572), .A(g30399) );
  INV_X1 NOT_13037( .ZN(g30573), .A(g30405) );
  INV_X1 NOT_13038( .ZN(g30574), .A(g30400) );
  INV_X1 NOT_13039( .ZN(g30575), .A(g30412) );
  INV_X1 NOT_13040( .ZN(II40288), .A(g30455) );
  INV_X1 NOT_13041( .ZN(g30578), .A(II40288) );
  INV_X1 NOT_13042( .ZN(II40291), .A(g30468) );
  INV_X1 NOT_13043( .ZN(g30579), .A(II40291) );
  INV_X1 NOT_13044( .ZN(II40294), .A(g30470) );
  INV_X1 NOT_13045( .ZN(g30580), .A(II40294) );
  INV_X1 NOT_13046( .ZN(II40297), .A(g30482) );
  INV_X1 NOT_13047( .ZN(g30581), .A(II40297) );
  INV_X1 NOT_13048( .ZN(II40300), .A(g30485) );
  INV_X1 NOT_13049( .ZN(g30582), .A(II40300) );
  INV_X1 NOT_13050( .ZN(II40303), .A(g30487) );
  INV_X1 NOT_13051( .ZN(g30583), .A(II40303) );
  INV_X1 NOT_13052( .ZN(II40307), .A(g30500) );
  INV_X1 NOT_13053( .ZN(g30585), .A(II40307) );
  INV_X1 NOT_13054( .ZN(II40310), .A(g30503) );
  INV_X1 NOT_13055( .ZN(g30586), .A(II40310) );
  INV_X1 NOT_13056( .ZN(II40313), .A(g30505) );
  INV_X1 NOT_13057( .ZN(g30587), .A(II40313) );
  INV_X1 NOT_13058( .ZN(II40317), .A(g30338) );
  INV_X1 NOT_13059( .ZN(g30591), .A(II40317) );
  INV_X1 NOT_13060( .ZN(II40320), .A(g30341) );
  INV_X1 NOT_13061( .ZN(g30592), .A(II40320) );
  INV_X1 NOT_13062( .ZN(II40326), .A(g30356) );
  INV_X1 NOT_13063( .ZN(g30600), .A(II40326) );
  INV_X1 NOT_13064( .ZN(II40420), .A(g30578) );
  INV_X1 NOT_13065( .ZN(g30710), .A(II40420) );
  INV_X1 NOT_13066( .ZN(II40423), .A(g30579) );
  INV_X1 NOT_13067( .ZN(g30711), .A(II40423) );
  INV_X1 NOT_13068( .ZN(II40426), .A(g30581) );
  INV_X1 NOT_13069( .ZN(g30712), .A(II40426) );
  INV_X1 NOT_13070( .ZN(II40429), .A(g30580) );
  INV_X1 NOT_13071( .ZN(g30713), .A(II40429) );
  INV_X1 NOT_13072( .ZN(II40432), .A(g30582) );
  INV_X1 NOT_13073( .ZN(g30714), .A(II40432) );
  INV_X1 NOT_13074( .ZN(II40435), .A(g30585) );
  INV_X1 NOT_13075( .ZN(g30715), .A(II40435) );
  INV_X1 NOT_13076( .ZN(II40438), .A(g30583) );
  INV_X1 NOT_13077( .ZN(g30716), .A(II40438) );
  INV_X1 NOT_13078( .ZN(II40441), .A(g30586) );
  INV_X1 NOT_13079( .ZN(g30717), .A(II40441) );
  INV_X1 NOT_13080( .ZN(II40444), .A(g30591) );
  INV_X1 NOT_13081( .ZN(g30718), .A(II40444) );
  INV_X1 NOT_13082( .ZN(II40447), .A(g30587) );
  INV_X1 NOT_13083( .ZN(g30719), .A(II40447) );
  INV_X1 NOT_13084( .ZN(II40450), .A(g30592) );
  INV_X1 NOT_13085( .ZN(g30720), .A(II40450) );
  INV_X1 NOT_13086( .ZN(II40453), .A(g30600) );
  INV_X1 NOT_13087( .ZN(g30721), .A(II40453) );
  INV_X1 NOT_13088( .ZN(II40456), .A(g30668) );
  INV_X1 NOT_13089( .ZN(g30722), .A(II40456) );
  INV_X1 NOT_13090( .ZN(II40459), .A(g30669) );
  INV_X1 NOT_13091( .ZN(g30723), .A(II40459) );
  INV_X1 NOT_13092( .ZN(II40462), .A(g30670) );
  INV_X1 NOT_13093( .ZN(g30724), .A(II40462) );
  INV_X1 NOT_13094( .ZN(II40465), .A(g30671) );
  INV_X1 NOT_13095( .ZN(g30725), .A(II40465) );
  INV_X1 NOT_13096( .ZN(II40468), .A(g30672) );
  INV_X1 NOT_13097( .ZN(g30726), .A(II40468) );
  INV_X1 NOT_13098( .ZN(II40471), .A(g30673) );
  INV_X1 NOT_13099( .ZN(g30727), .A(II40471) );
  INV_X1 NOT_13100( .ZN(II40475), .A(g30674) );
  INV_X1 NOT_13101( .ZN(g30729), .A(II40475) );
  INV_X1 NOT_13102( .ZN(II40478), .A(g30675) );
  INV_X1 NOT_13103( .ZN(g30730), .A(II40478) );
  INV_X1 NOT_13104( .ZN(II40481), .A(g30676) );
  INV_X1 NOT_13105( .ZN(g30731), .A(II40481) );
  INV_X1 NOT_13106( .ZN(II40484), .A(g30677) );
  INV_X1 NOT_13107( .ZN(g30732), .A(II40484) );
  INV_X1 NOT_13108( .ZN(II40487), .A(g30678) );
  INV_X1 NOT_13109( .ZN(g30733), .A(II40487) );
  INV_X1 NOT_13110( .ZN(II40490), .A(g30679) );
  INV_X1 NOT_13111( .ZN(g30734), .A(II40490) );
  INV_X1 NOT_13112( .ZN(II40495), .A(g30680) );
  INV_X1 NOT_13113( .ZN(g30737), .A(II40495) );
  INV_X1 NOT_13114( .ZN(II40498), .A(g30681) );
  INV_X1 NOT_13115( .ZN(g30738), .A(II40498) );
  INV_X1 NOT_13116( .ZN(II40501), .A(g30682) );
  INV_X1 NOT_13117( .ZN(g30739), .A(II40501) );
  INV_X1 NOT_13118( .ZN(II40504), .A(g30683) );
  INV_X1 NOT_13119( .ZN(g30740), .A(II40504) );
  INV_X1 NOT_13120( .ZN(II40507), .A(g30684) );
  INV_X1 NOT_13121( .ZN(g30741), .A(II40507) );
  INV_X1 NOT_13122( .ZN(II40510), .A(g30686) );
  INV_X1 NOT_13123( .ZN(g30742), .A(II40510) );
  INV_X1 NOT_13124( .ZN(II40515), .A(g30687) );
  INV_X1 NOT_13125( .ZN(g30745), .A(II40515) );
  INV_X1 NOT_13126( .ZN(II40518), .A(g30688) );
  INV_X1 NOT_13127( .ZN(g30746), .A(II40518) );
  INV_X1 NOT_13128( .ZN(II40521), .A(g30689) );
  INV_X1 NOT_13129( .ZN(g30747), .A(II40521) );
  INV_X1 NOT_13130( .ZN(II40524), .A(g30690) );
  INV_X1 NOT_13131( .ZN(g30748), .A(II40524) );
  INV_X1 NOT_13132( .ZN(II40527), .A(g30691) );
  INV_X1 NOT_13133( .ZN(g30749), .A(II40527) );
  INV_X1 NOT_13134( .ZN(II40531), .A(g30692) );
  INV_X1 NOT_13135( .ZN(g30751), .A(II40531) );
  INV_X1 NOT_13136( .ZN(II40534), .A(g30693) );
  INV_X1 NOT_13137( .ZN(g30752), .A(II40534) );
  INV_X1 NOT_13138( .ZN(II40537), .A(g30694) );
  INV_X1 NOT_13139( .ZN(g30753), .A(II40537) );
  INV_X1 NOT_13140( .ZN(II40542), .A(g30695) );
  INV_X1 NOT_13141( .ZN(g30756), .A(II40542) );
  INV_X1 NOT_13142( .ZN(g30765), .A(g30685) );
  INV_X1 NOT_13143( .ZN(II40555), .A(g30699) );
  INV_X1 NOT_13144( .ZN(g30767), .A(II40555) );
  INV_X1 NOT_13145( .ZN(II40565), .A(g30700) );
  INV_X1 NOT_13146( .ZN(g30769), .A(II40565) );
  INV_X1 NOT_13147( .ZN(II40568), .A(g30701) );
  INV_X1 NOT_13148( .ZN(g30770), .A(II40568) );
  INV_X1 NOT_13149( .ZN(II40578), .A(g30702) );
  INV_X1 NOT_13150( .ZN(g30772), .A(II40578) );
  INV_X1 NOT_13151( .ZN(II40581), .A(g30703) );
  INV_X1 NOT_13152( .ZN(g30773), .A(II40581) );
  INV_X1 NOT_13153( .ZN(II40584), .A(g30704) );
  INV_X1 NOT_13154( .ZN(g30774), .A(II40584) );
  INV_X1 NOT_13155( .ZN(II40594), .A(g30705) );
  INV_X1 NOT_13156( .ZN(g30776), .A(II40594) );
  INV_X1 NOT_13157( .ZN(II40597), .A(g30706) );
  INV_X1 NOT_13158( .ZN(g30777), .A(II40597) );
  INV_X1 NOT_13159( .ZN(II40600), .A(g30707) );
  INV_X1 NOT_13160( .ZN(g30778), .A(II40600) );
  INV_X1 NOT_13161( .ZN(II40611), .A(g30708) );
  INV_X1 NOT_13162( .ZN(g30781), .A(II40611) );
  INV_X1 NOT_13163( .ZN(II40614), .A(g30709) );
  INV_X1 NOT_13164( .ZN(g30782), .A(II40614) );
  INV_X1 NOT_13165( .ZN(II40618), .A(g30566) );
  INV_X1 NOT_13166( .ZN(g30784), .A(II40618) );
  INV_X1 NOT_13167( .ZN(II40634), .A(g30571) );
  INV_X1 NOT_13168( .ZN(g30792), .A(II40634) );
  INV_X1 NOT_13169( .ZN(II40637), .A(g30570) );
  INV_X1 NOT_13170( .ZN(g30793), .A(II40637) );
  INV_X1 NOT_13171( .ZN(II40640), .A(g30569) );
  INV_X1 NOT_13172( .ZN(g30794), .A(II40640) );
  INV_X1 NOT_13173( .ZN(II40643), .A(g30568) );
  INV_X1 NOT_13174( .ZN(g30795), .A(II40643) );
  INV_X1 NOT_13175( .ZN(II40647), .A(g30567) );
  INV_X1 NOT_13176( .ZN(g30797), .A(II40647) );
  INV_X1 NOT_13177( .ZN(II40651), .A(g30574) );
  INV_X1 NOT_13178( .ZN(g30799), .A(II40651) );
  INV_X1 NOT_13179( .ZN(II40654), .A(g30573) );
  INV_X1 NOT_13180( .ZN(g30800), .A(II40654) );
  INV_X1 NOT_13181( .ZN(II40658), .A(g30572) );
  INV_X1 NOT_13182( .ZN(g30802), .A(II40658) );
  INV_X1 NOT_13183( .ZN(II40661), .A(g30635) );
  INV_X1 NOT_13184( .ZN(g30803), .A(II40661) );
  INV_X1 NOT_13185( .ZN(II40664), .A(g30636) );
  INV_X1 NOT_13186( .ZN(g30804), .A(II40664) );
  INV_X1 NOT_13187( .ZN(II40667), .A(g30637) );
  INV_X1 NOT_13188( .ZN(g30805), .A(II40667) );
  INV_X1 NOT_13189( .ZN(II40670), .A(g30638) );
  INV_X1 NOT_13190( .ZN(g30806), .A(II40670) );
  INV_X1 NOT_13191( .ZN(II40673), .A(g30639) );
  INV_X1 NOT_13192( .ZN(g30807), .A(II40673) );
  INV_X1 NOT_13193( .ZN(II40676), .A(g30640) );
  INV_X1 NOT_13194( .ZN(g30808), .A(II40676) );
  INV_X1 NOT_13195( .ZN(II40679), .A(g30641) );
  INV_X1 NOT_13196( .ZN(g30809), .A(II40679) );
  INV_X1 NOT_13197( .ZN(II40682), .A(g30642) );
  INV_X1 NOT_13198( .ZN(g30810), .A(II40682) );
  INV_X1 NOT_13199( .ZN(II40685), .A(g30643) );
  INV_X1 NOT_13200( .ZN(g30811), .A(II40685) );
  INV_X1 NOT_13201( .ZN(II40688), .A(g30644) );
  INV_X1 NOT_13202( .ZN(g30812), .A(II40688) );
  INV_X1 NOT_13203( .ZN(II40691), .A(g30645) );
  INV_X1 NOT_13204( .ZN(g30813), .A(II40691) );
  INV_X32 NOT_13205( .ZN(II40694), .A(g30646) );
  INV_X32 NOT_13206( .ZN(g30814), .A(II40694) );
  INV_X1 NOT_13207( .ZN(II40697), .A(g30647) );
  INV_X1 NOT_13208( .ZN(g30815), .A(II40697) );
  INV_X1 NOT_13209( .ZN(II40700), .A(g30648) );
  INV_X1 NOT_13210( .ZN(g30816), .A(II40700) );
  INV_X1 NOT_13211( .ZN(II40703), .A(g30649) );
  INV_X1 NOT_13212( .ZN(g30817), .A(II40703) );
  INV_X1 NOT_13213( .ZN(II40706), .A(g30650) );
  INV_X1 NOT_13214( .ZN(g30818), .A(II40706) );
  INV_X1 NOT_13215( .ZN(II40709), .A(g30651) );
  INV_X1 NOT_13216( .ZN(g30819), .A(II40709) );
  INV_X1 NOT_13217( .ZN(II40712), .A(g30652) );
  INV_X1 NOT_13218( .ZN(g30820), .A(II40712) );
  INV_X1 NOT_13219( .ZN(II40715), .A(g30653) );
  INV_X1 NOT_13220( .ZN(g30821), .A(II40715) );
  INV_X1 NOT_13221( .ZN(II40718), .A(g30654) );
  INV_X1 NOT_13222( .ZN(g30822), .A(II40718) );
  INV_X1 NOT_13223( .ZN(II40721), .A(g30655) );
  INV_X1 NOT_13224( .ZN(g30823), .A(II40721) );
  INV_X1 NOT_13225( .ZN(II40724), .A(g30656) );
  INV_X1 NOT_13226( .ZN(g30824), .A(II40724) );
  INV_X1 NOT_13227( .ZN(II40727), .A(g30657) );
  INV_X1 NOT_13228( .ZN(g30825), .A(II40727) );
  INV_X1 NOT_13229( .ZN(II40730), .A(g30658) );
  INV_X1 NOT_13230( .ZN(g30826), .A(II40730) );
  INV_X1 NOT_13231( .ZN(II40733), .A(g30659) );
  INV_X1 NOT_13232( .ZN(g30827), .A(II40733) );
  INV_X1 NOT_13233( .ZN(II40736), .A(g30660) );
  INV_X1 NOT_13234( .ZN(g30828), .A(II40736) );
  INV_X1 NOT_13235( .ZN(II40739), .A(g30661) );
  INV_X1 NOT_13236( .ZN(g30829), .A(II40739) );
  INV_X1 NOT_13237( .ZN(II40742), .A(g30662) );
  INV_X1 NOT_13238( .ZN(g30830), .A(II40742) );
  INV_X1 NOT_13239( .ZN(II40745), .A(g30663) );
  INV_X1 NOT_13240( .ZN(g30831), .A(II40745) );
  INV_X1 NOT_13241( .ZN(II40748), .A(g30664) );
  INV_X1 NOT_13242( .ZN(g30832), .A(II40748) );
  INV_X1 NOT_13243( .ZN(II40751), .A(g30665) );
  INV_X1 NOT_13244( .ZN(g30833), .A(II40751) );
  INV_X1 NOT_13245( .ZN(II40754), .A(g30666) );
  INV_X1 NOT_13246( .ZN(g30834), .A(II40754) );
  INV_X1 NOT_13247( .ZN(II40757), .A(g30667) );
  INV_X1 NOT_13248( .ZN(g30835), .A(II40757) );
  INV_X1 NOT_13249( .ZN(II40760), .A(g30722) );
  INV_X1 NOT_13250( .ZN(g30836), .A(II40760) );
  INV_X1 NOT_13251( .ZN(II40763), .A(g30729) );
  INV_X1 NOT_13252( .ZN(g30837), .A(II40763) );
  INV_X1 NOT_13253( .ZN(II40766), .A(g30737) );
  INV_X1 NOT_13254( .ZN(g30838), .A(II40766) );
  INV_X1 NOT_13255( .ZN(II40769), .A(g30803) );
  INV_X1 NOT_13256( .ZN(g30839), .A(II40769) );
  INV_X1 NOT_13257( .ZN(II40772), .A(g30804) );
  INV_X1 NOT_13258( .ZN(g30840), .A(II40772) );
  INV_X1 NOT_13259( .ZN(II40775), .A(g30807) );
  INV_X1 NOT_13260( .ZN(g30841), .A(II40775) );
  INV_X1 NOT_13261( .ZN(II40778), .A(g30805) );
  INV_X1 NOT_13262( .ZN(g30842), .A(II40778) );
  INV_X1 NOT_13263( .ZN(II40781), .A(g30808) );
  INV_X1 NOT_13264( .ZN(g30843), .A(II40781) );
  INV_X1 NOT_13265( .ZN(II40784), .A(g30813) );
  INV_X1 NOT_13266( .ZN(g30844), .A(II40784) );
  INV_X1 NOT_13267( .ZN(II40787), .A(g30809) );
  INV_X1 NOT_13268( .ZN(g30845), .A(II40787) );
  INV_X1 NOT_13269( .ZN(II40790), .A(g30814) );
  INV_X1 NOT_13270( .ZN(g30846), .A(II40790) );
  INV_X1 NOT_13271( .ZN(II40793), .A(g30821) );
  INV_X1 NOT_13272( .ZN(g30847), .A(II40793) );
  INV_X1 NOT_13273( .ZN(II40796), .A(g30829) );
  INV_X1 NOT_13274( .ZN(g30848), .A(II40796) );
  INV_X1 NOT_13275( .ZN(II40799), .A(g30723) );
  INV_X1 NOT_13276( .ZN(g30849), .A(II40799) );
  INV_X1 NOT_13277( .ZN(II40802), .A(g30730) );
  INV_X1 NOT_13278( .ZN(g30850), .A(II40802) );
  INV_X1 NOT_13279( .ZN(II40805), .A(g30767) );
  INV_X1 NOT_13280( .ZN(g30851), .A(II40805) );
  INV_X1 NOT_13281( .ZN(II40808), .A(g30769) );
  INV_X1 NOT_13282( .ZN(g30852), .A(II40808) );
  INV_X1 NOT_13283( .ZN(II40811), .A(g30772) );
  INV_X1 NOT_13284( .ZN(g30853), .A(II40811) );
  INV_X1 NOT_13285( .ZN(II40814), .A(g30731) );
  INV_X1 NOT_13286( .ZN(g30854), .A(II40814) );
  INV_X1 NOT_13287( .ZN(II40817), .A(g30738) );
  INV_X1 NOT_13288( .ZN(g30855), .A(II40817) );
  INV_X1 NOT_13289( .ZN(II40820), .A(g30745) );
  INV_X1 NOT_13290( .ZN(g30856), .A(II40820) );
  INV_X1 NOT_13291( .ZN(II40823), .A(g30806) );
  INV_X1 NOT_13292( .ZN(g30857), .A(II40823) );
  INV_X1 NOT_13293( .ZN(II40826), .A(g30810) );
  INV_X1 NOT_13294( .ZN(g30858), .A(II40826) );
  INV_X1 NOT_13295( .ZN(II40829), .A(g30815) );
  INV_X1 NOT_13296( .ZN(g30859), .A(II40829) );
  INV_X1 NOT_13297( .ZN(II40832), .A(g30811) );
  INV_X1 NOT_13298( .ZN(g30860), .A(II40832) );
  INV_X1 NOT_13299( .ZN(II40835), .A(g30816) );
  INV_X1 NOT_13300( .ZN(g30861), .A(II40835) );
  INV_X1 NOT_13301( .ZN(II40838), .A(g30822) );
  INV_X1 NOT_13302( .ZN(g30862), .A(II40838) );
  INV_X1 NOT_13303( .ZN(II40841), .A(g30817) );
  INV_X1 NOT_13304( .ZN(g30863), .A(II40841) );
  INV_X1 NOT_13305( .ZN(II40844), .A(g30823) );
  INV_X1 NOT_13306( .ZN(g30864), .A(II40844) );
  INV_X1 NOT_13307( .ZN(II40847), .A(g30830) );
  INV_X1 NOT_13308( .ZN(g30865), .A(II40847) );
  INV_X1 NOT_13309( .ZN(II40850), .A(g30724) );
  INV_X1 NOT_13310( .ZN(g30866), .A(II40850) );
  INV_X1 NOT_13311( .ZN(II40853), .A(g30732) );
  INV_X1 NOT_13312( .ZN(g30867), .A(II40853) );
  INV_X1 NOT_13313( .ZN(II40856), .A(g30739) );
  INV_X1 NOT_13314( .ZN(g30868), .A(II40856) );
  INV_X1 NOT_13315( .ZN(II40859), .A(g30770) );
  INV_X1 NOT_13316( .ZN(g30869), .A(II40859) );
  INV_X1 NOT_13317( .ZN(II40862), .A(g30773) );
  INV_X1 NOT_13318( .ZN(g30870), .A(II40862) );
  INV_X1 NOT_13319( .ZN(II40865), .A(g30776) );
  INV_X1 NOT_13320( .ZN(g30871), .A(II40865) );
  INV_X1 NOT_13321( .ZN(II40868), .A(g30740) );
  INV_X1 NOT_13322( .ZN(g30872), .A(II40868) );
  INV_X1 NOT_13323( .ZN(II40871), .A(g30746) );
  INV_X1 NOT_13324( .ZN(g30873), .A(II40871) );
  INV_X1 NOT_13325( .ZN(II40874), .A(g30751) );
  INV_X1 NOT_13326( .ZN(g30874), .A(II40874) );
  INV_X1 NOT_13327( .ZN(II40877), .A(g30812) );
  INV_X1 NOT_13328( .ZN(g30875), .A(II40877) );
  INV_X1 NOT_13329( .ZN(II40880), .A(g30818) );
  INV_X1 NOT_13330( .ZN(g30876), .A(II40880) );
  INV_X1 NOT_13331( .ZN(II40883), .A(g30824) );
  INV_X1 NOT_13332( .ZN(g30877), .A(II40883) );
  INV_X1 NOT_13333( .ZN(II40886), .A(g30819) );
  INV_X1 NOT_13334( .ZN(g30878), .A(II40886) );
  INV_X1 NOT_13335( .ZN(II40889), .A(g30825) );
  INV_X1 NOT_13336( .ZN(g30879), .A(II40889) );
  INV_X1 NOT_13337( .ZN(II40892), .A(g30831) );
  INV_X1 NOT_13338( .ZN(g30880), .A(II40892) );
  INV_X1 NOT_13339( .ZN(II40895), .A(g30826) );
  INV_X1 NOT_13340( .ZN(g30881), .A(II40895) );
  INV_X1 NOT_13341( .ZN(II40898), .A(g30832) );
  INV_X1 NOT_13342( .ZN(g30882), .A(II40898) );
  INV_X1 NOT_13343( .ZN(II40901), .A(g30725) );
  INV_X1 NOT_13344( .ZN(g30883), .A(II40901) );
  INV_X1 NOT_13345( .ZN(II40904), .A(g30733) );
  INV_X1 NOT_13346( .ZN(g30884), .A(II40904) );
  INV_X1 NOT_13347( .ZN(II40907), .A(g30741) );
  INV_X1 NOT_13348( .ZN(g30885), .A(II40907) );
  INV_X1 NOT_13349( .ZN(II40910), .A(g30747) );
  INV_X1 NOT_13350( .ZN(g30886), .A(II40910) );
  INV_X1 NOT_13351( .ZN(II40913), .A(g30774) );
  INV_X1 NOT_13352( .ZN(g30887), .A(II40913) );
  INV_X1 NOT_13353( .ZN(II40916), .A(g30777) );
  INV_X1 NOT_13354( .ZN(g30888), .A(II40916) );
  INV_X1 NOT_13355( .ZN(II40919), .A(g30781) );
  INV_X1 NOT_13356( .ZN(g30889), .A(II40919) );
  INV_X1 NOT_13357( .ZN(II40922), .A(g30748) );
  INV_X1 NOT_13358( .ZN(g30890), .A(II40922) );
  INV_X1 NOT_13359( .ZN(II40925), .A(g30752) );
  INV_X1 NOT_13360( .ZN(g30891), .A(II40925) );
  INV_X1 NOT_13361( .ZN(II40928), .A(g30756) );
  INV_X1 NOT_13362( .ZN(g30892), .A(II40928) );
  INV_X1 NOT_13363( .ZN(II40931), .A(g30820) );
  INV_X1 NOT_13364( .ZN(g30893), .A(II40931) );
  INV_X1 NOT_13365( .ZN(II40934), .A(g30827) );
  INV_X1 NOT_13366( .ZN(g30894), .A(II40934) );
  INV_X1 NOT_13367( .ZN(II40937), .A(g30833) );
  INV_X1 NOT_13368( .ZN(g30895), .A(II40937) );
  INV_X1 NOT_13369( .ZN(II40940), .A(g30828) );
  INV_X1 NOT_13370( .ZN(g30896), .A(II40940) );
  INV_X1 NOT_13371( .ZN(II40943), .A(g30834) );
  INV_X1 NOT_13372( .ZN(g30897), .A(II40943) );
  INV_X1 NOT_13373( .ZN(II40946), .A(g30726) );
  INV_X1 NOT_13374( .ZN(g30898), .A(II40946) );
  INV_X1 NOT_13375( .ZN(II40949), .A(g30835) );
  INV_X1 NOT_13376( .ZN(g30899), .A(II40949) );
  INV_X8 NOT_13377( .ZN(II40952), .A(g30727) );
  INV_X8 NOT_13378( .ZN(g30900), .A(II40952) );
  INV_X8 NOT_13379( .ZN(II40955), .A(g30734) );
  INV_X8 NOT_13380( .ZN(g30901), .A(II40955) );
  INV_X1 NOT_13381( .ZN(II40958), .A(g30742) );
  INV_X1 NOT_13382( .ZN(g30902), .A(II40958) );
  INV_X1 NOT_13383( .ZN(II40961), .A(g30749) );
  INV_X1 NOT_13384( .ZN(g30903), .A(II40961) );
  INV_X1 NOT_13385( .ZN(II40964), .A(g30753) );
  INV_X1 NOT_13386( .ZN(g30904), .A(II40964) );
  INV_X1 NOT_13387( .ZN(II40967), .A(g30778) );
  INV_X1 NOT_13388( .ZN(g30905), .A(II40967) );
  INV_X1 NOT_13389( .ZN(II40970), .A(g30782) );
  INV_X1 NOT_13390( .ZN(g30906), .A(II40970) );
  INV_X1 NOT_13391( .ZN(II40973), .A(g30784) );
  INV_X1 NOT_13392( .ZN(g30907), .A(II40973) );
  INV_X1 NOT_13393( .ZN(II40976), .A(g30799) );
  INV_X1 NOT_13394( .ZN(g30908), .A(II40976) );
  INV_X1 NOT_13395( .ZN(II40979), .A(g30800) );
  INV_X1 NOT_13396( .ZN(g30909), .A(II40979) );
  INV_X1 NOT_13397( .ZN(II40982), .A(g30802) );
  INV_X1 NOT_13398( .ZN(g30910), .A(II40982) );
  INV_X1 NOT_13399( .ZN(II40985), .A(g30792) );
  INV_X1 NOT_13400( .ZN(g30911), .A(II40985) );
  INV_X1 NOT_13401( .ZN(II40988), .A(g30793) );
  INV_X1 NOT_13402( .ZN(g30912), .A(II40988) );
  INV_X1 NOT_13403( .ZN(II40991), .A(g30794) );
  INV_X1 NOT_13404( .ZN(g30913), .A(II40991) );
  INV_X1 NOT_13405( .ZN(II40994), .A(g30795) );
  INV_X1 NOT_13406( .ZN(g30914), .A(II40994) );
  INV_X1 NOT_13407( .ZN(II40997), .A(g30797) );
  INV_X1 NOT_13408( .ZN(g30915), .A(II40997) );
  INV_X1 NOT_13409( .ZN(II41024), .A(g30765) );
  INV_X1 NOT_13410( .ZN(g30928), .A(II41024) );
  INV_X1 NOT_13411( .ZN(II41035), .A(g30796) );
  INV_X1 NOT_13412( .ZN(g30937), .A(II41035) );
  INV_X1 NOT_13413( .ZN(II41038), .A(g30798) );
  INV_X1 NOT_13414( .ZN(g30938), .A(II41038) );
  INV_X1 NOT_13415( .ZN(II41041), .A(g30801) );
  INV_X1 NOT_13416( .ZN(g30939), .A(II41041) );
  INV_X1 NOT_13417( .ZN(II41044), .A(g30928) );
  INV_X1 NOT_13418( .ZN(g30940), .A(II41044) );
  INV_X1 NOT_13419( .ZN(II41047), .A(g30937) );
  INV_X1 NOT_13420( .ZN(g30941), .A(II41047) );
  INV_X1 NOT_13421( .ZN(II41050), .A(g30938) );
  INV_X1 NOT_13422( .ZN(g30942), .A(II41050) );
  INV_X1 NOT_13423( .ZN(II41053), .A(g30939) );
  INV_X1 NOT_13424( .ZN(g30943), .A(II41053) );
  INV_X1 NOT_13425( .ZN(g30962), .A(g30958) );
  INV_X1 NOT_13426( .ZN(g30963), .A(g30957) );
  INV_X1 NOT_13427( .ZN(g30964), .A(g30961) );
  INV_X1 NOT_13428( .ZN(g30965), .A(g30959) );
  INV_X1 NOT_13429( .ZN(g30966), .A(g30956) );
  INV_X1 NOT_13430( .ZN(g30967), .A(g30954) );
  INV_X1 NOT_13431( .ZN(g30968), .A(g30960) );
  INV_X1 NOT_13432( .ZN(g30969), .A(g30955) );
  INV_X1 NOT_13433( .ZN(g30971), .A(g30970) );
  INV_X1 NOT_13434( .ZN(II41090), .A(g30965) );
  INV_X1 NOT_13435( .ZN(g30972), .A(II41090) );
  INV_X1 NOT_13436( .ZN(II41093), .A(g30964) );
  INV_X1 NOT_13437( .ZN(g30973), .A(II41093) );
  INV_X1 NOT_13438( .ZN(II41096), .A(g30963) );
  INV_X1 NOT_13439( .ZN(g30974), .A(II41096) );
  INV_X1 NOT_13440( .ZN(II41099), .A(g30962) );
  INV_X1 NOT_13441( .ZN(g30975), .A(II41099) );
  INV_X1 NOT_13442( .ZN(II41102), .A(g30969) );
  INV_X1 NOT_13443( .ZN(g30976), .A(II41102) );
  INV_X1 NOT_13444( .ZN(II41105), .A(g30968) );
  INV_X1 NOT_13445( .ZN(g30977), .A(II41105) );
  INV_X1 NOT_13446( .ZN(II41108), .A(g30967) );
  INV_X1 NOT_13447( .ZN(g30978), .A(II41108) );
  INV_X1 NOT_13448( .ZN(II41111), .A(g30966) );
  INV_X1 NOT_13449( .ZN(g30979), .A(II41111) );
  INV_X1 NOT_13450( .ZN(II41114), .A(g30976) );
  INV_X1 NOT_13451( .ZN(g30980), .A(II41114) );
  INV_X1 NOT_13452( .ZN(II41117), .A(g30977) );
  INV_X1 NOT_13453( .ZN(g30981), .A(II41117) );
  INV_X1 NOT_13454( .ZN(II41120), .A(g30978) );
  INV_X1 NOT_13455( .ZN(g30982), .A(II41120) );
  INV_X1 NOT_13456( .ZN(II41123), .A(g30979) );
  INV_X1 NOT_13457( .ZN(g30983), .A(II41123) );
  INV_X1 NOT_13458( .ZN(II41126), .A(g30972) );
  INV_X1 NOT_13459( .ZN(g30984), .A(II41126) );
  INV_X1 NOT_13460( .ZN(II41129), .A(g30973) );
  INV_X1 NOT_13461( .ZN(g30985), .A(II41129) );
  INV_X1 NOT_13462( .ZN(II41132), .A(g30974) );
  INV_X1 NOT_13463( .ZN(g30986), .A(II41132) );
  INV_X1 NOT_13464( .ZN(II41135), .A(g30975) );
  INV_X1 NOT_13465( .ZN(g30987), .A(II41135) );
  INV_X1 NOT_13466( .ZN(II41138), .A(g30971) );
  INV_X1 NOT_13467( .ZN(g30988), .A(II41138) );
  INV_X1 NOT_13468( .ZN(II41141), .A(g30988) );
  INV_X1 NOT_13469( .ZN(g30989), .A(II41141) );
  AND2_X1 AND2_0( .ZN(g5630), .A1(g325), .A2(g349) );
  AND2_X1 AND2_1( .ZN(g5649), .A1(g331), .A2(g351) );
  AND2_X1 AND2_2( .ZN(g5650), .A1(g325), .A2(g364) );
  AND2_X1 AND2_3( .ZN(g5658), .A1(g1012), .A2(g1036) );
  AND2_X1 AND2_4( .ZN(g5676), .A1(g337), .A2(g353) );
  AND2_X1 AND2_5( .ZN(g5677), .A1(g331), .A2(g366) );
  AND2_X1 AND2_6( .ZN(g5678), .A1(g325), .A2(g379) );
  AND2_X1 AND2_7( .ZN(g5687), .A1(g1018), .A2(g1038) );
  AND2_X1 AND2_8( .ZN(g5688), .A1(g1012), .A2(g1051) );
  AND2_X1 AND2_9( .ZN(g5696), .A1(g1706), .A2(g1730) );
  AND2_X1 AND2_10( .ZN(g5709), .A1(g337), .A2(g368) );
  AND2_X1 AND2_11( .ZN(g5710), .A1(g331), .A2(g381) );
  AND2_X1 AND2_12( .ZN(g5711), .A1(g325), .A2(g394) );
  AND2_X1 AND2_13( .ZN(g5728), .A1(g1024), .A2(g1040) );
  AND2_X1 AND2_14( .ZN(g5729), .A1(g1018), .A2(g1053) );
  AND2_X1 AND2_15( .ZN(g5730), .A1(g1012), .A2(g1066) );
  AND2_X1 AND2_16( .ZN(g5739), .A1(g1712), .A2(g1732) );
  AND2_X1 AND2_17( .ZN(g5740), .A1(g1706), .A2(g1745) );
  AND2_X1 AND2_18( .ZN(g5748), .A1(g2400), .A2(g2424) );
  AND2_X1 AND2_19( .ZN(g5757), .A1(g337), .A2(g383) );
  AND2_X1 AND2_20( .ZN(g5758), .A1(g331), .A2(g396) );
  AND2_X1 AND2_21( .ZN(g5767), .A1(g1024), .A2(g1055) );
  AND2_X1 AND2_22( .ZN(g5768), .A1(g1018), .A2(g1068) );
  AND2_X1 AND2_23( .ZN(g5769), .A1(g1012), .A2(g1081) );
  AND2_X1 AND2_24( .ZN(g5786), .A1(g1718), .A2(g1734) );
  AND2_X1 AND2_25( .ZN(g5787), .A1(g1712), .A2(g1747) );
  AND2_X1 AND2_26( .ZN(g5788), .A1(g1706), .A2(g1760) );
  AND2_X1 AND2_27( .ZN(g5797), .A1(g2406), .A2(g2426) );
  AND2_X1 AND2_28( .ZN(g5798), .A1(g2400), .A2(g2439) );
  AND2_X1 AND2_29( .ZN(g5807), .A1(g337), .A2(g324) );
  AND2_X1 AND2_30( .ZN(g5816), .A1(g1024), .A2(g1070) );
  AND2_X1 AND2_31( .ZN(g5817), .A1(g1018), .A2(g1083) );
  AND2_X1 AND2_32( .ZN(g5826), .A1(g1718), .A2(g1749) );
  AND2_X1 AND2_33( .ZN(g5827), .A1(g1712), .A2(g1762) );
  AND2_X1 AND2_34( .ZN(g5828), .A1(g1706), .A2(g1775) );
  AND2_X1 AND2_35( .ZN(g5845), .A1(g2412), .A2(g2428) );
  AND2_X1 AND2_36( .ZN(g5846), .A1(g2406), .A2(g2441) );
  AND2_X1 AND2_37( .ZN(g5847), .A1(g2400), .A2(g2454) );
  AND2_X1 AND2_38( .ZN(g5863), .A1(g1024), .A2(g1011) );
  AND2_X1 AND2_39( .ZN(g5872), .A1(g1718), .A2(g1764) );
  AND2_X1 AND2_40( .ZN(g5873), .A1(g1712), .A2(g1777) );
  AND2_X1 AND2_41( .ZN(g5882), .A1(g2412), .A2(g2443) );
  AND2_X1 AND2_42( .ZN(g5883), .A1(g2406), .A2(g2456) );
  AND2_X1 AND2_43( .ZN(g5884), .A1(g2400), .A2(g2469) );
  AND2_X1 AND2_44( .ZN(g5910), .A1(g1718), .A2(g1705) );
  AND2_X1 AND2_45( .ZN(g5919), .A1(g2412), .A2(g2458) );
  AND2_X1 AND2_46( .ZN(g5920), .A1(g2406), .A2(g2471) );
  AND2_X1 AND2_47( .ZN(g5949), .A1(g2412), .A2(g2399) );
  AND2_X1 AND2_48( .ZN(g8327), .A1(g3254), .A2(g219) );
  AND2_X1 AND2_49( .ZN(g8328), .A1(g6314), .A2(g225) );
  AND2_X1 AND2_50( .ZN(g8329), .A1(g6232), .A2(g231) );
  AND2_X1 AND2_51( .ZN(g8339), .A1(g6519), .A2(g903) );
  AND2_X1 AND2_52( .ZN(g8340), .A1(g6369), .A2(g909) );
  AND2_X1 AND2_53( .ZN(g8350), .A1(g6574), .A2(g1594) );
  AND2_X1 AND2_54( .ZN(g8385), .A1(g3254), .A2(g228) );
  AND2_X1 AND2_55( .ZN(g8386), .A1(g6314), .A2(g234) );
  AND2_X1 AND2_56( .ZN(g8387), .A1(g6232), .A2(g240) );
  AND2_X1 AND2_57( .ZN(g8394), .A1(g3410), .A2(g906) );
  AND2_X1 AND2_58( .ZN(g8395), .A1(g6519), .A2(g912) );
  AND2_X1 AND2_59( .ZN(g8396), .A1(g6369), .A2(g918) );
  AND2_X1 AND2_60( .ZN(g8406), .A1(g6783), .A2(g1597) );
  AND2_X1 AND2_61( .ZN(g8407), .A1(g6574), .A2(g1603) );
  AND2_X1 AND2_62( .ZN(g8417), .A1(g6838), .A2(g2288) );
  AND2_X1 AND2_63( .ZN(g8431), .A1(g3254), .A2(g237) );
  AND2_X1 AND2_64( .ZN(g8432), .A1(g6314), .A2(g243) );
  AND2_X1 AND2_65( .ZN(g8433), .A1(g6232), .A2(g249) );
  AND2_X1 AND2_66( .ZN(g8437), .A1(g3410), .A2(g915) );
  AND2_X1 AND2_67( .ZN(g8438), .A1(g6519), .A2(g921) );
  AND2_X1 AND2_68( .ZN(g8439), .A1(g6369), .A2(g927) );
  AND2_X1 AND2_69( .ZN(g8446), .A1(g3566), .A2(g1600) );
  AND2_X1 AND2_70( .ZN(g8447), .A1(g6783), .A2(g1606) );
  AND2_X1 AND2_71( .ZN(g8448), .A1(g6574), .A2(g1612) );
  AND2_X1 AND2_72( .ZN(g8458), .A1(g7085), .A2(g2291) );
  AND2_X1 AND2_73( .ZN(g8459), .A1(g6838), .A2(g2297) );
  AND2_X1 AND2_74( .ZN(g8463), .A1(g3254), .A2(g246) );
  AND2_X1 AND2_75( .ZN(g8464), .A1(g6314), .A2(g252) );
  AND2_X1 AND2_76( .ZN(g8465), .A1(g6232), .A2(g258) );
  AND2_X1 AND2_77( .ZN(g8466), .A1(g3410), .A2(g924) );
  AND2_X1 AND2_78( .ZN(g8467), .A1(g6519), .A2(g930) );
  AND2_X1 AND2_79( .ZN(g8468), .A1(g6369), .A2(g936) );
  AND2_X1 AND2_80( .ZN(g8472), .A1(g3566), .A2(g1609) );
  AND2_X1 AND2_81( .ZN(g8473), .A1(g6783), .A2(g1615) );
  AND2_X1 AND2_82( .ZN(g8474), .A1(g6574), .A2(g1621) );
  AND2_X1 AND2_83( .ZN(g8481), .A1(g3722), .A2(g2294) );
  AND2_X1 AND2_84( .ZN(g8482), .A1(g7085), .A2(g2300) );
  AND2_X1 AND2_85( .ZN(g8483), .A1(g6838), .A2(g2306) );
  AND2_X1 AND2_86( .ZN(g8484), .A1(g6232), .A2(g186) );
  AND2_X1 AND2_87( .ZN(g8485), .A1(g3254), .A2(g255) );
  AND2_X1 AND2_88( .ZN(g8486), .A1(g6314), .A2(g261) );
  AND2_X1 AND2_89( .ZN(g8487), .A1(g6232), .A2(g267) );
  AND2_X1 AND2_90( .ZN(g8488), .A1(g3410), .A2(g933) );
  AND2_X1 AND2_91( .ZN(g8489), .A1(g6519), .A2(g939) );
  AND2_X1 AND2_92( .ZN(g8490), .A1(g6369), .A2(g945) );
  AND2_X1 AND2_93( .ZN(g8491), .A1(g3566), .A2(g1618) );
  AND2_X1 AND2_94( .ZN(g8492), .A1(g6783), .A2(g1624) );
  AND2_X1 AND2_95( .ZN(g8493), .A1(g6574), .A2(g1630) );
  AND2_X1 AND2_96( .ZN(g8497), .A1(g3722), .A2(g2303) );
  AND2_X1 AND2_97( .ZN(g8498), .A1(g7085), .A2(g2309) );
  AND2_X1 AND2_98( .ZN(g8499), .A1(g6838), .A2(g2315) );
  AND2_X1 AND2_99( .ZN(g8500), .A1(g6314), .A2(g189) );
  AND2_X1 AND2_100( .ZN(g8501), .A1(g6232), .A2(g195) );
  AND2_X1 AND2_101( .ZN(g8502), .A1(g3254), .A2(g264) );
  AND2_X1 AND2_102( .ZN(g8503), .A1(g6314), .A2(g270) );
  AND2_X1 AND2_103( .ZN(g8504), .A1(g6369), .A2(g873) );
  AND2_X1 AND2_104( .ZN(g8505), .A1(g3410), .A2(g942) );
  AND2_X1 AND2_105( .ZN(g8506), .A1(g6519), .A2(g948) );
  AND2_X1 AND2_106( .ZN(g8507), .A1(g6369), .A2(g954) );
  AND2_X1 AND2_107( .ZN(g8508), .A1(g3566), .A2(g1627) );
  AND2_X1 AND2_108( .ZN(g8509), .A1(g6783), .A2(g1633) );
  AND2_X1 AND2_109( .ZN(g8510), .A1(g6574), .A2(g1639) );
  AND2_X1 AND2_110( .ZN(g8511), .A1(g3722), .A2(g2312) );
  AND2_X1 AND2_111( .ZN(g8512), .A1(g7085), .A2(g2318) );
  AND2_X1 AND2_112( .ZN(g8513), .A1(g6838), .A2(g2324) );
  AND2_X1 AND2_113( .ZN(g8515), .A1(g3254), .A2(g192) );
  AND2_X1 AND2_114( .ZN(g8516), .A1(g6314), .A2(g198) );
  AND2_X1 AND2_115( .ZN(g8517), .A1(g6232), .A2(g204) );
  AND2_X1 AND2_116( .ZN(g8518), .A1(g3254), .A2(g273) );
  AND2_X1 AND2_117( .ZN(g8519), .A1(g6519), .A2(g876) );
  AND2_X1 AND2_118( .ZN(g8520), .A1(g6369), .A2(g882) );
  AND2_X1 AND2_119( .ZN(g8521), .A1(g3410), .A2(g951) );
  AND2_X1 AND2_120( .ZN(g8522), .A1(g6519), .A2(g957) );
  AND2_X1 AND2_121( .ZN(g8523), .A1(g6574), .A2(g1567) );
  AND2_X1 AND2_122( .ZN(g8524), .A1(g3566), .A2(g1636) );
  AND2_X1 AND2_123( .ZN(g8525), .A1(g6783), .A2(g1642) );
  AND2_X1 AND2_124( .ZN(g8526), .A1(g6574), .A2(g1648) );
  AND2_X1 AND2_125( .ZN(g8527), .A1(g3722), .A2(g2321) );
  AND2_X1 AND2_126( .ZN(g8528), .A1(g7085), .A2(g2327) );
  AND2_X2 AND2_127( .ZN(g8529), .A1(g6838), .A2(g2333) );
  AND2_X2 AND2_128( .ZN(g8531), .A1(g3254), .A2(g201) );
  AND2_X1 AND2_129( .ZN(g8532), .A1(g6314), .A2(g207) );
  AND2_X1 AND2_130( .ZN(g8534), .A1(g3410), .A2(g879) );
  AND2_X1 AND2_131( .ZN(g8535), .A1(g6519), .A2(g885) );
  AND2_X1 AND2_132( .ZN(g8536), .A1(g6369), .A2(g891) );
  AND2_X1 AND2_133( .ZN(g8537), .A1(g3410), .A2(g960) );
  AND2_X1 AND2_134( .ZN(g8538), .A1(g6783), .A2(g1570) );
  AND2_X1 AND2_135( .ZN(g8539), .A1(g6574), .A2(g1576) );
  AND2_X1 AND2_136( .ZN(g8540), .A1(g3566), .A2(g1645) );
  AND2_X1 AND2_137( .ZN(g8541), .A1(g6783), .A2(g1651) );
  AND2_X1 AND2_138( .ZN(g8542), .A1(g6838), .A2(g2261) );
  AND2_X1 AND2_139( .ZN(g8543), .A1(g3722), .A2(g2330) );
  AND2_X1 AND2_140( .ZN(g8544), .A1(g7085), .A2(g2336) );
  AND2_X1 AND2_141( .ZN(g8545), .A1(g6838), .A2(g2342) );
  AND2_X1 AND2_142( .ZN(g8546), .A1(g3254), .A2(g210) );
  AND2_X1 AND2_143( .ZN(g8548), .A1(g3410), .A2(g888) );
  AND2_X1 AND2_144( .ZN(g8549), .A1(g6519), .A2(g894) );
  AND2_X1 AND2_145( .ZN(g8551), .A1(g3566), .A2(g1573) );
  AND2_X1 AND2_146( .ZN(g8552), .A1(g6783), .A2(g1579) );
  AND2_X1 AND2_147( .ZN(g8553), .A1(g6574), .A2(g1585) );
  AND2_X1 AND2_148( .ZN(g8554), .A1(g3566), .A2(g1654) );
  AND2_X1 AND2_149( .ZN(g8555), .A1(g7085), .A2(g2264) );
  AND2_X1 AND2_150( .ZN(g8556), .A1(g6838), .A2(g2270) );
  AND2_X1 AND2_151( .ZN(g8557), .A1(g3722), .A2(g2339) );
  AND2_X1 AND2_152( .ZN(g8558), .A1(g7085), .A2(g2345) );
  AND2_X1 AND2_153( .ZN(g8559), .A1(g3410), .A2(g897) );
  AND2_X1 AND2_154( .ZN(g8561), .A1(g3566), .A2(g1582) );
  AND2_X1 AND2_155( .ZN(g8562), .A1(g6783), .A2(g1588) );
  AND2_X1 AND2_156( .ZN(g8564), .A1(g3722), .A2(g2267) );
  AND2_X1 AND2_157( .ZN(g8565), .A1(g7085), .A2(g2273) );
  AND2_X1 AND2_158( .ZN(g8566), .A1(g6838), .A2(g2279) );
  AND2_X1 AND2_159( .ZN(g8567), .A1(g3722), .A2(g2348) );
  AND2_X1 AND2_160( .ZN(g8570), .A1(g3566), .A2(g1591) );
  AND2_X1 AND2_161( .ZN(g8572), .A1(g3722), .A2(g2276) );
  AND2_X1 AND2_162( .ZN(g8573), .A1(g7085), .A2(g2282) );
  AND2_X1 AND2_163( .ZN(g8576), .A1(g3722), .A2(g2285) );
  AND2_X1 AND2_164( .ZN(g8601), .A1(g6643), .A2(g7153) );
  AND2_X1 AND2_165( .ZN(g8612), .A1(g3338), .A2(g6908) );
  AND2_X1 AND2_166( .ZN(g8613), .A1(g6945), .A2(g7349) );
  AND2_X1 AND2_167( .ZN(g8621), .A1(g6486), .A2(g6672) );
  AND2_X1 AND2_168( .ZN(g8625), .A1(g3494), .A2(g7158) );
  AND2_X1 AND2_169( .ZN(g8626), .A1(g7195), .A2(g7479) );
  AND2_X1 AND2_170( .ZN(g8631), .A1(g6751), .A2(g6974) );
  AND2_X1 AND2_171( .ZN(g8635), .A1(g3650), .A2(g7354) );
  AND2_X1 AND2_172( .ZN(g8636), .A1(g7391), .A2(g7535) );
  AND2_X1 AND2_173( .ZN(g8650), .A1(g7053), .A2(g7224) );
  AND2_X1 AND2_174( .ZN(g8654), .A1(g3806), .A2(g7484) );
  AND2_X1 AND2_175( .ZN(g8666), .A1(g7303), .A2(g7420) );
  AND2_X1 AND2_176( .ZN(g8676), .A1(g6643), .A2(g7838) );
  AND2_X1 AND2_177( .ZN(g8687), .A1(g3338), .A2(g7827) );
  AND2_X1 AND2_178( .ZN(g8688), .A1(g6945), .A2(g7858) );
  AND2_X1 AND2_179( .ZN(g8703), .A1(g6486), .A2(g7819) );
  AND2_X1 AND2_180( .ZN(g8704), .A1(g6643), .A2(g7996) );
  AND2_X1 AND2_181( .ZN(g8705), .A1(g3494), .A2(g7842) );
  AND2_X1 AND2_182( .ZN(g8706), .A1(g7195), .A2(g7888) );
  AND2_X1 AND2_183( .ZN(g8717), .A1(g3338), .A2(g7953) );
  AND2_X1 AND2_184( .ZN(g8722), .A1(g6751), .A2(g7830) );
  AND2_X1 AND2_185( .ZN(g8723), .A1(g6945), .A2(g8071) );
  AND2_X1 AND2_186( .ZN(g8724), .A1(g3650), .A2(g7862) );
  AND2_X1 AND2_187( .ZN(g8725), .A1(g7391), .A2(g7912) );
  AND2_X1 AND2_188( .ZN(g8751), .A1(g6486), .A2(g7906) );
  AND2_X1 AND2_189( .ZN(g8755), .A1(g3494), .A2(g8004) );
  AND2_X1 AND2_190( .ZN(g8760), .A1(g7053), .A2(g7845) );
  AND2_X1 AND2_191( .ZN(g8761), .A1(g7195), .A2(g8156) );
  AND2_X1 AND2_192( .ZN(g8762), .A1(g3806), .A2(g7892) );
  AND2_X1 AND2_193( .ZN(g8774), .A1(g6751), .A2(g7958) );
  AND2_X1 AND2_194( .ZN(g8778), .A1(g3650), .A2(g8079) );
  AND2_X2 AND2_195( .ZN(g8783), .A1(g7303), .A2(g7865) );
  AND2_X2 AND2_196( .ZN(g8784), .A1(g7391), .A2(g8242) );
  AND2_X2 AND2_197( .ZN(g8797), .A1(g7053), .A2(g8009) );
  AND2_X1 AND2_198( .ZN(g8801), .A1(g3806), .A2(g8164) );
  AND2_X1 AND2_199( .ZN(g8816), .A1(g7303), .A2(g8084) );
  AND2_X1 AND2_200( .ZN(g8841), .A1(g6486), .A2(g490) );
  AND2_X1 AND2_201( .ZN(g8842), .A1(g6512), .A2(g5508) );
  AND2_X1 AND2_202( .ZN(g8861), .A1(g6643), .A2(g493) );
  AND2_X1 AND2_203( .ZN(g8868), .A1(g6751), .A2(g1177) );
  AND2_X1 AND2_204( .ZN(g8869), .A1(g6776), .A2(g5552) );
  AND2_X1 AND2_205( .ZN(g8892), .A1(g3338), .A2(g496) );
  AND2_X1 AND2_206( .ZN(g8899), .A1(g6945), .A2(g1180) );
  AND2_X1 AND2_207( .ZN(g8906), .A1(g7053), .A2(g1871) );
  AND2_X1 AND2_208( .ZN(g8907), .A1(g7078), .A2(g5598) );
  AND2_X1 AND2_209( .ZN(g8932), .A1(g3494), .A2(g1183) );
  AND2_X1 AND2_210( .ZN(g8939), .A1(g7195), .A2(g1874) );
  AND2_X1 AND2_211( .ZN(g8946), .A1(g7303), .A2(g2565) );
  AND2_X1 AND2_212( .ZN(g8947), .A1(g7328), .A2(g5615) );
  AND2_X1 AND2_213( .ZN(g8972), .A1(g3650), .A2(g1877) );
  AND2_X1 AND2_214( .ZN(g8979), .A1(g7391), .A2(g2568) );
  AND2_X1 AND2_215( .ZN(g9004), .A1(g3806), .A2(g2571) );
  AND2_X1 AND2_216( .ZN(g9009), .A1(g6486), .A2(g565) );
  AND2_X1 AND2_217( .ZN(g9026), .A1(g5438), .A2(g7610) );
  AND2_X1 AND2_218( .ZN(g9033), .A1(g6643), .A2(g567) );
  AND2_X1 AND2_219( .ZN(g9034), .A1(g6751), .A2(g1251) );
  AND2_X1 AND2_220( .ZN(g9047), .A1(g6448), .A2(g7616) );
  AND2_X1 AND2_221( .ZN(g9048), .A1(g3338), .A2(g489) );
  AND2_X1 AND2_222( .ZN(g9049), .A1(g5473), .A2(g7619) );
  AND2_X1 AND2_223( .ZN(g9056), .A1(g6945), .A2(g1253) );
  AND2_X1 AND2_224( .ZN(g9057), .A1(g7053), .A2(g1945) );
  AND2_X1 AND2_225( .ZN(g9061), .A1(g3306), .A2(g7623) );
  AND2_X1 AND2_226( .ZN(g9062), .A1(g5438), .A2(g7626) );
  AND2_X1 AND2_227( .ZN(g9063), .A1(g5438), .A2(g7629) );
  AND2_X1 AND2_228( .ZN(g9064), .A1(g6713), .A2(g7632) );
  AND2_X1 AND2_229( .ZN(g9065), .A1(g3494), .A2(g1176) );
  AND2_X1 AND2_230( .ZN(g9066), .A1(g5512), .A2(g7635) );
  AND2_X1 AND2_231( .ZN(g9073), .A1(g7195), .A2(g1947) );
  AND2_X1 AND2_232( .ZN(g9074), .A1(g7303), .A2(g2639) );
  AND2_X1 AND2_233( .ZN(g9075), .A1(g6448), .A2(g7643) );
  AND2_X1 AND2_234( .ZN(g9076), .A1(g5438), .A2(g7646) );
  AND2_X1 AND2_235( .ZN(g9077), .A1(g6448), .A2(g7649) );
  AND2_X1 AND2_236( .ZN(g9078), .A1(g3462), .A2(g7652) );
  AND2_X1 AND2_237( .ZN(g9079), .A1(g5473), .A2(g7655) );
  AND2_X1 AND2_238( .ZN(g9080), .A1(g5473), .A2(g7658) );
  AND2_X1 AND2_239( .ZN(g9081), .A1(g7015), .A2(g7661) );
  AND2_X1 AND2_240( .ZN(g9082), .A1(g3650), .A2(g1870) );
  AND2_X1 AND2_241( .ZN(g9083), .A1(g5556), .A2(g7664) );
  AND2_X1 AND2_242( .ZN(g9090), .A1(g7391), .A2(g2641) );
  AND2_X1 AND2_243( .ZN(g9091), .A1(g3306), .A2(g7670) );
  AND2_X1 AND2_244( .ZN(g9092), .A1(g6448), .A2(g7673) );
  AND2_X1 AND2_245( .ZN(g9093), .A1(g3306), .A2(g7676) );
  AND2_X1 AND2_246( .ZN(g9094), .A1(g6713), .A2(g7679) );
  AND2_X1 AND2_247( .ZN(g9095), .A1(g5473), .A2(g7682) );
  AND2_X1 AND2_248( .ZN(g9096), .A1(g6713), .A2(g7685) );
  AND2_X1 AND2_249( .ZN(g9097), .A1(g3618), .A2(g7688) );
  AND2_X1 AND2_250( .ZN(g9098), .A1(g5512), .A2(g7691) );
  AND2_X1 AND2_251( .ZN(g9099), .A1(g5512), .A2(g7694) );
  AND2_X1 AND2_252( .ZN(g9100), .A1(g7265), .A2(g7697) );
  AND2_X1 AND2_253( .ZN(g9101), .A1(g3806), .A2(g2564) );
  AND2_X1 AND2_254( .ZN(g9102), .A1(g3306), .A2(g7703) );
  AND2_X1 AND2_255( .ZN(g9103), .A1(g3462), .A2(g7706) );
  AND2_X1 AND2_256( .ZN(g9104), .A1(g6713), .A2(g7709) );
  AND2_X1 AND2_257( .ZN(g9105), .A1(g3462), .A2(g7712) );
  AND2_X1 AND2_258( .ZN(g9106), .A1(g7015), .A2(g7715) );
  AND2_X1 AND2_259( .ZN(g9107), .A1(g5512), .A2(g7718) );
  AND2_X1 AND2_260( .ZN(g9108), .A1(g7015), .A2(g7721) );
  AND2_X1 AND2_261( .ZN(g9109), .A1(g3774), .A2(g7724) );
  AND2_X1 AND2_262( .ZN(g9110), .A1(g5556), .A2(g7727) );
  AND2_X1 AND2_263( .ZN(g9111), .A1(g5556), .A2(g7730) );
  AND2_X1 AND2_264( .ZN(g9112), .A1(g3462), .A2(g7733) );
  AND2_X1 AND2_265( .ZN(g9113), .A1(g3618), .A2(g7736) );
  AND2_X1 AND2_266( .ZN(g9114), .A1(g7015), .A2(g7739) );
  AND2_X1 AND2_267( .ZN(g9115), .A1(g3618), .A2(g7742) );
  AND2_X1 AND2_268( .ZN(g9116), .A1(g7265), .A2(g7745) );
  AND2_X1 AND2_269( .ZN(g9117), .A1(g5556), .A2(g7748) );
  AND2_X1 AND2_270( .ZN(g9118), .A1(g7265), .A2(g7751) );
  AND2_X1 AND2_271( .ZN(g9119), .A1(g5438), .A2(g7754) );
  AND2_X1 AND2_272( .ZN(g9120), .A1(g3618), .A2(g7757) );
  AND2_X1 AND2_273( .ZN(g9121), .A1(g3774), .A2(g7760) );
  AND2_X1 AND2_274( .ZN(g9122), .A1(g7265), .A2(g7763) );
  AND2_X1 AND2_275( .ZN(g9123), .A1(g3774), .A2(g7766) );
  AND2_X1 AND2_276( .ZN(g9124), .A1(g6448), .A2(g7769) );
  AND2_X1 AND2_277( .ZN(g9125), .A1(g5473), .A2(g7776) );
  AND2_X1 AND2_278( .ZN(g9126), .A1(g3774), .A2(g7779) );
  AND2_X1 AND2_279( .ZN(g9127), .A1(g3306), .A2(g7782) );
  AND2_X1 AND2_280( .ZN(g9131), .A1(g6713), .A2(g7785) );
  AND2_X1 AND2_281( .ZN(g9132), .A1(g5512), .A2(g7792) );
  AND2_X1 AND2_282( .ZN(g9133), .A1(g3462), .A2(g7796) );
  AND2_X1 AND2_283( .ZN(g9137), .A1(g7015), .A2(g7799) );
  AND2_X1 AND2_284( .ZN(g9138), .A1(g5556), .A2(g7806) );
  AND2_X1 AND2_285( .ZN(g9139), .A1(g3618), .A2(g7809) );
  AND2_X1 AND2_286( .ZN(g9143), .A1(g7265), .A2(g7812) );
  AND2_X1 AND2_287( .ZN(g9145), .A1(g3774), .A2(g7823) );
  AND2_X1 AND2_288( .ZN(g9241), .A1(g6232), .A2(g7950) );
  AND2_X1 AND2_289( .ZN(g9301), .A1(g6314), .A2(g7990) );
  AND2_X1 AND2_290( .ZN(g9302), .A1(g6232), .A2(g7993) );
  AND2_X1 AND2_291( .ZN(g9319), .A1(g6369), .A2(g8001) );
  AND2_X1 AND2_292( .ZN(g9364), .A1(g3254), .A2(g8053) );
  AND2_X1 AND2_293( .ZN(g9365), .A1(g6314), .A2(g8056) );
  AND2_X1 AND2_294( .ZN(g9366), .A1(g6232), .A2(g8059) );
  AND2_X1 AND2_295( .ZN(g9367), .A1(g6232), .A2(g8062) );
  AND2_X1 AND2_296( .ZN(g9382), .A1(g6519), .A2(g8065) );
  AND2_X1 AND2_297( .ZN(g9383), .A1(g6369), .A2(g8068) );
  AND2_X1 AND2_298( .ZN(g9400), .A1(g6574), .A2(g8076) );
  AND2_X1 AND2_299( .ZN(g9438), .A1(g3254), .A2(g8123) );
  AND2_X1 AND2_300( .ZN(g9439), .A1(g6314), .A2(g8126) );
  AND2_X1 AND2_301( .ZN(g9440), .A1(g6232), .A2(g8129) );
  AND2_X1 AND2_302( .ZN(g9441), .A1(g6314), .A2(g8132) );
  AND2_X1 AND2_303( .ZN(g9442), .A1(g6232), .A2(g8135) );
  AND2_X1 AND2_304( .ZN(g9461), .A1(g3410), .A2(g8138) );
  AND2_X1 AND2_305( .ZN(g9462), .A1(g6519), .A2(g8141) );
  AND2_X1 AND2_306( .ZN(g9463), .A1(g6369), .A2(g8144) );
  AND2_X1 AND2_307( .ZN(g9464), .A1(g6369), .A2(g8147) );
  AND2_X1 AND2_308( .ZN(g9479), .A1(g6783), .A2(g8150) );
  AND2_X1 AND2_309( .ZN(g9480), .A1(g6574), .A2(g8153) );
  AND2_X1 AND2_310( .ZN(g9497), .A1(g6838), .A2(g8161) );
  AND2_X1 AND2_311( .ZN(g9518), .A1(g3254), .A2(g8191) );
  AND2_X1 AND2_312( .ZN(g9519), .A1(g6314), .A2(g8194) );
  AND2_X1 AND2_313( .ZN(g9520), .A1(g6232), .A2(g8197) );
  AND2_X1 AND2_314( .ZN(g9521), .A1(g3254), .A2(g8200) );
  AND2_X2 AND2_315( .ZN(g9522), .A1(g6314), .A2(g8203) );
  AND2_X2 AND2_316( .ZN(g9523), .A1(g6232), .A2(g8206) );
  AND3_X1 AND3_0( .ZN(g9534), .A1(g7772), .A2(g6135), .A3(g538) );
  AND2_X1 AND2_317( .ZN(g9580), .A1(g3410), .A2(g8209) );
  AND2_X1 AND2_318( .ZN(g9581), .A1(g6519), .A2(g8212) );
  AND2_X1 AND2_319( .ZN(g9582), .A1(g6369), .A2(g8215) );
  AND2_X1 AND2_320( .ZN(g9583), .A1(g6519), .A2(g8218) );
  AND2_X1 AND2_321( .ZN(g9584), .A1(g6369), .A2(g8221) );
  AND2_X1 AND2_322( .ZN(g9603), .A1(g3566), .A2(g8224) );
  AND2_X1 AND2_323( .ZN(g9604), .A1(g6783), .A2(g8227) );
  AND2_X1 AND2_324( .ZN(g9605), .A1(g6574), .A2(g8230) );
  AND2_X1 AND2_325( .ZN(g9606), .A1(g6574), .A2(g8233) );
  AND2_X1 AND2_326( .ZN(g9621), .A1(g7085), .A2(g8236) );
  AND2_X1 AND2_327( .ZN(g9622), .A1(g6838), .A2(g8239) );
  AND2_X1 AND2_328( .ZN(g9630), .A1(g3254), .A2(g3922) );
  AND2_X1 AND2_329( .ZN(g9631), .A1(g6314), .A2(g3925) );
  AND2_X1 AND2_330( .ZN(g9632), .A1(g6232), .A2(g3928) );
  AND2_X1 AND2_331( .ZN(g9633), .A1(g3254), .A2(g3931) );
  AND2_X1 AND2_332( .ZN(g9634), .A1(g6314), .A2(g3934) );
  AND2_X1 AND2_333( .ZN(g9635), .A1(g6232), .A2(g3937) );
  AND4_X1 AND4_0( .ZN(II16735), .A1(g5856), .A2(g4338), .A3(g4339), .A4(g5141) );
  AND4_X1 AND4_1( .ZN(II16736), .A1(g5713), .A2(g5958), .A3(g4735), .A4(g4736) );
  AND2_X1 AND2_334( .ZN(g9636), .A1(II16735), .A2(II16736) );
  AND2_X1 AND2_335( .ZN(g9639), .A1(g5438), .A2(g408) );
  AND2_X1 AND2_336( .ZN(g9647), .A1(g6678), .A2(g3942) );
  AND2_X1 AND2_337( .ZN(g9648), .A1(g6678), .A2(g3945) );
  AND2_X1 AND2_338( .ZN(g9660), .A1(g3410), .A2(g3948) );
  AND2_X1 AND2_339( .ZN(g9661), .A1(g6519), .A2(g3951) );
  AND2_X1 AND2_340( .ZN(g9662), .A1(g6369), .A2(g3954) );
  AND2_X1 AND2_341( .ZN(g9663), .A1(g3410), .A2(g3957) );
  AND2_X1 AND2_342( .ZN(g9664), .A1(g6519), .A2(g3960) );
  AND2_X1 AND2_343( .ZN(g9665), .A1(g6369), .A2(g3963) );
  AND3_X1 AND3_1( .ZN(g9676), .A1(g7788), .A2(g6145), .A3(g1224) );
  AND2_X1 AND2_344( .ZN(g9722), .A1(g3566), .A2(g3966) );
  AND2_X1 AND2_345( .ZN(g9723), .A1(g6783), .A2(g3969) );
  AND2_X1 AND2_346( .ZN(g9724), .A1(g6574), .A2(g3972) );
  AND2_X1 AND2_347( .ZN(g9725), .A1(g6783), .A2(g3975) );
  AND2_X1 AND2_348( .ZN(g9726), .A1(g6574), .A2(g3978) );
  AND2_X1 AND2_349( .ZN(g9745), .A1(g3722), .A2(g3981) );
  AND2_X1 AND2_350( .ZN(g9746), .A1(g7085), .A2(g3984) );
  AND2_X1 AND2_351( .ZN(g9747), .A1(g6838), .A2(g3987) );
  AND2_X1 AND2_352( .ZN(g9748), .A1(g6838), .A2(g3990) );
  AND2_X1 AND2_353( .ZN(g9759), .A1(g3254), .A2(g4000) );
  AND2_X1 AND2_354( .ZN(g9760), .A1(g6314), .A2(g4003) );
  AND2_X1 AND2_355( .ZN(g9761), .A1(g6232), .A2(g4006) );
  AND2_X1 AND2_356( .ZN(g9762), .A1(g3254), .A2(g4009) );
  AND2_X1 AND2_357( .ZN(g9763), .A1(g6314), .A2(g4012) );
  AND2_X1 AND2_358( .ZN(g9764), .A1(g6448), .A2(g411) );
  AND2_X1 AND2_359( .ZN(g9765), .A1(g5438), .A2(g417) );
  AND2_X1 AND2_360( .ZN(g9766), .A1(g5438), .A2(g4017) );
  AND2_X1 AND2_361( .ZN(g9773), .A1(g6912), .A2(g4020) );
  AND2_X1 AND2_362( .ZN(g9774), .A1(g6678), .A2(g4023) );
  AND2_X1 AND2_363( .ZN(g9775), .A1(g6912), .A2(g4026) );
  AND2_X1 AND2_364( .ZN(g9776), .A1(g3410), .A2(g4029) );
  AND2_X1 AND2_365( .ZN(g9777), .A1(g6519), .A2(g4032) );
  AND2_X1 AND2_366( .ZN(g9778), .A1(g6369), .A2(g4035) );
  AND2_X1 AND2_367( .ZN(g9779), .A1(g3410), .A2(g4038) );
  AND2_X1 AND2_368( .ZN(g9780), .A1(g6519), .A2(g4041) );
  AND2_X1 AND2_369( .ZN(g9781), .A1(g6369), .A2(g4044) );
  AND4_X1 AND4_2( .ZN(II16826), .A1(g5903), .A2(g4507), .A3(g4508), .A4(g5234) );
  AND4_X1 AND4_3( .ZN(II16827), .A1(g5771), .A2(g5987), .A3(g4911), .A4(g4912) );
  AND2_X1 AND2_370( .ZN(g9782), .A1(II16826), .A2(II16827) );
  AND2_X1 AND2_371( .ZN(g9785), .A1(g5473), .A2(g1095) );
  AND2_X1 AND2_372( .ZN(g9793), .A1(g6980), .A2(g4049) );
  AND2_X1 AND2_373( .ZN(g9794), .A1(g6980), .A2(g4052) );
  AND2_X1 AND2_374( .ZN(g9806), .A1(g3566), .A2(g4055) );
  AND2_X1 AND2_375( .ZN(g9807), .A1(g6783), .A2(g4058) );
  AND2_X1 AND2_376( .ZN(g9808), .A1(g6574), .A2(g4061) );
  AND2_X1 AND2_377( .ZN(g9809), .A1(g3566), .A2(g4064) );
  AND2_X1 AND2_378( .ZN(g9810), .A1(g6783), .A2(g4067) );
  AND2_X1 AND2_379( .ZN(g9811), .A1(g6574), .A2(g4070) );
  AND3_X1 AND3_2( .ZN(g9822), .A1(g7802), .A2(g6166), .A3(g1918) );
  AND2_X1 AND2_380( .ZN(g9868), .A1(g3722), .A2(g4073) );
  AND2_X1 AND2_381( .ZN(g9869), .A1(g7085), .A2(g4076) );
  AND2_X1 AND2_382( .ZN(g9870), .A1(g6838), .A2(g4079) );
  AND2_X1 AND2_383( .ZN(g9871), .A1(g7085), .A2(g4082) );
  AND2_X1 AND2_384( .ZN(g9872), .A1(g6838), .A2(g4085) );
  AND2_X1 AND2_385( .ZN(g9887), .A1(g6232), .A2(g4095) );
  AND2_X1 AND2_386( .ZN(g9888), .A1(g3254), .A2(g4098) );
  AND2_X1 AND2_387( .ZN(g9889), .A1(g6314), .A2(g4101) );
  AND2_X1 AND2_388( .ZN(g9890), .A1(g6232), .A2(g4104) );
  AND2_X1 AND2_389( .ZN(g9891), .A1(g3254), .A2(g4107) );
  AND2_X1 AND2_390( .ZN(g9892), .A1(g3306), .A2(g414) );
  AND2_X1 AND2_391( .ZN(g9893), .A1(g6448), .A2(g420) );
  AND2_X1 AND2_392( .ZN(g9894), .A1(g6448), .A2(g4112) );
  AND2_X1 AND2_393( .ZN(g9901), .A1(g3366), .A2(g4115) );
  AND2_X1 AND2_394( .ZN(g9902), .A1(g6912), .A2(g4118) );
  AND2_X1 AND2_395( .ZN(g9903), .A1(g6678), .A2(g4121) );
  AND2_X1 AND2_396( .ZN(g9904), .A1(g3366), .A2(g4124) );
  AND2_X1 AND2_397( .ZN(g9905), .A1(g3410), .A2(g4127) );
  AND2_X1 AND2_398( .ZN(g9906), .A1(g6519), .A2(g4130) );
  AND2_X1 AND2_399( .ZN(g9907), .A1(g6369), .A2(g4133) );
  AND2_X1 AND2_400( .ZN(g9908), .A1(g3410), .A2(g4136) );
  AND2_X1 AND2_401( .ZN(g9909), .A1(g6519), .A2(g4139) );
  AND2_X1 AND2_402( .ZN(g9910), .A1(g6713), .A2(g1098) );
  AND2_X1 AND2_403( .ZN(g9911), .A1(g5473), .A2(g1104) );
  AND2_X1 AND2_404( .ZN(g9912), .A1(g5473), .A2(g4144) );
  AND2_X1 AND2_405( .ZN(g9919), .A1(g7162), .A2(g4147) );
  AND2_X1 AND2_406( .ZN(g9920), .A1(g6980), .A2(g4150) );
  AND2_X1 AND2_407( .ZN(g9921), .A1(g7162), .A2(g4153) );
  AND2_X1 AND2_408( .ZN(g9922), .A1(g3566), .A2(g4156) );
  AND2_X2 AND2_409( .ZN(g9923), .A1(g6783), .A2(g4159) );
  AND2_X2 AND2_410( .ZN(g9924), .A1(g6574), .A2(g4162) );
  AND2_X1 AND2_411( .ZN(g9925), .A1(g3566), .A2(g4165) );
  AND2_X1 AND2_412( .ZN(g9926), .A1(g6783), .A2(g4168) );
  AND2_X1 AND2_413( .ZN(g9927), .A1(g6574), .A2(g4171) );
  AND4_X1 AND4_4( .ZN(II16930), .A1(g5942), .A2(g4683), .A3(g4684), .A4(g5297) );
  AND4_X1 AND4_5( .ZN(II16931), .A1(g5830), .A2(g6024), .A3(g5070), .A4(g5071) );
  AND2_X1 AND2_414( .ZN(g9928), .A1(II16930), .A2(II16931) );
  AND2_X1 AND2_415( .ZN(g9931), .A1(g5512), .A2(g1789) );
  AND2_X1 AND2_416( .ZN(g9939), .A1(g7230), .A2(g4176) );
  AND2_X1 AND2_417( .ZN(g9940), .A1(g7230), .A2(g4179) );
  AND2_X1 AND2_418( .ZN(g9952), .A1(g3722), .A2(g4182) );
  AND2_X1 AND2_419( .ZN(g9953), .A1(g7085), .A2(g4185) );
  AND2_X1 AND2_420( .ZN(g9954), .A1(g6838), .A2(g4188) );
  AND2_X1 AND2_421( .ZN(g9955), .A1(g3722), .A2(g4191) );
  AND2_X1 AND2_422( .ZN(g9956), .A1(g7085), .A2(g4194) );
  AND2_X1 AND2_423( .ZN(g9957), .A1(g6838), .A2(g4197) );
  AND3_X1 AND3_3( .ZN(g9968), .A1(g7815), .A2(g6193), .A3(g2612) );
  AND2_X1 AND2_424( .ZN(g10007), .A1(g6314), .A2(g4205) );
  AND2_X1 AND2_425( .ZN(g10008), .A1(g6232), .A2(g4208) );
  AND2_X1 AND2_426( .ZN(g10009), .A1(g3254), .A2(g4211) );
  AND2_X1 AND2_427( .ZN(g10010), .A1(g6314), .A2(g4214) );
  AND2_X1 AND2_428( .ZN(g10011), .A1(g5438), .A2(g4217) );
  AND2_X1 AND2_429( .ZN(g10012), .A1(g3306), .A2(g423) );
  AND2_X1 AND2_430( .ZN(g10013), .A1(g3306), .A2(g4221) );
  AND2_X1 AND2_431( .ZN(g10014), .A1(g5438), .A2(g429) );
  AND2_X1 AND2_432( .ZN(g10024), .A1(g3398), .A2(g6912) );
  AND2_X1 AND2_433( .ZN(g10035), .A1(g3366), .A2(g4225) );
  AND2_X1 AND2_434( .ZN(g10036), .A1(g6912), .A2(g4228) );
  AND2_X1 AND2_435( .ZN(g10037), .A1(g6678), .A2(g4231) );
  AND2_X1 AND2_436( .ZN(g10041), .A1(g6369), .A2(g4234) );
  AND2_X1 AND2_437( .ZN(g10042), .A1(g3410), .A2(g4237) );
  AND2_X1 AND2_438( .ZN(g10043), .A1(g6519), .A2(g4240) );
  AND2_X1 AND2_439( .ZN(g10044), .A1(g6369), .A2(g4243) );
  AND2_X1 AND2_440( .ZN(g10045), .A1(g3410), .A2(g4246) );
  AND2_X1 AND2_441( .ZN(g10046), .A1(g3462), .A2(g1101) );
  AND2_X1 AND2_442( .ZN(g10047), .A1(g6713), .A2(g1107) );
  AND2_X1 AND2_443( .ZN(g10048), .A1(g6713), .A2(g4251) );
  AND2_X1 AND2_444( .ZN(g10055), .A1(g3522), .A2(g4254) );
  AND2_X1 AND2_445( .ZN(g10056), .A1(g7162), .A2(g4257) );
  AND2_X1 AND2_446( .ZN(g10057), .A1(g6980), .A2(g4260) );
  AND2_X1 AND2_447( .ZN(g10058), .A1(g3522), .A2(g4263) );
  AND2_X1 AND2_448( .ZN(g10059), .A1(g3566), .A2(g4266) );
  AND2_X1 AND2_449( .ZN(g10060), .A1(g6783), .A2(g4269) );
  AND2_X1 AND2_450( .ZN(g10061), .A1(g6574), .A2(g4272) );
  AND2_X1 AND2_451( .ZN(g10062), .A1(g3566), .A2(g4275) );
  AND2_X1 AND2_452( .ZN(g10063), .A1(g6783), .A2(g4278) );
  AND2_X1 AND2_453( .ZN(g10064), .A1(g7015), .A2(g1792) );
  AND2_X1 AND2_454( .ZN(g10065), .A1(g5512), .A2(g1798) );
  AND2_X1 AND2_455( .ZN(g10066), .A1(g5512), .A2(g4283) );
  AND2_X1 AND2_456( .ZN(g10073), .A1(g7358), .A2(g4286) );
  AND2_X1 AND2_457( .ZN(g10074), .A1(g7230), .A2(g4289) );
  AND2_X1 AND2_458( .ZN(g10075), .A1(g7358), .A2(g4292) );
  AND2_X1 AND2_459( .ZN(g10076), .A1(g3722), .A2(g4295) );
  AND2_X1 AND2_460( .ZN(g10077), .A1(g7085), .A2(g4298) );
  AND2_X1 AND2_461( .ZN(g10078), .A1(g6838), .A2(g4301) );
  AND2_X1 AND2_462( .ZN(g10079), .A1(g3722), .A2(g4304) );
  AND2_X1 AND2_463( .ZN(g10080), .A1(g7085), .A2(g4307) );
  AND2_X1 AND2_464( .ZN(g10081), .A1(g6838), .A2(g4310) );
  AND4_X1 AND4_6( .ZN(II17042), .A1(g5976), .A2(g4860), .A3(g4861), .A4(g5334) );
  AND4_X1 AND4_7( .ZN(II17043), .A1(g5886), .A2(g6040), .A3(g5199), .A4(g5200) );
  AND2_X1 AND2_465( .ZN(g10082), .A1(II17042), .A2(II17043) );
  AND2_X1 AND2_466( .ZN(g10085), .A1(g5556), .A2(g2483) );
  AND2_X1 AND2_467( .ZN(g10093), .A1(g7426), .A2(g4315) );
  AND2_X1 AND2_468( .ZN(g10094), .A1(g7426), .A2(g4318) );
  AND2_X1 AND2_469( .ZN(g10101), .A1(g3254), .A2(g4329) );
  AND2_X1 AND2_470( .ZN(g10102), .A1(g6314), .A2(g4332) );
  AND2_X1 AND2_471( .ZN(g10103), .A1(g3254), .A2(g4335) );
  AND2_X1 AND2_472( .ZN(g10104), .A1(g6448), .A2(g4340) );
  AND2_X1 AND2_473( .ZN(g10105), .A1(g5438), .A2(g4343) );
  AND2_X1 AND2_474( .ZN(g10106), .A1(g6448), .A2(g432) );
  AND2_X1 AND2_475( .ZN(g10107), .A1(g5438), .A2(g438) );
  AND2_X1 AND2_476( .ZN(g10108), .A1(g6486), .A2(g569) );
  AND2_X1 AND2_477( .ZN(g10112), .A1(g3366), .A2(g4348) );
  AND2_X1 AND2_478( .ZN(g10113), .A1(g6912), .A2(g4351) );
  AND2_X1 AND2_479( .ZN(g10114), .A1(g6678), .A2(g4354) );
  AND2_X1 AND2_480( .ZN(g10115), .A1(g6678), .A2(g4357) );
  AND2_X1 AND2_481( .ZN(g10116), .A1(g6519), .A2(g4360) );
  AND2_X1 AND2_482( .ZN(g10117), .A1(g6369), .A2(g4363) );
  AND2_X1 AND2_483( .ZN(g10118), .A1(g3410), .A2(g4366) );
  AND2_X1 AND2_484( .ZN(g10119), .A1(g6519), .A2(g4369) );
  AND2_X1 AND2_485( .ZN(g10120), .A1(g5473), .A2(g4372) );
  AND2_X1 AND2_486( .ZN(g10121), .A1(g3462), .A2(g1110) );
  AND2_X1 AND2_487( .ZN(g10122), .A1(g3462), .A2(g4376) );
  AND2_X1 AND2_488( .ZN(g10123), .A1(g5473), .A2(g1116) );
  AND2_X1 AND2_489( .ZN(g10133), .A1(g3554), .A2(g7162) );
  AND2_X1 AND2_490( .ZN(g10144), .A1(g3522), .A2(g4380) );
  AND2_X1 AND2_491( .ZN(g10145), .A1(g7162), .A2(g4383) );
  AND2_X1 AND2_492( .ZN(g10146), .A1(g6980), .A2(g4386) );
  AND2_X1 AND2_493( .ZN(g10150), .A1(g6574), .A2(g4389) );
  AND2_X1 AND2_494( .ZN(g10151), .A1(g3566), .A2(g4392) );
  AND2_X1 AND2_495( .ZN(g10152), .A1(g6783), .A2(g4395) );
  AND2_X1 AND2_496( .ZN(g10153), .A1(g6574), .A2(g4398) );
  AND2_X1 AND2_497( .ZN(g10154), .A1(g3566), .A2(g4401) );
  AND2_X1 AND2_498( .ZN(g10155), .A1(g3618), .A2(g1795) );
  AND2_X1 AND2_499( .ZN(g10156), .A1(g7015), .A2(g1801) );
  AND2_X1 AND2_500( .ZN(g10157), .A1(g7015), .A2(g4406) );
  AND2_X1 AND2_501( .ZN(g10164), .A1(g3678), .A2(g4409) );
  AND2_X1 AND2_502( .ZN(g10165), .A1(g7358), .A2(g4412) );
  AND2_X1 AND2_503( .ZN(g10166), .A1(g7230), .A2(g4415) );
  AND2_X1 AND2_504( .ZN(g10167), .A1(g3678), .A2(g4418) );
  AND2_X1 AND2_505( .ZN(g10168), .A1(g3722), .A2(g4421) );
  AND2_X1 AND2_506( .ZN(g10169), .A1(g7085), .A2(g4424) );
  AND2_X1 AND2_507( .ZN(g10170), .A1(g6838), .A2(g4427) );
  AND2_X1 AND2_508( .ZN(g10171), .A1(g3722), .A2(g4430) );
  AND2_X1 AND2_509( .ZN(g10172), .A1(g7085), .A2(g4433) );
  AND2_X1 AND2_510( .ZN(g10173), .A1(g7265), .A2(g2486) );
  AND2_X1 AND2_511( .ZN(g10174), .A1(g5556), .A2(g2492) );
  AND2_X1 AND2_512( .ZN(g10175), .A1(g5556), .A2(g4438) );
  AND2_X1 AND2_513( .ZN(g10182), .A1(g7488), .A2(g4441) );
  AND2_X1 AND2_514( .ZN(g10183), .A1(g7426), .A2(g4444) );
  AND2_X1 AND2_515( .ZN(g10184), .A1(g7488), .A2(g4447) );
  AND4_X1 AND4_8( .ZN(II17156), .A1(g6898), .A2(g2998), .A3(g6901), .A4(g3002) );
  AND4_X1 AND4_9( .ZN(g10186), .A1(g3013), .A2(g7466), .A3(g3024), .A4(II17156) );
  AND2_X1 AND2_516( .ZN(g10192), .A1(g3254), .A2(g4453) );
  AND2_X1 AND2_517( .ZN(g10193), .A1(g3306), .A2(g4465) );
  AND2_X1 AND2_518( .ZN(g10194), .A1(g6448), .A2(g4468) );
  AND2_X1 AND2_519( .ZN(g10195), .A1(g5438), .A2(g4471) );
  AND2_X1 AND2_520( .ZN(g10196), .A1(g3306), .A2(g435) );
  AND2_X1 AND2_521( .ZN(g10197), .A1(g6448), .A2(g441) );
  AND2_X1 AND2_522( .ZN(g10198), .A1(g6643), .A2(g571) );
  AND2_X1 AND2_523( .ZN(g10199), .A1(g6486), .A2(g4476) );
  AND2_X1 AND2_524( .ZN(g10200), .A1(g6486), .A2(g587) );
  AND2_X1 AND2_525( .ZN(g10201), .A1(g3366), .A2(g4480) );
  AND2_X1 AND2_526( .ZN(g10202), .A1(g6912), .A2(g4483) );
  AND2_X1 AND2_527( .ZN(g10203), .A1(g6678), .A2(g4486) );
  AND2_X1 AND2_528( .ZN(g10204), .A1(g6912), .A2(g4489) );
  AND2_X1 AND2_529( .ZN(g10205), .A1(g6678), .A2(g4492) );
  AND2_X1 AND2_530( .ZN(g10206), .A1(g3410), .A2(g4498) );
  AND2_X1 AND2_531( .ZN(g10207), .A1(g6519), .A2(g4501) );
  AND2_X1 AND2_532( .ZN(g10208), .A1(g3410), .A2(g4504) );
  AND2_X1 AND2_533( .ZN(g10209), .A1(g6713), .A2(g4509) );
  AND2_X1 AND2_534( .ZN(g10210), .A1(g5473), .A2(g4512) );
  AND2_X1 AND2_535( .ZN(g10211), .A1(g6713), .A2(g1119) );
  AND2_X1 AND2_536( .ZN(g10212), .A1(g5473), .A2(g1125) );
  AND2_X1 AND2_537( .ZN(g10213), .A1(g6751), .A2(g1255) );
  AND2_X1 AND2_538( .ZN(g10217), .A1(g3522), .A2(g4517) );
  AND2_X1 AND2_539( .ZN(g10218), .A1(g7162), .A2(g4520) );
  AND2_X1 AND2_540( .ZN(g10219), .A1(g6980), .A2(g4523) );
  AND2_X1 AND2_541( .ZN(g10220), .A1(g6980), .A2(g4526) );
  AND2_X2 AND2_542( .ZN(g10221), .A1(g6783), .A2(g4529) );
  AND2_X2 AND2_543( .ZN(g10222), .A1(g6574), .A2(g4532) );
  AND2_X1 AND2_544( .ZN(g10223), .A1(g3566), .A2(g4535) );
  AND2_X1 AND2_545( .ZN(g10224), .A1(g6783), .A2(g4538) );
  AND2_X1 AND2_546( .ZN(g10225), .A1(g5512), .A2(g4541) );
  AND2_X1 AND2_547( .ZN(g10226), .A1(g3618), .A2(g1804) );
  AND2_X1 AND2_548( .ZN(g10227), .A1(g3618), .A2(g4545) );
  AND2_X1 AND2_549( .ZN(g10228), .A1(g5512), .A2(g1810) );
  AND2_X1 AND2_550( .ZN(g10238), .A1(g3710), .A2(g7358) );
  AND2_X1 AND2_551( .ZN(g10249), .A1(g3678), .A2(g4549) );
  AND2_X1 AND2_552( .ZN(g10250), .A1(g7358), .A2(g4552) );
  AND2_X1 AND2_553( .ZN(g10251), .A1(g7230), .A2(g4555) );
  AND2_X1 AND2_554( .ZN(g10255), .A1(g6838), .A2(g4558) );
  AND2_X1 AND2_555( .ZN(g10256), .A1(g3722), .A2(g4561) );
  AND2_X1 AND2_556( .ZN(g10257), .A1(g7085), .A2(g4564) );
  AND2_X1 AND2_557( .ZN(g10258), .A1(g6838), .A2(g4567) );
  AND2_X1 AND2_558( .ZN(g10259), .A1(g3722), .A2(g4570) );
  AND2_X1 AND2_559( .ZN(g10260), .A1(g3774), .A2(g2489) );
  AND2_X1 AND2_560( .ZN(g10261), .A1(g7265), .A2(g2495) );
  AND2_X1 AND2_561( .ZN(g10262), .A1(g7265), .A2(g4575) );
  AND2_X1 AND2_562( .ZN(g10269), .A1(g3834), .A2(g4578) );
  AND2_X1 AND2_563( .ZN(g10270), .A1(g7488), .A2(g4581) );
  AND2_X1 AND2_564( .ZN(g10271), .A1(g7426), .A2(g4584) );
  AND2_X1 AND2_565( .ZN(g10272), .A1(g3834), .A2(g4587) );
  AND2_X1 AND2_566( .ZN(g10279), .A1(g3306), .A2(g4592) );
  AND2_X1 AND2_567( .ZN(g10280), .A1(g6448), .A2(g4595) );
  AND2_X1 AND2_568( .ZN(g10281), .A1(g5438), .A2(g4598) );
  AND2_X1 AND2_569( .ZN(g10282), .A1(g3306), .A2(g444) );
  AND2_X1 AND2_570( .ZN(g10283), .A1(g3338), .A2(g573) );
  AND2_X1 AND2_571( .ZN(g10284), .A1(g6643), .A2(g4603) );
  AND2_X1 AND2_572( .ZN(g10285), .A1(g6486), .A2(g4606) );
  AND2_X1 AND2_573( .ZN(g10286), .A1(g6643), .A2(g590) );
  AND2_X1 AND2_574( .ZN(g10287), .A1(g6486), .A2(g596) );
  AND2_X1 AND2_575( .ZN(g10288), .A1(g3366), .A2(g4611) );
  AND2_X1 AND2_576( .ZN(g10289), .A1(g6912), .A2(g4614) );
  AND2_X1 AND2_577( .ZN(g10290), .A1(g6678), .A2(g4617) );
  AND2_X1 AND2_578( .ZN(g10291), .A1(g3366), .A2(g4620) );
  AND2_X1 AND2_579( .ZN(g10292), .A1(g6912), .A2(g4623) );
  AND2_X1 AND2_580( .ZN(g10293), .A1(g6678), .A2(g4626) );
  AND2_X1 AND2_581( .ZN(g10294), .A1(g3410), .A2(g4629) );
  AND2_X1 AND2_582( .ZN(g10295), .A1(g3462), .A2(g4641) );
  AND2_X1 AND2_583( .ZN(g10296), .A1(g6713), .A2(g4644) );
  AND2_X1 AND2_584( .ZN(g10297), .A1(g5473), .A2(g4647) );
  AND2_X1 AND2_585( .ZN(g10298), .A1(g3462), .A2(g1122) );
  AND2_X1 AND2_586( .ZN(g10299), .A1(g6713), .A2(g1128) );
  AND2_X1 AND2_587( .ZN(g10300), .A1(g6945), .A2(g1257) );
  AND2_X1 AND2_588( .ZN(g10301), .A1(g6751), .A2(g4652) );
  AND2_X1 AND2_589( .ZN(g10302), .A1(g6751), .A2(g1273) );
  AND2_X1 AND2_590( .ZN(g10303), .A1(g3522), .A2(g4656) );
  AND2_X1 AND2_591( .ZN(g10304), .A1(g7162), .A2(g4659) );
  AND2_X1 AND2_592( .ZN(g10305), .A1(g6980), .A2(g4662) );
  AND2_X1 AND2_593( .ZN(g10306), .A1(g7162), .A2(g4665) );
  AND2_X1 AND2_594( .ZN(g10307), .A1(g6980), .A2(g4668) );
  AND2_X1 AND2_595( .ZN(g10308), .A1(g3566), .A2(g4674) );
  AND2_X1 AND2_596( .ZN(g10309), .A1(g6783), .A2(g4677) );
  AND2_X1 AND2_597( .ZN(g10310), .A1(g3566), .A2(g4680) );
  AND2_X1 AND2_598( .ZN(g10311), .A1(g7015), .A2(g4685) );
  AND2_X1 AND2_599( .ZN(g10312), .A1(g5512), .A2(g4688) );
  AND2_X1 AND2_600( .ZN(g10313), .A1(g7015), .A2(g1813) );
  AND2_X1 AND2_601( .ZN(g10314), .A1(g5512), .A2(g1819) );
  AND2_X1 AND2_602( .ZN(g10315), .A1(g7053), .A2(g1949) );
  AND2_X1 AND2_603( .ZN(g10319), .A1(g3678), .A2(g4693) );
  AND2_X1 AND2_604( .ZN(g10320), .A1(g7358), .A2(g4696) );
  AND2_X1 AND2_605( .ZN(g10321), .A1(g7230), .A2(g4699) );
  AND2_X1 AND2_606( .ZN(g10322), .A1(g7230), .A2(g4702) );
  AND2_X1 AND2_607( .ZN(g10323), .A1(g7085), .A2(g4705) );
  AND2_X1 AND2_608( .ZN(g10324), .A1(g6838), .A2(g4708) );
  AND2_X1 AND2_609( .ZN(g10325), .A1(g3722), .A2(g4711) );
  AND2_X1 AND2_610( .ZN(g10326), .A1(g7085), .A2(g4714) );
  AND2_X1 AND2_611( .ZN(g10327), .A1(g5556), .A2(g4717) );
  AND2_X1 AND2_612( .ZN(g10328), .A1(g3774), .A2(g2498) );
  AND2_X1 AND2_613( .ZN(g10329), .A1(g3774), .A2(g4721) );
  AND2_X1 AND2_614( .ZN(g10330), .A1(g5556), .A2(g2504) );
  AND2_X1 AND2_615( .ZN(g10340), .A1(g3866), .A2(g7488) );
  AND2_X1 AND2_616( .ZN(g10351), .A1(g3834), .A2(g4725) );
  AND2_X1 AND2_617( .ZN(g10352), .A1(g7488), .A2(g4728) );
  AND2_X1 AND2_618( .ZN(g10353), .A1(g7426), .A2(g4731) );
  AND2_X1 AND2_619( .ZN(g10360), .A1(g3306), .A2(g4737) );
  AND2_X1 AND2_620( .ZN(g10361), .A1(g6448), .A2(g4740) );
  AND2_X1 AND2_621( .ZN(g10362), .A1(g3338), .A2(g4743) );
  AND2_X1 AND2_622( .ZN(g10363), .A1(g6643), .A2(g4746) );
  AND2_X1 AND2_623( .ZN(g10364), .A1(g6486), .A2(g4749) );
  AND2_X1 AND2_624( .ZN(g10365), .A1(g3338), .A2(g593) );
  AND2_X1 AND2_625( .ZN(g10366), .A1(g6643), .A2(g599) );
  AND2_X1 AND2_626( .ZN(g10367), .A1(g3366), .A2(g4754) );
  AND2_X1 AND2_627( .ZN(g10368), .A1(g6912), .A2(g4757) );
  AND2_X1 AND2_628( .ZN(g10369), .A1(g6678), .A2(g4760) );
  AND2_X1 AND2_629( .ZN(g10370), .A1(g3366), .A2(g4763) );
  AND2_X1 AND2_630( .ZN(g10371), .A1(g6912), .A2(g4766) );
  AND2_X1 AND2_631( .ZN(g10372), .A1(g3462), .A2(g4769) );
  AND2_X1 AND2_632( .ZN(g10373), .A1(g6713), .A2(g4772) );
  AND2_X1 AND2_633( .ZN(g10374), .A1(g5473), .A2(g4775) );
  AND2_X1 AND2_634( .ZN(g10375), .A1(g3462), .A2(g1131) );
  AND2_X1 AND2_635( .ZN(g10376), .A1(g3494), .A2(g1259) );
  AND2_X1 AND2_636( .ZN(g10377), .A1(g6945), .A2(g4780) );
  AND2_X1 AND2_637( .ZN(g10378), .A1(g6751), .A2(g4783) );
  AND2_X1 AND2_638( .ZN(g10379), .A1(g6945), .A2(g1276) );
  AND2_X1 AND2_639( .ZN(g10380), .A1(g6751), .A2(g1282) );
  AND2_X1 AND2_640( .ZN(g10381), .A1(g3522), .A2(g4788) );
  AND2_X1 AND2_641( .ZN(g10382), .A1(g7162), .A2(g4791) );
  AND2_X1 AND2_642( .ZN(g10383), .A1(g6980), .A2(g4794) );
  AND2_X1 AND2_643( .ZN(g10384), .A1(g3522), .A2(g4797) );
  AND2_X2 AND2_644( .ZN(g10385), .A1(g7162), .A2(g4800) );
  AND2_X2 AND2_645( .ZN(g10386), .A1(g6980), .A2(g4803) );
  AND2_X1 AND2_646( .ZN(g10387), .A1(g3566), .A2(g4806) );
  AND2_X1 AND2_647( .ZN(g10388), .A1(g3618), .A2(g4818) );
  AND2_X1 AND2_648( .ZN(g10389), .A1(g7015), .A2(g4821) );
  AND2_X1 AND2_649( .ZN(g10390), .A1(g5512), .A2(g4824) );
  AND2_X1 AND2_650( .ZN(g10391), .A1(g3618), .A2(g1816) );
  AND2_X1 AND2_651( .ZN(g10392), .A1(g7015), .A2(g1822) );
  AND2_X1 AND2_652( .ZN(g10393), .A1(g7195), .A2(g1951) );
  AND2_X1 AND2_653( .ZN(g10394), .A1(g7053), .A2(g4829) );
  AND2_X1 AND2_654( .ZN(g10395), .A1(g7053), .A2(g1967) );
  AND2_X1 AND2_655( .ZN(g10396), .A1(g3678), .A2(g4833) );
  AND2_X1 AND2_656( .ZN(g10397), .A1(g7358), .A2(g4836) );
  AND2_X1 AND2_657( .ZN(g10398), .A1(g7230), .A2(g4839) );
  AND2_X1 AND2_658( .ZN(g10399), .A1(g7358), .A2(g4842) );
  AND2_X1 AND2_659( .ZN(g10400), .A1(g7230), .A2(g4845) );
  AND2_X1 AND2_660( .ZN(g10401), .A1(g3722), .A2(g4851) );
  AND2_X1 AND2_661( .ZN(g10402), .A1(g7085), .A2(g4854) );
  AND2_X1 AND2_662( .ZN(g10403), .A1(g3722), .A2(g4857) );
  AND2_X1 AND2_663( .ZN(g10404), .A1(g7265), .A2(g4862) );
  AND2_X1 AND2_664( .ZN(g10405), .A1(g5556), .A2(g4865) );
  AND2_X1 AND2_665( .ZN(g10406), .A1(g7265), .A2(g2507) );
  AND2_X1 AND2_666( .ZN(g10407), .A1(g5556), .A2(g2513) );
  AND2_X1 AND2_667( .ZN(g10408), .A1(g7303), .A2(g2643) );
  AND2_X1 AND2_668( .ZN(g10412), .A1(g3834), .A2(g4870) );
  AND2_X1 AND2_669( .ZN(g10413), .A1(g7488), .A2(g4873) );
  AND2_X1 AND2_670( .ZN(g10414), .A1(g7426), .A2(g4876) );
  AND2_X1 AND2_671( .ZN(g10415), .A1(g7426), .A2(g4879) );
  AND2_X1 AND2_672( .ZN(g10422), .A1(g3306), .A2(g4882) );
  AND2_X1 AND2_673( .ZN(g10423), .A1(g5438), .A2(g4885) );
  AND2_X1 AND2_674( .ZN(g10430), .A1(g3338), .A2(g4888) );
  AND2_X1 AND2_675( .ZN(g10431), .A1(g6643), .A2(g4891) );
  AND2_X1 AND2_676( .ZN(g10432), .A1(g6486), .A2(g4894) );
  AND2_X1 AND2_677( .ZN(g10433), .A1(g3338), .A2(g602) );
  AND2_X1 AND2_678( .ZN(g10434), .A1(g6486), .A2(g605) );
  AND2_X1 AND2_679( .ZN(g10435), .A1(g3366), .A2(g4899) );
  AND2_X1 AND2_680( .ZN(g10436), .A1(g6912), .A2(g4902) );
  AND2_X1 AND2_681( .ZN(g10437), .A1(g6678), .A2(g4905) );
  AND2_X1 AND2_682( .ZN(g10438), .A1(g3366), .A2(g4908) );
  AND2_X1 AND2_683( .ZN(g10439), .A1(g3462), .A2(g4913) );
  AND2_X1 AND2_684( .ZN(g10440), .A1(g6713), .A2(g4916) );
  AND2_X1 AND2_685( .ZN(g10441), .A1(g3494), .A2(g4919) );
  AND2_X1 AND2_686( .ZN(g10442), .A1(g6945), .A2(g4922) );
  AND2_X1 AND2_687( .ZN(g10443), .A1(g6751), .A2(g4925) );
  AND2_X1 AND2_688( .ZN(g10444), .A1(g3494), .A2(g1279) );
  AND2_X1 AND2_689( .ZN(g10445), .A1(g6945), .A2(g1285) );
  AND2_X1 AND2_690( .ZN(g10446), .A1(g3522), .A2(g4930) );
  AND2_X1 AND2_691( .ZN(g10447), .A1(g7162), .A2(g4933) );
  AND2_X1 AND2_692( .ZN(g10448), .A1(g6980), .A2(g4936) );
  AND2_X1 AND2_693( .ZN(g10449), .A1(g3522), .A2(g4939) );
  AND2_X1 AND2_694( .ZN(g10450), .A1(g7162), .A2(g4942) );
  AND2_X1 AND2_695( .ZN(g10451), .A1(g3618), .A2(g4945) );
  AND2_X1 AND2_696( .ZN(g10452), .A1(g7015), .A2(g4948) );
  AND2_X1 AND2_697( .ZN(g10453), .A1(g5512), .A2(g4951) );
  AND2_X1 AND2_698( .ZN(g10454), .A1(g3618), .A2(g1825) );
  AND2_X1 AND2_699( .ZN(g10455), .A1(g3650), .A2(g1953) );
  AND2_X1 AND2_700( .ZN(g10456), .A1(g7195), .A2(g4956) );
  AND2_X1 AND2_701( .ZN(g10457), .A1(g7053), .A2(g4959) );
  AND2_X1 AND2_702( .ZN(g10458), .A1(g7195), .A2(g1970) );
  AND2_X1 AND2_703( .ZN(g10459), .A1(g7053), .A2(g1976) );
  AND2_X1 AND2_704( .ZN(g10460), .A1(g3678), .A2(g4964) );
  AND2_X1 AND2_705( .ZN(g10461), .A1(g7358), .A2(g4967) );
  AND2_X1 AND2_706( .ZN(g10462), .A1(g7230), .A2(g4970) );
  AND2_X1 AND2_707( .ZN(g10463), .A1(g3678), .A2(g4973) );
  AND2_X1 AND2_708( .ZN(g10464), .A1(g7358), .A2(g4976) );
  AND2_X1 AND2_709( .ZN(g10465), .A1(g7230), .A2(g4979) );
  AND2_X1 AND2_710( .ZN(g10466), .A1(g3722), .A2(g4982) );
  AND2_X1 AND2_711( .ZN(g10467), .A1(g3774), .A2(g4994) );
  AND2_X1 AND2_712( .ZN(g10468), .A1(g7265), .A2(g4997) );
  AND2_X1 AND2_713( .ZN(g10469), .A1(g5556), .A2(g5000) );
  AND2_X1 AND2_714( .ZN(g10470), .A1(g3774), .A2(g2510) );
  AND2_X1 AND2_715( .ZN(g10471), .A1(g7265), .A2(g2516) );
  AND2_X1 AND2_716( .ZN(g10472), .A1(g7391), .A2(g2645) );
  AND2_X1 AND2_717( .ZN(g10473), .A1(g7303), .A2(g5005) );
  AND2_X1 AND2_718( .ZN(g10474), .A1(g7303), .A2(g2661) );
  AND2_X1 AND2_719( .ZN(g10475), .A1(g3834), .A2(g5009) );
  AND2_X1 AND2_720( .ZN(g10476), .A1(g7488), .A2(g5012) );
  AND2_X1 AND2_721( .ZN(g10477), .A1(g7426), .A2(g5015) );
  AND2_X1 AND2_722( .ZN(g10478), .A1(g7488), .A2(g5018) );
  AND2_X1 AND2_723( .ZN(g10479), .A1(g7426), .A2(g5021) );
  AND3_X1 AND3_4( .ZN(II17429), .A1(g6901), .A2(g7338), .A3(g7146) );
  AND3_X1 AND3_5( .ZN(g10480), .A1(g7466), .A2(g7342), .A3(II17429) );
  AND2_X1 AND2_724( .ZN(g10485), .A1(g6448), .A2(g5024) );
  AND2_X1 AND2_725( .ZN(g10492), .A1(g3338), .A2(g5027) );
  AND2_X1 AND2_726( .ZN(g10493), .A1(g6643), .A2(g5030) );
  AND2_X1 AND2_727( .ZN(g10494), .A1(g6643), .A2(g608) );
  AND2_X1 AND2_728( .ZN(g10495), .A1(g6486), .A2(g614) );
  AND2_X1 AND2_729( .ZN(g10496), .A1(g3366), .A2(g5035) );
  AND2_X1 AND2_730( .ZN(g10497), .A1(g6912), .A2(g5038) );
  AND2_X1 AND2_731( .ZN(g10498), .A1(g3462), .A2(g5041) );
  AND2_X1 AND2_732( .ZN(g10499), .A1(g5473), .A2(g5044) );
  AND2_X1 AND2_733( .ZN(g10506), .A1(g3494), .A2(g5047) );
  AND2_X1 AND2_734( .ZN(g10507), .A1(g6945), .A2(g5050) );
  AND2_X1 AND2_735( .ZN(g10508), .A1(g6751), .A2(g5053) );
  AND2_X1 AND2_736( .ZN(g10509), .A1(g3494), .A2(g1288) );
  AND2_X1 AND2_737( .ZN(g10510), .A1(g6751), .A2(g1291) );
  AND2_X1 AND2_738( .ZN(g10511), .A1(g3522), .A2(g5058) );
  AND2_X1 AND2_739( .ZN(g10512), .A1(g7162), .A2(g5061) );
  AND2_X1 AND2_740( .ZN(g10513), .A1(g6980), .A2(g5064) );
  AND2_X1 AND2_741( .ZN(g10514), .A1(g3522), .A2(g5067) );
  AND2_X1 AND2_742( .ZN(g10515), .A1(g3618), .A2(g5072) );
  AND2_X1 AND2_743( .ZN(g10516), .A1(g7015), .A2(g5075) );
  AND2_X1 AND2_744( .ZN(g10517), .A1(g3650), .A2(g5078) );
  AND2_X1 AND2_745( .ZN(g10518), .A1(g7195), .A2(g5081) );
  AND2_X1 AND2_746( .ZN(g10519), .A1(g7053), .A2(g5084) );
  AND2_X1 AND2_747( .ZN(g10520), .A1(g3650), .A2(g1973) );
  AND2_X1 AND2_748( .ZN(g10521), .A1(g7195), .A2(g1979) );
  AND2_X1 AND2_749( .ZN(g10522), .A1(g3678), .A2(g5089) );
  AND2_X1 AND2_750( .ZN(g10523), .A1(g7358), .A2(g5092) );
  AND2_X1 AND2_751( .ZN(g10524), .A1(g7230), .A2(g5095) );
  AND2_X1 AND2_752( .ZN(g10525), .A1(g3678), .A2(g5098) );
  AND2_X1 AND2_753( .ZN(g10526), .A1(g7358), .A2(g5101) );
  AND2_X1 AND2_754( .ZN(g10527), .A1(g3774), .A2(g5104) );
  AND2_X1 AND2_755( .ZN(g10528), .A1(g7265), .A2(g5107) );
  AND2_X1 AND2_756( .ZN(g10529), .A1(g5556), .A2(g5110) );
  AND2_X1 AND2_757( .ZN(g10530), .A1(g3774), .A2(g2519) );
  AND2_X1 AND2_758( .ZN(g10531), .A1(g3806), .A2(g2647) );
  AND2_X2 AND2_759( .ZN(g10532), .A1(g7391), .A2(g5115) );
  AND2_X2 AND2_760( .ZN(g10533), .A1(g7303), .A2(g5118) );
  AND2_X1 AND2_761( .ZN(g10534), .A1(g7391), .A2(g2664) );
  AND2_X1 AND2_762( .ZN(g10535), .A1(g7303), .A2(g2670) );
  AND2_X1 AND2_763( .ZN(g10536), .A1(g3834), .A2(g5123) );
  AND2_X1 AND2_764( .ZN(g10537), .A1(g7488), .A2(g5126) );
  AND2_X1 AND2_765( .ZN(g10538), .A1(g7426), .A2(g5129) );
  AND2_X1 AND2_766( .ZN(g10539), .A1(g3834), .A2(g5132) );
  AND2_X1 AND2_767( .ZN(g10540), .A1(g7488), .A2(g5135) );
  AND2_X1 AND2_768( .ZN(g10541), .A1(g7426), .A2(g5138) );
  AND2_X1 AND2_769( .ZN(g10548), .A1(g3306), .A2(g5142) );
  AND2_X1 AND2_770( .ZN(g10555), .A1(g3338), .A2(g5145) );
  AND2_X1 AND2_771( .ZN(g10556), .A1(g3338), .A2(g611) );
  AND2_X1 AND2_772( .ZN(g10557), .A1(g6643), .A2(g617) );
  AND2_X1 AND2_773( .ZN(g10558), .A1(g3366), .A2(g5150) );
  AND2_X1 AND2_774( .ZN(g10559), .A1(g6713), .A2(g5153) );
  AND2_X1 AND2_775( .ZN(g10566), .A1(g3494), .A2(g5156) );
  AND2_X1 AND2_776( .ZN(g10567), .A1(g6945), .A2(g5159) );
  AND2_X1 AND2_777( .ZN(g10568), .A1(g6945), .A2(g1294) );
  AND2_X1 AND2_778( .ZN(g10569), .A1(g6751), .A2(g1300) );
  AND2_X1 AND2_779( .ZN(g10570), .A1(g3522), .A2(g5164) );
  AND2_X1 AND2_780( .ZN(g10571), .A1(g7162), .A2(g5167) );
  AND2_X1 AND2_781( .ZN(g10572), .A1(g3618), .A2(g5170) );
  AND2_X1 AND2_782( .ZN(g10573), .A1(g5512), .A2(g5173) );
  AND2_X1 AND2_783( .ZN(g10580), .A1(g3650), .A2(g5176) );
  AND2_X1 AND2_784( .ZN(g10581), .A1(g7195), .A2(g5179) );
  AND2_X1 AND2_785( .ZN(g10582), .A1(g7053), .A2(g5182) );
  AND2_X1 AND2_786( .ZN(g10583), .A1(g3650), .A2(g1982) );
  AND2_X1 AND2_787( .ZN(g10584), .A1(g7053), .A2(g1985) );
  AND2_X1 AND2_788( .ZN(g10585), .A1(g3678), .A2(g5187) );
  AND2_X1 AND2_789( .ZN(g10586), .A1(g7358), .A2(g5190) );
  AND2_X1 AND2_790( .ZN(g10587), .A1(g7230), .A2(g5193) );
  AND2_X1 AND2_791( .ZN(g10588), .A1(g3678), .A2(g5196) );
  AND2_X1 AND2_792( .ZN(g10589), .A1(g3774), .A2(g5201) );
  AND2_X1 AND2_793( .ZN(g10590), .A1(g7265), .A2(g5204) );
  AND2_X1 AND2_794( .ZN(g10591), .A1(g3806), .A2(g5207) );
  AND2_X1 AND2_795( .ZN(g10592), .A1(g7391), .A2(g5210) );
  AND2_X1 AND2_796( .ZN(g10593), .A1(g7303), .A2(g5213) );
  AND2_X1 AND2_797( .ZN(g10594), .A1(g3806), .A2(g2667) );
  AND2_X1 AND2_798( .ZN(g10595), .A1(g7391), .A2(g2673) );
  AND2_X1 AND2_799( .ZN(g10596), .A1(g3834), .A2(g5218) );
  AND2_X1 AND2_800( .ZN(g10597), .A1(g7488), .A2(g5221) );
  AND2_X1 AND2_801( .ZN(g10598), .A1(g7426), .A2(g5224) );
  AND2_X1 AND2_802( .ZN(g10599), .A1(g3834), .A2(g5227) );
  AND2_X1 AND2_803( .ZN(g10600), .A1(g7488), .A2(g5230) );
  AND2_X1 AND2_804( .ZN(g10604), .A1(g3338), .A2(g620) );
  AND2_X1 AND2_805( .ZN(g10605), .A1(g3462), .A2(g5235) );
  AND2_X1 AND2_806( .ZN(g10612), .A1(g3494), .A2(g5238) );
  AND2_X1 AND2_807( .ZN(g10613), .A1(g3494), .A2(g1297) );
  AND2_X1 AND2_808( .ZN(g10614), .A1(g6945), .A2(g1303) );
  AND2_X1 AND2_809( .ZN(g10615), .A1(g3522), .A2(g5243) );
  AND2_X1 AND2_810( .ZN(g10616), .A1(g7015), .A2(g5246) );
  AND2_X1 AND2_811( .ZN(g10623), .A1(g3650), .A2(g5249) );
  AND2_X1 AND2_812( .ZN(g10624), .A1(g7195), .A2(g5252) );
  AND2_X1 AND2_813( .ZN(g10625), .A1(g7195), .A2(g1988) );
  AND2_X1 AND2_814( .ZN(g10626), .A1(g7053), .A2(g1994) );
  AND2_X1 AND2_815( .ZN(g10627), .A1(g3678), .A2(g5257) );
  AND2_X1 AND2_816( .ZN(g10628), .A1(g7358), .A2(g5260) );
  AND2_X1 AND2_817( .ZN(g10629), .A1(g3774), .A2(g5263) );
  AND2_X1 AND2_818( .ZN(g10630), .A1(g5556), .A2(g5266) );
  AND2_X1 AND2_819( .ZN(g10637), .A1(g3806), .A2(g5269) );
  AND2_X1 AND2_820( .ZN(g10638), .A1(g7391), .A2(g5272) );
  AND2_X1 AND2_821( .ZN(g10639), .A1(g7303), .A2(g5275) );
  AND2_X1 AND2_822( .ZN(g10640), .A1(g3806), .A2(g2676) );
  AND2_X1 AND2_823( .ZN(g10641), .A1(g7303), .A2(g2679) );
  AND2_X1 AND2_824( .ZN(g10642), .A1(g3834), .A2(g5280) );
  AND2_X1 AND2_825( .ZN(g10643), .A1(g7488), .A2(g5283) );
  AND2_X1 AND2_826( .ZN(g10644), .A1(g7426), .A2(g5286) );
  AND2_X1 AND2_827( .ZN(g10645), .A1(g3834), .A2(g5289) );
  AND2_X1 AND2_828( .ZN(g10650), .A1(g6678), .A2(g5293) );
  AND2_X1 AND2_829( .ZN(g10651), .A1(g3494), .A2(g1306) );
  AND2_X1 AND2_830( .ZN(g10652), .A1(g3618), .A2(g5298) );
  AND2_X1 AND2_831( .ZN(g10659), .A1(g3650), .A2(g5301) );
  AND2_X1 AND2_832( .ZN(g10660), .A1(g3650), .A2(g1991) );
  AND2_X1 AND2_833( .ZN(g10661), .A1(g7195), .A2(g1997) );
  AND2_X1 AND2_834( .ZN(g10662), .A1(g3678), .A2(g5306) );
  AND2_X1 AND2_835( .ZN(g10663), .A1(g7265), .A2(g5309) );
  AND2_X1 AND2_836( .ZN(g10670), .A1(g3806), .A2(g5312) );
  AND2_X1 AND2_837( .ZN(g10671), .A1(g7391), .A2(g5315) );
  AND2_X1 AND2_838( .ZN(g10672), .A1(g7391), .A2(g2682) );
  AND2_X1 AND2_839( .ZN(g10673), .A1(g7303), .A2(g2688) );
  AND2_X1 AND2_840( .ZN(g10674), .A1(g3834), .A2(g5320) );
  AND2_X1 AND2_841( .ZN(g10675), .A1(g7488), .A2(g5323) );
  AND2_X1 AND2_842( .ZN(g10678), .A1(g6912), .A2(g5327) );
  AND2_X1 AND2_843( .ZN(g10680), .A1(g6980), .A2(g5330) );
  AND2_X1 AND2_844( .ZN(g10681), .A1(g3650), .A2(g2000) );
  AND2_X1 AND2_845( .ZN(g10682), .A1(g3774), .A2(g5335) );
  AND2_X1 AND2_846( .ZN(g10689), .A1(g3806), .A2(g5338) );
  AND2_X1 AND2_847( .ZN(g10690), .A1(g3806), .A2(g2685) );
  AND2_X1 AND2_848( .ZN(g10691), .A1(g7391), .A2(g2691) );
  AND2_X1 AND2_849( .ZN(g10692), .A1(g3834), .A2(g5343) );
  AND4_X1 AND4_10( .ZN(g10693), .A1(g7462), .A2(g7522), .A3(g2924), .A4(g7545) );
  AND2_X1 AND2_850( .ZN(g10704), .A1(g3366), .A2(g5352) );
  AND2_X1 AND2_851( .ZN(g10707), .A1(g7162), .A2(g5355) );
  AND2_X1 AND2_852( .ZN(g10709), .A1(g7230), .A2(g5358) );
  AND2_X1 AND2_853( .ZN(g10710), .A1(g3806), .A2(g2694) );
  AND3_X1 AND3_6( .ZN(II17599), .A1(g7566), .A2(g7583), .A3(g7587) );
  AND3_X4 AND3_7( .ZN(g10711), .A1(g7595), .A2(g7600), .A3(II17599) );
  AND2_X1 AND2_854( .ZN(g10724), .A1(g3522), .A2(g5369) );
  AND2_X1 AND2_855( .ZN(g10727), .A1(g7358), .A2(g5372) );
  AND2_X1 AND2_856( .ZN(g10729), .A1(g7426), .A2(g5375) );
  AND2_X1 AND2_857( .ZN(g10745), .A1(g3678), .A2(g5382) );
  AND2_X1 AND2_858( .ZN(g10748), .A1(g7488), .A2(g5385) );
  AND2_X1 AND2_859( .ZN(g10764), .A1(g3834), .A2(g5391) );
  AND2_X1 AND2_860( .ZN(g11347), .A1(g6232), .A2(g213) );
  AND2_X1 AND2_861( .ZN(g11420), .A1(g6314), .A2(g216) );
  AND2_X1 AND2_862( .ZN(g11421), .A1(g6232), .A2(g222) );
  AND2_X1 AND2_863( .ZN(g11431), .A1(g6369), .A2(g900) );
  AND2_X1 AND2_864( .ZN(g11607), .A1(g5871), .A2(g8360) );
  AND2_X1 AND2_865( .ZN(g11612), .A1(g5881), .A2(g8378) );
  AND2_X1 AND2_866( .ZN(g11637), .A1(g5918), .A2(g8427) );
  AND2_X1 AND2_867( .ZN(g11771), .A1(g554), .A2(g8622) );
  AND2_X1 AND2_868( .ZN(g11788), .A1(g1240), .A2(g8632) );
  AND2_X1 AND2_869( .ZN(g11805), .A1(g6173), .A2(g8643) );
  AND2_X1 AND2_870( .ZN(g11814), .A1(g1934), .A2(g8651) );
  AND2_X1 AND2_871( .ZN(g11816), .A1(g7869), .A2(g8655) );
  AND2_X1 AND2_872( .ZN(g11838), .A1(g6205), .A2(g8659) );
  AND2_X1 AND2_873( .ZN(g11847), .A1(g2628), .A2(g8667) );
  AND2_X1 AND2_874( .ZN(g11851), .A1(g7849), .A2(g8670) );
  AND2_X2 AND2_875( .ZN(g11880), .A1(g6294), .A2(g8678) );
  AND2_X2 AND2_876( .ZN(g11885), .A1(g7834), .A2(g8684) );
  AND2_X1 AND2_877( .ZN(g11922), .A1(g6431), .A2(g8690) );
  AND2_X1 AND2_878( .ZN(g11926), .A1(g8169), .A2(g8696) );
  AND2_X1 AND2_879( .ZN(g11966), .A1(g8090), .A2(g8708) );
  AND2_X1 AND2_880( .ZN(g11967), .A1(g7967), .A2(g8711) );
  AND2_X1 AND2_881( .ZN(g12012), .A1(g8015), .A2(g8745) );
  AND2_X1 AND2_882( .ZN(g12069), .A1(g7964), .A2(g8763) );
  AND2_X1 AND2_883( .ZN(g12070), .A1(g8018), .A2(g8766) );
  AND2_X1 AND2_884( .ZN(g12128), .A1(g7916), .A2(g8785) );
  AND2_X1 AND2_885( .ZN(g12129), .A1(g7872), .A2(g8788) );
  AND2_X1 AND2_886( .ZN(g12186), .A1(g8093), .A2(g8805) );
  AND2_X1 AND2_887( .ZN(g12273), .A1(g8172), .A2(g8829) );
  AND2_X1 AND2_888( .ZN(g12274), .A1(g7900), .A2(g8832) );
  AND2_X1 AND2_889( .ZN(g12307), .A1(g7919), .A2(g8853) );
  AND2_X1 AND2_890( .ZN(g12330), .A1(g8246), .A2(g8879) );
  AND2_X1 AND2_891( .ZN(g12331), .A1(g7927), .A2(g8882) );
  AND2_X1 AND2_892( .ZN(g12353), .A1(g7852), .A2(g8915) );
  AND2_X1 AND2_893( .ZN(g12376), .A1(g7974), .A2(g8949) );
  AND2_X1 AND2_894( .ZN(g12419), .A1(g8028), .A2(g9006) );
  AND2_X1 AND2_895( .ZN(g12429), .A1(g8101), .A2(g9044) );
  AND2_X1 AND2_896( .ZN(g12477), .A1(g7822), .A2(g9128) );
  AND2_X1 AND2_897( .ZN(g12494), .A1(g7833), .A2(g9134) );
  AND2_X1 AND2_898( .ZN(g12514), .A1(g7848), .A2(g9140) );
  AND2_X1 AND2_899( .ZN(g12531), .A1(g7868), .A2(g9146) );
  AND2_X1 AND2_900( .ZN(g12650), .A1(g6149), .A2(g9290) );
  AND4_X1 AND4_11( .ZN(II19937), .A1(g9507), .A2(g9427), .A3(g9356), .A4(g9293) );
  AND4_X1 AND4_12( .ZN(II19938), .A1(g9232), .A2(g9187), .A3(g9161), .A4(g9150) );
  AND2_X1 AND2_901( .ZN(g12876), .A1(II19937), .A2(II19938) );
  AND2_X1 AND2_902( .ZN(g12908), .A1(g7899), .A2(g10004) );
  AND4_X1 AND4_13( .ZN(II19971), .A1(g9649), .A2(g9569), .A3(g9453), .A4(g9374) );
  AND4_X1 AND4_14( .ZN(II19972), .A1(g9310), .A2(g9248), .A3(g9203), .A4(g9174) );
  AND2_X1 AND2_903( .ZN(g12916), .A1(II19971), .A2(II19972) );
  AND2_X1 AND2_904( .ZN(g12938), .A1(g8179), .A2(g10096) );
  AND4_X1 AND4_15( .ZN(II19996), .A1(g9795), .A2(g9711), .A3(g9595), .A4(g9471) );
  AND4_X1 AND4_16( .ZN(II19997), .A1(g9391), .A2(g9326), .A3(g9264), .A4(g9216) );
  AND2_X1 AND2_905( .ZN(g12945), .A1(II19996), .A2(II19997) );
  AND2_X1 AND2_906( .ZN(g12966), .A1(g7926), .A2(g10189) );
  AND4_X1 AND4_17( .ZN(II20021), .A1(g9941), .A2(g9857), .A3(g9737), .A4(g9613) );
  AND4_X1 AND4_18( .ZN(II20022), .A1(g9488), .A2(g9407), .A3(g9342), .A4(g9277) );
  AND2_X1 AND2_907( .ZN(g12974), .A1(II20021), .A2(II20022) );
  AND2_X1 AND2_908( .ZN(g12989), .A1(g8254), .A2(g10273) );
  AND2_X1 AND2_909( .ZN(g12990), .A1(g8180), .A2(g10276) );
  AND2_X1 AND2_910( .ZN(g13000), .A1(g7973), .A2(g10357) );
  AND2_X1 AND2_911( .ZN(g13004), .A1(g10186), .A2(g8317) );
  AND2_X1 AND2_912( .ZN(g13009), .A1(g3995), .A2(g10416) );
  AND2_X1 AND2_913( .ZN(g13010), .A1(g8255), .A2(g10419) );
  AND2_X1 AND2_914( .ZN(g13023), .A1(g8027), .A2(g10482) );
  AND2_X1 AND2_915( .ZN(g13031), .A1(g7879), .A2(g10542) );
  AND2_X1 AND2_916( .ZN(g13032), .A1(g3996), .A2(g10545) );
  AND2_X1 AND2_917( .ZN(g13042), .A1(g8100), .A2(g10601) );
  AND3_X1 AND3_8( .ZN(II20100), .A1(g10186), .A2(g3018), .A3(g3028) );
  AND3_X1 AND3_9( .ZN(g13055), .A1(g7471), .A2(g7570), .A3(II20100) );
  AND2_X1 AND2_918( .ZN(g13056), .A1(g4092), .A2(g10646) );
  AND4_X1 AND4_19( .ZN(II20131), .A1(g8313), .A2(g7542), .A3(g2888), .A4(g7566) );
  AND4_X1 AND4_20( .ZN(II20132), .A1(g2892), .A2(g2903), .A3(g7595), .A4(g2908) );
  AND2_X1 AND2_919( .ZN(g13082), .A1(II20131), .A2(II20132) );
  AND4_X1 AND4_21( .ZN(g13110), .A1(g10693), .A2(g2883), .A3(g7562), .A4(g10711) );
  AND2_X2 AND2_920( .ZN(g13247), .A1(g298), .A2(g11032) );
  AND2_X2 AND2_921( .ZN(g13266), .A1(g5628), .A2(g11088) );
  AND2_X1 AND2_922( .ZN(g13270), .A1(g985), .A2(g11102) );
  AND2_X1 AND2_923( .ZN(g13289), .A1(g5647), .A2(g11141) );
  AND2_X1 AND2_924( .ZN(g13291), .A1(g5656), .A2(g11154) );
  AND2_X1 AND2_925( .ZN(g13295), .A1(g1679), .A2(g11170) );
  AND2_X1 AND2_926( .ZN(g13316), .A1(g5675), .A2(g11210) );
  AND2_X1 AND2_927( .ZN(g13320), .A1(g5685), .A2(g11225) );
  AND2_X1 AND2_928( .ZN(g13322), .A1(g5694), .A2(g11240) );
  AND2_X1 AND2_929( .ZN(g13326), .A1(g2373), .A2(g11256) );
  AND2_X1 AND2_930( .ZN(g13335), .A1(g5708), .A2(g11278) );
  AND2_X1 AND2_931( .ZN(g13340), .A1(g5727), .A2(g11294) );
  AND2_X1 AND2_932( .ZN(g13343), .A1(g5737), .A2(g11309) );
  AND2_X1 AND2_933( .ZN(g13345), .A1(g5746), .A2(g11324) );
  AND2_X1 AND2_934( .ZN(g13355), .A1(g5756), .A2(g11355) );
  AND2_X1 AND2_935( .ZN(g13360), .A1(g5766), .A2(g11373) );
  AND2_X1 AND2_936( .ZN(g13365), .A1(g5785), .A2(g11389) );
  AND2_X1 AND2_937( .ZN(g13368), .A1(g5795), .A2(g11404) );
  AND2_X1 AND2_938( .ZN(g13385), .A1(g5815), .A2(g11441) );
  AND2_X1 AND2_939( .ZN(g13390), .A1(g5825), .A2(g11459) );
  AND2_X1 AND2_940( .ZN(g13395), .A1(g5844), .A2(g11475) );
  AND2_X1 AND2_941( .ZN(g13477), .A1(g6016), .A2(g12191) );
  AND2_X1 AND2_942( .ZN(g13479), .A1(g6017), .A2(g12196) );
  AND2_X1 AND2_943( .ZN(g13480), .A1(g6018), .A2(g12197) );
  AND2_X1 AND2_944( .ZN(g13481), .A1(g5864), .A2(g11603) );
  AND2_X1 AND2_945( .ZN(g13483), .A1(g6020), .A2(g12209) );
  AND2_X1 AND2_946( .ZN(g13484), .A1(g6021), .A2(g12210) );
  AND2_X1 AND2_947( .ZN(g13485), .A1(g6022), .A2(g12211) );
  AND2_X1 AND2_948( .ZN(g13486), .A1(g6023), .A2(g12212) );
  AND2_X1 AND2_949( .ZN(g13487), .A1(g5874), .A2(g11608) );
  AND2_X1 AND2_950( .ZN(g13488), .A1(g6025), .A2(g12218) );
  AND2_X1 AND2_951( .ZN(g13489), .A1(g6026), .A2(g12219) );
  AND2_X1 AND2_952( .ZN(g13490), .A1(g6027), .A2(g12220) );
  AND2_X1 AND2_953( .ZN(g13491), .A1(g6028), .A2(g12221) );
  AND2_X1 AND2_954( .ZN(g13492), .A1(g2371), .A2(g12222) );
  AND2_X1 AND2_955( .ZN(g13493), .A1(g5887), .A2(g11613) );
  AND2_X1 AND2_956( .ZN(g13496), .A1(g6032), .A2(g12246) );
  AND2_X1 AND2_957( .ZN(g13498), .A1(g6033), .A2(g12251) );
  AND2_X1 AND2_958( .ZN(g13499), .A1(g6034), .A2(g12252) );
  AND2_X1 AND2_959( .ZN(g13500), .A1(g5911), .A2(g11633) );
  AND2_X1 AND2_960( .ZN(g13502), .A1(g6036), .A2(g12264) );
  AND2_X1 AND2_961( .ZN(g13503), .A1(g6037), .A2(g12265) );
  AND2_X1 AND2_962( .ZN(g13504), .A1(g6038), .A2(g12266) );
  AND2_X1 AND2_963( .ZN(g13505), .A1(g6039), .A2(g12267) );
  AND2_X1 AND2_964( .ZN(g13506), .A1(g5921), .A2(g11638) );
  AND2_X1 AND2_965( .ZN(g13513), .A1(g6043), .A2(g12289) );
  AND2_X1 AND2_966( .ZN(g13515), .A1(g6044), .A2(g12294) );
  AND2_X1 AND2_967( .ZN(g13516), .A1(g6045), .A2(g12295) );
  AND2_X1 AND2_968( .ZN(g13517), .A1(g5950), .A2(g11656) );
  AND2_X1 AND2_969( .ZN(g13527), .A1(g6047), .A2(g12325) );
  AND2_X1 AND2_970( .ZN(g13609), .A1(g6141), .A2(g12456) );
  AND2_X1 AND2_971( .ZN(g13619), .A1(g6162), .A2(g12466) );
  AND2_X1 AND2_972( .ZN(g13623), .A1(g5428), .A2(g12472) );
  AND2_X1 AND2_973( .ZN(g13625), .A1(g6173), .A2(g12476) );
  AND2_X1 AND2_974( .ZN(g13631), .A1(g6189), .A2(g12481) );
  AND2_X1 AND2_975( .ZN(g13634), .A1(g12776), .A2(g8617) );
  AND2_X1 AND2_976( .ZN(g13636), .A1(g6205), .A2(g12493) );
  AND2_X1 AND2_977( .ZN(g13642), .A1(g6221), .A2(g12498) );
  AND2_X1 AND2_978( .ZN(g13643), .A1(g5431), .A2(g12502) );
  AND2_X1 AND2_979( .ZN(g13645), .A1(g6281), .A2(g12504) );
  AND2_X2 AND2_980( .ZN(g13646), .A1(g7772), .A2(g12505) );
  AND2_X2 AND2_981( .ZN(g13648), .A1(g6294), .A2(g12513) );
  AND2_X2 AND2_982( .ZN(g13654), .A1(g8093), .A2(g11791) );
  AND2_X1 AND2_983( .ZN(g13655), .A1(g7540), .A2(g12518) );
  AND2_X1 AND2_984( .ZN(g13656), .A1(g12776), .A2(g8640) );
  AND2_X1 AND2_985( .ZN(g13671), .A1(g6418), .A2(g12521) );
  AND2_X1 AND2_986( .ZN(g13672), .A1(g7788), .A2(g12522) );
  AND2_X1 AND2_987( .ZN(g13674), .A1(g6431), .A2(g12530) );
  AND2_X1 AND2_988( .ZN(g13675), .A1(g7561), .A2(g12532) );
  AND2_X1 AND2_989( .ZN(g13676), .A1(g5434), .A2(g12533) );
  AND2_X1 AND2_990( .ZN(g13701), .A1(g6623), .A2(g12536) );
  AND2_X1 AND2_991( .ZN(g13702), .A1(g7802), .A2(g12537) );
  AND2_X1 AND2_992( .ZN(g13703), .A1(g8018), .A2(g11848) );
  AND2_X1 AND2_993( .ZN(g13704), .A1(g7581), .A2(g12542) );
  AND2_X1 AND2_994( .ZN(g13705), .A1(g12776), .A2(g8673) );
  AND2_X1 AND2_995( .ZN(g13738), .A1(g6887), .A2(g12545) );
  AND2_X1 AND2_996( .ZN(g13739), .A1(g7815), .A2(g12546) );
  AND2_X1 AND2_997( .ZN(g13740), .A1(g6636), .A2(g12547) );
  AND2_X1 AND2_998( .ZN(g13755), .A1(g7347), .A2(g12551) );
  AND2_X1 AND2_999( .ZN(g13787), .A1(g7967), .A2(g11923) );
  AND2_X1 AND2_1000( .ZN(g13788), .A1(g6897), .A2(g12553) );
  AND2_X1 AND2_1001( .ZN(g13789), .A1(g7140), .A2(g12554) );
  AND2_X1 AND2_1002( .ZN(g13790), .A1(g7475), .A2(g12558) );
  AND2_X1 AND2_1003( .ZN(g13796), .A1(g7477), .A2(g12559) );
  AND2_X1 AND2_1004( .ZN(g13815), .A1(g7139), .A2(g12560) );
  AND2_X1 AND2_1005( .ZN(g13816), .A1(g7530), .A2(g12596) );
  AND2_X1 AND2_1006( .ZN(g13818), .A1(g7531), .A2(g12597) );
  AND2_X1 AND2_1007( .ZN(g13824), .A1(g7533), .A2(g12598) );
  AND2_X1 AND2_1008( .ZN(g13833), .A1(g7919), .A2(g12009) );
  AND2_X1 AND2_1009( .ZN(g13834), .A1(g7336), .A2(g12599) );
  AND2_X1 AND2_1010( .ZN(g13835), .A1(g7461), .A2(g12600) );
  AND2_X1 AND2_1011( .ZN(g13837), .A1(g7556), .A2(g12642) );
  AND2_X1 AND2_1012( .ZN(g13839), .A1(g7557), .A2(g12643) );
  AND2_X1 AND2_1013( .ZN(g13845), .A1(g7559), .A2(g12644) );
  AND2_X1 AND2_1014( .ZN(g13846), .A1(g7460), .A2(g12645) );
  AND2_X1 AND2_1015( .ZN(g13847), .A1(g7521), .A2(g12646) );
  AND2_X1 AND2_1016( .ZN(g13851), .A1(g7579), .A2(g12688) );
  AND2_X1 AND2_1017( .ZN(g13853), .A1(g7580), .A2(g12689) );
  AND2_X1 AND2_1018( .ZN(g13854), .A1(g5349), .A2(g12690) );
  AND2_X1 AND2_1019( .ZN(g13855), .A1(g7541), .A2(g12691) );
  AND2_X1 AND2_1020( .ZN(g13860), .A1(g7593), .A2(g12742) );
  AND2_X1 AND2_1021( .ZN(g13862), .A1(g5366), .A2(g12743) );
  AND2_X1 AND2_1022( .ZN(g13865), .A1(g548), .A2(g12748) );
  AND2_X1 AND2_1023( .ZN(g13870), .A1(g7582), .A2(g12768) );
  AND2_X1 AND2_1024( .ZN(g13871), .A1(g7898), .A2(g12775) );
  AND2_X1 AND2_1025( .ZN(g13878), .A1(g7610), .A2(g12782) );
  AND2_X1 AND2_1026( .ZN(g13880), .A1(g1234), .A2(g12790) );
  AND2_X1 AND2_1027( .ZN(g13884), .A1(g7594), .A2(g12807) );
  AND2_X1 AND2_1028( .ZN(g13892), .A1(g7616), .A2(g12815) );
  AND2_X1 AND2_1029( .ZN(g13900), .A1(g7619), .A2(g12821) );
  AND2_X1 AND2_1030( .ZN(g13902), .A1(g1928), .A2(g12829) );
  AND2_X1 AND2_1031( .ZN(g13904), .A1(g7337), .A2(g12843) );
  AND2_X1 AND2_1032( .ZN(g13905), .A1(g7925), .A2(g12847) );
  AND2_X1 AND2_1033( .ZN(g13913), .A1(g7623), .A2(g12850) );
  AND2_X1 AND2_1034( .ZN(g13914), .A1(g7626), .A2(g12851) );
  AND2_X1 AND2_1035( .ZN(g13933), .A1(g7632), .A2(g12853) );
  AND2_X1 AND2_1036( .ZN(g13941), .A1(g7635), .A2(g12859) );
  AND2_X1 AND2_1037( .ZN(g13943), .A1(g2622), .A2(g12867) );
  AND2_X1 AND2_1038( .ZN(g13944), .A1(g7141), .A2(g12874) );
  AND2_X1 AND2_1039( .ZN(g13952), .A1(g7643), .A2(g12881) );
  AND2_X1 AND2_1040( .ZN(g13953), .A1(g7646), .A2(g12882) );
  AND2_X1 AND2_1041( .ZN(g13969), .A1(g7652), .A2(g12891) );
  AND2_X1 AND2_1042( .ZN(g13970), .A1(g7655), .A2(g12892) );
  AND2_X1 AND2_1043( .ZN(g13989), .A1(g7661), .A2(g12894) );
  AND2_X1 AND2_1044( .ZN(g13997), .A1(g7664), .A2(g12900) );
  AND2_X1 AND2_1045( .ZN(g13998), .A1(g7972), .A2(g12907) );
  AND2_X1 AND2_1046( .ZN(g14006), .A1(g7670), .A2(g12914) );
  AND2_X1 AND2_1047( .ZN(g14007), .A1(g7673), .A2(g12915) );
  AND2_X1 AND2_1048( .ZN(g14022), .A1(g7679), .A2(g12921) );
  AND2_X1 AND2_1049( .ZN(g14023), .A1(g7682), .A2(g12922) );
  AND2_X1 AND2_1050( .ZN(g14039), .A1(g7688), .A2(g12931) );
  AND2_X1 AND2_1051( .ZN(g14040), .A1(g7691), .A2(g12932) );
  AND2_X1 AND2_1052( .ZN(g14059), .A1(g7697), .A2(g12934) );
  AND2_X1 AND2_1053( .ZN(g14067), .A1(g7703), .A2(g12940) );
  AND2_X1 AND2_1054( .ZN(g14097), .A1(g7706), .A2(g12943) );
  AND2_X1 AND2_1055( .ZN(g14098), .A1(g7709), .A2(g12944) );
  AND2_X1 AND2_1056( .ZN(g14113), .A1(g7715), .A2(g12950) );
  AND2_X1 AND2_1057( .ZN(g14114), .A1(g7718), .A2(g12951) );
  AND2_X1 AND2_1058( .ZN(g14130), .A1(g7724), .A2(g12960) );
  AND2_X1 AND2_1059( .ZN(g14131), .A1(g7727), .A2(g12961) );
  AND2_X1 AND2_1060( .ZN(g14143), .A1(g8026), .A2(g12965) );
  AND2_X1 AND2_1061( .ZN(g14182), .A1(g7733), .A2(g12969) );
  AND2_X1 AND2_1062( .ZN(g14212), .A1(g7736), .A2(g12972) );
  AND2_X1 AND2_1063( .ZN(g14213), .A1(g7739), .A2(g12973) );
  AND2_X1 AND2_1064( .ZN(g14228), .A1(g7745), .A2(g12979) );
  AND2_X1 AND2_1065( .ZN(g14229), .A1(g7748), .A2(g12980) );
  AND2_X1 AND2_1066( .ZN(g14297), .A1(g7757), .A2(g12993) );
  AND2_X1 AND2_1067( .ZN(g14327), .A1(g7760), .A2(g12996) );
  AND2_X1 AND2_1068( .ZN(g14328), .A1(g7763), .A2(g12997) );
  AND2_X1 AND2_1069( .ZN(g14336), .A1(g8099), .A2(g12998) );
  AND2_X1 AND2_1070( .ZN(g14419), .A1(g7779), .A2(g13003) );
  AND2_X1 AND2_1071( .ZN(g14690), .A1(g7841), .A2(g13101) );
  AND2_X1 AND2_1072( .ZN(g14724), .A1(g7861), .A2(g13117) );
  AND2_X1 AND2_1073( .ZN(g14752), .A1(g7891), .A2(g13130) );
  AND2_X1 AND2_1074( .ZN(g14767), .A1(g13245), .A2(g10765) );
  AND2_X1 AND2_1075( .ZN(g14773), .A1(g7915), .A2(g13141) );
  AND2_X1 AND2_1076( .ZN(g14884), .A1(g8169), .A2(g12548) );
  AND2_X1 AND2_1077( .ZN(g14894), .A1(g3940), .A2(g13148) );
  AND2_X1 AND2_1078( .ZN(g14956), .A1(g11059), .A2(g13151) );
  AND2_X1 AND2_1079( .ZN(g14957), .A1(g4015), .A2(g13152) );
  AND2_X1 AND2_1080( .ZN(g14958), .A1(g4016), .A2(g13153) );
  AND2_X1 AND2_1081( .ZN(g14975), .A1(g4047), .A2(g13154) );
  AND2_X1 AND2_1082( .ZN(g15020), .A1(g8090), .A2(g12561) );
  AND2_X1 AND2_1083( .ZN(g15030), .A1(g4110), .A2(g13158) );
  AND2_X1 AND2_1084( .ZN(g15031), .A1(g4111), .A2(g13159) );
  AND2_X1 AND2_1085( .ZN(g15046), .A1(g4142), .A2(g13161) );
  AND2_X1 AND2_1086( .ZN(g15047), .A1(g4143), .A2(g13162) );
  AND2_X1 AND2_1087( .ZN(g15064), .A1(g4174), .A2(g13163) );
  AND2_X1 AND2_1088( .ZN(g15093), .A1(g7869), .A2(g12601) );
  AND2_X1 AND2_1089( .ZN(g15094), .A1(g7872), .A2(g12604) );
  AND2_X1 AND2_1090( .ZN(g15104), .A1(g4220), .A2(g13167) );
  AND2_X1 AND2_1091( .ZN(g15105), .A1(g4224), .A2(g13168) );
  AND2_X1 AND2_1092( .ZN(g15126), .A1(g4249), .A2(g13169) );
  AND2_X1 AND2_1093( .ZN(g15127), .A1(g4250), .A2(g13170) );
  AND2_X1 AND2_1094( .ZN(g15142), .A1(g4281), .A2(g13172) );
  AND2_X1 AND2_1095( .ZN(g15143), .A1(g4282), .A2(g13173) );
  AND2_X1 AND2_1096( .ZN(g15160), .A1(g4313), .A2(g13174) );
  AND2_X1 AND2_1097( .ZN(g15171), .A1(g8015), .A2(g12647) );
  AND2_X1 AND2_1098( .ZN(g15172), .A1(g4346), .A2(g13176) );
  AND2_X1 AND2_1099( .ZN(g15173), .A1(g4347), .A2(g13177) );
  AND2_X1 AND2_1100( .ZN(g15178), .A1(g640), .A2(g12651) );
  AND2_X1 AND2_1101( .ZN(g15196), .A1(g4375), .A2(g13178) );
  AND2_X1 AND2_1102( .ZN(g15197), .A1(g4379), .A2(g13179) );
  AND2_X1 AND2_1103( .ZN(g15218), .A1(g4404), .A2(g13180) );
  AND2_X1 AND2_1104( .ZN(g15219), .A1(g4405), .A2(g13181) );
  AND2_X1 AND2_1105( .ZN(g15234), .A1(g4436), .A2(g13183) );
  AND2_X1 AND2_1106( .ZN(g15235), .A1(g4437), .A2(g13184) );
  AND2_X1 AND2_1107( .ZN(g15243), .A1(g7849), .A2(g12692) );
  AND2_X1 AND2_1108( .ZN(g15244), .A1(g7852), .A2(g12695) );
  AND2_X1 AND2_1109( .ZN(g15245), .A1(g4474), .A2(g13185) );
  AND2_X1 AND2_1110( .ZN(g15246), .A1(g4475), .A2(g13186) );
  AND2_X1 AND2_1111( .ZN(g15247), .A1(g4479), .A2(g13187) );
  AND2_X1 AND2_1112( .ZN(g15257), .A1(g4357), .A2(g12702) );
  AND2_X1 AND2_1113( .ZN(g15258), .A1(g4515), .A2(g13188) );
  AND2_X1 AND2_1114( .ZN(g15259), .A1(g4516), .A2(g13189) );
  AND2_X1 AND2_1115( .ZN(g15264), .A1(g1326), .A2(g12705) );
  AND2_X1 AND2_1116( .ZN(g15282), .A1(g4544), .A2(g13190) );
  AND2_X1 AND2_1117( .ZN(g15283), .A1(g4548), .A2(g13191) );
  AND2_X1 AND2_1118( .ZN(g15304), .A1(g4573), .A2(g13192) );
  AND2_X1 AND2_1119( .ZN(g15305), .A1(g4574), .A2(g13193) );
  AND2_X1 AND2_1120( .ZN(g15320), .A1(g7964), .A2(g12744) );
  AND2_X1 AND2_1121( .ZN(g15321), .A1(g4601), .A2(g13195) );
  AND2_X1 AND2_1122( .ZN(g15324), .A1(g4609), .A2(g13196) );
  AND2_X1 AND2_1123( .ZN(g15325), .A1(g4610), .A2(g13197) );
  AND2_X1 AND2_1124( .ZN(g15335), .A1(g4489), .A2(g12749) );
  AND2_X1 AND2_1125( .ZN(g15336), .A1(g4492), .A2(g12752) );
  AND2_X1 AND2_1126( .ZN(g15337), .A1(g4650), .A2(g13198) );
  AND2_X1 AND2_1127( .ZN(g15338), .A1(g4651), .A2(g13199) );
  AND2_X1 AND2_1128( .ZN(g15339), .A1(g4655), .A2(g13200) );
  AND2_X1 AND2_1129( .ZN(g15349), .A1(g4526), .A2(g12759) );
  AND2_X1 AND2_1130( .ZN(g15350), .A1(g4691), .A2(g13201) );
  AND2_X1 AND2_1131( .ZN(g15351), .A1(g4692), .A2(g13202) );
  AND2_X1 AND2_1132( .ZN(g15356), .A1(g2020), .A2(g12762) );
  AND2_X1 AND2_1133( .ZN(g15374), .A1(g4720), .A2(g13203) );
  AND2_X1 AND2_1134( .ZN(g15375), .A1(g4724), .A2(g13204) );
  AND2_X1 AND2_1135( .ZN(g15388), .A1(g7834), .A2(g12769) );
  AND2_X1 AND2_1136( .ZN(g15389), .A1(g8246), .A2(g12772) );
  AND2_X1 AND2_1137( .ZN(g15391), .A1(g4752), .A2(g13205) );
  AND2_X1 AND2_1138( .ZN(g15392), .A1(g4753), .A2(g13206) );
  AND2_X1 AND2_1139( .ZN(g15402), .A1(g4620), .A2(g12783) );
  AND2_X1 AND2_1140( .ZN(g15403), .A1(g4623), .A2(g12786) );
  AND2_X1 AND2_1141( .ZN(g15407), .A1(g4778), .A2(g13207) );
  AND2_X1 AND2_1142( .ZN(g15410), .A1(g4786), .A2(g13208) );
  AND2_X1 AND2_1143( .ZN(g15411), .A1(g4787), .A2(g13209) );
  AND2_X1 AND2_1144( .ZN(g15421), .A1(g4665), .A2(g12791) );
  AND2_X1 AND2_1145( .ZN(g15422), .A1(g4668), .A2(g12794) );
  AND2_X1 AND2_1146( .ZN(g15423), .A1(g4827), .A2(g13210) );
  AND2_X1 AND2_1147( .ZN(g15424), .A1(g4828), .A2(g13211) );
  AND2_X2 AND2_1148( .ZN(g15425), .A1(g4832), .A2(g13212) );
  AND2_X2 AND2_1149( .ZN(g15435), .A1(g4702), .A2(g12801) );
  AND2_X1 AND2_1150( .ZN(g15436), .A1(g4868), .A2(g13213) );
  AND2_X1 AND2_1151( .ZN(g15437), .A1(g4869), .A2(g13214) );
  AND2_X1 AND2_1152( .ZN(g15442), .A1(g2714), .A2(g12804) );
  AND2_X1 AND2_1153( .ZN(g15452), .A1(g7916), .A2(g12808) );
  AND2_X1 AND2_1154( .ZN(g15453), .A1(g6898), .A2(g12811) );
  AND2_X1 AND2_1155( .ZN(g15459), .A1(g4897), .A2(g13218) );
  AND2_X1 AND2_1156( .ZN(g15460), .A1(g4898), .A2(g13219) );
  AND2_X1 AND2_1157( .ZN(g15470), .A1(g4763), .A2(g12816) );
  AND2_X1 AND2_1158( .ZN(g15475), .A1(g4928), .A2(g13220) );
  AND2_X1 AND2_1159( .ZN(g15476), .A1(g4929), .A2(g13221) );
  AND2_X1 AND2_1160( .ZN(g15486), .A1(g4797), .A2(g12822) );
  AND2_X1 AND2_1161( .ZN(g15487), .A1(g4800), .A2(g12825) );
  AND2_X1 AND2_1162( .ZN(g15491), .A1(g4954), .A2(g13222) );
  AND2_X1 AND2_1163( .ZN(g15494), .A1(g4962), .A2(g13223) );
  AND2_X1 AND2_1164( .ZN(g15495), .A1(g4963), .A2(g13224) );
  AND2_X1 AND2_1165( .ZN(g15505), .A1(g4842), .A2(g12830) );
  AND2_X1 AND2_1166( .ZN(g15506), .A1(g4845), .A2(g12833) );
  AND2_X1 AND2_1167( .ZN(g15507), .A1(g5003), .A2(g13225) );
  AND2_X1 AND2_1168( .ZN(g15508), .A1(g5004), .A2(g13226) );
  AND2_X1 AND2_1169( .ZN(g15509), .A1(g5008), .A2(g13227) );
  AND2_X1 AND2_1170( .ZN(g15519), .A1(g4879), .A2(g12840) );
  AND2_X1 AND2_1171( .ZN(g15520), .A1(g8172), .A2(g12844) );
  AND2_X1 AND2_1172( .ZN(g15526), .A1(g5033), .A2(g13232) );
  AND2_X1 AND2_1173( .ZN(g15527), .A1(g5034), .A2(g13233) );
  AND2_X1 AND2_1174( .ZN(g15545), .A1(g5056), .A2(g13237) );
  AND2_X1 AND2_1175( .ZN(g15546), .A1(g5057), .A2(g13238) );
  AND2_X1 AND2_1176( .ZN(g15556), .A1(g4939), .A2(g12854) );
  AND2_X1 AND2_1177( .ZN(g15561), .A1(g5087), .A2(g13239) );
  AND2_X1 AND2_1178( .ZN(g15562), .A1(g5088), .A2(g13240) );
  AND2_X1 AND2_1179( .ZN(g15572), .A1(g4973), .A2(g12860) );
  AND2_X1 AND2_1180( .ZN(g15573), .A1(g4976), .A2(g12863) );
  AND2_X1 AND2_1181( .ZN(g15577), .A1(g5113), .A2(g13241) );
  AND2_X1 AND2_1182( .ZN(g15580), .A1(g5121), .A2(g13242) );
  AND2_X1 AND2_1183( .ZN(g15581), .A1(g5122), .A2(g13243) );
  AND2_X1 AND2_1184( .ZN(g15591), .A1(g5018), .A2(g12868) );
  AND2_X1 AND2_1185( .ZN(g15592), .A1(g5021), .A2(g12871) );
  AND2_X1 AND2_1186( .ZN(g15593), .A1(g7897), .A2(g13244) );
  AND2_X1 AND2_1187( .ZN(g15594), .A1(g5148), .A2(g13249) );
  AND2_X1 AND2_1188( .ZN(g15595), .A1(g5149), .A2(g13250) );
  AND2_X1 AND2_1189( .ZN(g15604), .A1(g5162), .A2(g13255) );
  AND2_X1 AND2_1190( .ZN(g15605), .A1(g5163), .A2(g13256) );
  AND2_X1 AND2_1191( .ZN(g15623), .A1(g5185), .A2(g13260) );
  AND2_X1 AND2_1192( .ZN(g15624), .A1(g5186), .A2(g13261) );
  AND2_X1 AND2_1193( .ZN(g15634), .A1(g5098), .A2(g12895) );
  AND2_X1 AND2_1194( .ZN(g15639), .A1(g5216), .A2(g13262) );
  AND2_X1 AND2_1195( .ZN(g15640), .A1(g5217), .A2(g13263) );
  AND2_X1 AND2_1196( .ZN(g15650), .A1(g5132), .A2(g12901) );
  AND2_X1 AND2_1197( .ZN(g15651), .A1(g5135), .A2(g12904) );
  AND2_X1 AND2_1198( .ZN(g15658), .A1(g8177), .A2(g13264) );
  AND2_X1 AND2_1199( .ZN(g15666), .A1(g5233), .A2(g13268) );
  AND2_X1 AND2_1200( .ZN(g15670), .A1(g5241), .A2(g13272) );
  AND2_X1 AND2_1201( .ZN(g15671), .A1(g5242), .A2(g13273) );
  AND2_X1 AND2_1202( .ZN(g15680), .A1(g5255), .A2(g13278) );
  AND2_X1 AND2_1203( .ZN(g15681), .A1(g5256), .A2(g13279) );
  AND2_X1 AND2_1204( .ZN(g15699), .A1(g5278), .A2(g13283) );
  AND2_X1 AND2_1205( .ZN(g15700), .A1(g5279), .A2(g13284) );
  AND2_X1 AND2_1206( .ZN(g15710), .A1(g5227), .A2(g12935) );
  AND2_X1 AND2_1207( .ZN(g15717), .A1(g7924), .A2(g13285) );
  AND2_X1 AND2_1208( .ZN(g15725), .A1(g5296), .A2(g13293) );
  AND2_X1 AND2_1209( .ZN(g15729), .A1(g5304), .A2(g13297) );
  AND2_X1 AND2_1210( .ZN(g15730), .A1(g5305), .A2(g13298) );
  AND2_X1 AND2_1211( .ZN(g15739), .A1(g5318), .A2(g13303) );
  AND2_X1 AND2_1212( .ZN(g15740), .A1(g5319), .A2(g13304) );
  AND2_X1 AND2_1213( .ZN(g15753), .A1(g7542), .A2(g12962) );
  AND2_X1 AND2_1214( .ZN(g15754), .A1(g7837), .A2(g13308) );
  AND2_X1 AND2_1215( .ZN(g15755), .A1(g8178), .A2(g13309) );
  AND2_X1 AND2_1216( .ZN(g15765), .A1(g5333), .A2(g13324) );
  AND2_X1 AND2_1217( .ZN(g15769), .A1(g5341), .A2(g13328) );
  AND2_X1 AND2_1218( .ZN(g15770), .A1(g5342), .A2(g13329) );
  AND3_X2 AND3_10( .ZN(II22028), .A1(g13004), .A2(g3018), .A3(g7549) );
  AND3_X4 AND3_11( .ZN(g15780), .A1(g7471), .A2(g3032), .A3(II22028) );
  AND2_X1 AND2_1219( .ZN(g15781), .A1(g7971), .A2(g13330) );
  AND2_X1 AND2_1220( .ZN(g15793), .A1(g5361), .A2(g13347) );
  AND2_X1 AND2_1221( .ZN(g15801), .A1(g7856), .A2(g13351) );
  AND2_X1 AND2_1222( .ZN(g15802), .A1(g8253), .A2(g13352) );
  AND2_X1 AND2_1223( .ZN(g15817), .A1(g8025), .A2(g13373) );
  AND2_X1 AND2_1224( .ZN(g15828), .A1(g7877), .A2(g13398) );
  AND2_X1 AND2_1225( .ZN(g15829), .A1(g7857), .A2(g13400) );
  AND2_X1 AND2_1226( .ZN(g15840), .A1(g8098), .A2(g11620) );
  AND2_X1 AND2_1227( .ZN(g15852), .A1(g7878), .A2(g11642) );
  AND3_X1 AND3_12( .ZN(II22136), .A1(g13082), .A2(g2912), .A3(g7522) );
  AND3_X1 AND3_13( .ZN(g15902), .A1(g7607), .A2(g2920), .A3(II22136) );
  AND2_X1 AND2_1228( .ZN(g15998), .A1(g5469), .A2(g11732) );
  AND2_X1 AND2_1229( .ZN(g16003), .A1(g12013), .A2(g10826) );
  AND2_X1 AND2_1230( .ZN(g16004), .A1(g5587), .A2(g11734) );
  AND2_X1 AND2_1231( .ZN(g16008), .A1(g5504), .A2(g11735) );
  AND2_X1 AND2_1232( .ZN(g16009), .A1(g12071), .A2(g10843) );
  AND2_X1 AND2_1233( .ZN(g16010), .A1(g7639), .A2(g11736) );
  AND2_X1 AND2_1234( .ZN(g16015), .A1(g12013), .A2(g10859) );
  AND2_X1 AND2_1235( .ZN(g16016), .A1(g5601), .A2(g11740) );
  AND2_X1 AND2_1236( .ZN(g16017), .A1(g12130), .A2(g10862) );
  AND2_X1 AND2_1237( .ZN(g16018), .A1(g6149), .A2(g11741) );
  AND2_X1 AND2_1238( .ZN(g16019), .A1(g5507), .A2(g11742) );
  AND2_X1 AND2_1239( .ZN(g16028), .A1(g5543), .A2(g11745) );
  AND2_X1 AND2_1240( .ZN(g16029), .A1(g12071), .A2(g10877) );
  AND2_X1 AND2_1241( .ZN(g16030), .A1(g7667), .A2(g11746) );
  AND2_X1 AND2_1242( .ZN(g16031), .A1(g6227), .A2(g11747) );
  AND2_X1 AND2_1243( .ZN(g16032), .A1(g12187), .A2(g10883) );
  AND2_X1 AND2_1244( .ZN(g16033), .A1(g5546), .A2(g11748) );
  AND2_X1 AND2_1245( .ZN(g16045), .A1(g12013), .A2(g10892) );
  AND2_X1 AND2_1246( .ZN(g16046), .A1(g5618), .A2(g11761) );
  AND2_X1 AND2_1247( .ZN(g16047), .A1(g12130), .A2(g10895) );
  AND2_X1 AND2_1248( .ZN(g16048), .A1(g6170), .A2(g11762) );
  AND2_X1 AND2_1249( .ZN(g16049), .A1(g6638), .A2(g11763) );
  AND2_X1 AND2_1250( .ZN(g16050), .A1(g5590), .A2(g11764) );
  AND2_X1 AND2_1251( .ZN(g16051), .A1(g12235), .A2(g10901) );
  AND2_X1 AND2_1252( .ZN(g16052), .A1(g5591), .A2(g11765) );
  AND2_X1 AND2_1253( .ZN(g16053), .A1(g297), .A2(g11770) );
  AND2_X1 AND2_1254( .ZN(g16066), .A1(g12071), .A2(g10912) );
  AND2_X1 AND2_1255( .ZN(g16067), .A1(g7700), .A2(g11774) );
  AND2_X1 AND2_1256( .ZN(g16068), .A1(g6310), .A2(g11775) );
  AND2_X1 AND2_1257( .ZN(g16069), .A1(g5346), .A2(g11776) );
  AND2_X1 AND2_1258( .ZN(g16070), .A1(g12187), .A2(g10921) );
  AND2_X1 AND2_1259( .ZN(g16071), .A1(g5604), .A2(g11777) );
  AND2_X1 AND2_1260( .ZN(g16072), .A1(g12275), .A2(g10924) );
  AND2_X1 AND2_1261( .ZN(g16073), .A1(g5605), .A2(g11778) );
  AND2_X1 AND2_1262( .ZN(g16074), .A1(g5646), .A2(g11782) );
  AND2_X1 AND2_1263( .ZN(g16081), .A1(g3304), .A2(g11783) );
  AND2_X1 AND2_1264( .ZN(g16089), .A1(g984), .A2(g11787) );
  AND2_X1 AND2_1265( .ZN(g16100), .A1(g12130), .A2(g10937) );
  AND2_X1 AND2_1266( .ZN(g16101), .A1(g6197), .A2(g11794) );
  AND2_X1 AND2_1267( .ZN(g16102), .A1(g6905), .A2(g11795) );
  AND2_X1 AND2_1268( .ZN(g16103), .A1(g5621), .A2(g11796) );
  AND2_X1 AND2_1269( .ZN(g16104), .A1(g12235), .A2(g10946) );
  AND2_X1 AND2_1270( .ZN(g16105), .A1(g5622), .A2(g11797) );
  AND2_X1 AND2_1271( .ZN(g16106), .A1(g12308), .A2(g10949) );
  AND2_X1 AND2_1272( .ZN(g16107), .A1(g5666), .A2(g11801) );
  AND2_X1 AND2_1273( .ZN(g16108), .A1(g5667), .A2(g11802) );
  AND2_X1 AND2_1274( .ZN(g16109), .A1(g8277), .A2(g11803) );
  AND2_X1 AND2_1275( .ZN(g16110), .A1(g516), .A2(g11804) );
  AND2_X1 AND2_1276( .ZN(g16111), .A1(g5551), .A2(g13215) );
  AND2_X1 AND2_1277( .ZN(g16112), .A1(g5684), .A2(g11808) );
  AND2_X1 AND2_1278( .ZN(g16119), .A1(g3460), .A2(g11809) );
  AND2_X1 AND2_1279( .ZN(g16127), .A1(g1678), .A2(g11813) );
  AND2_X1 AND2_1280( .ZN(g16133), .A1(g6444), .A2(g11817) );
  AND2_X1 AND2_1281( .ZN(g16134), .A1(g5363), .A2(g11818) );
  AND2_X1 AND2_1282( .ZN(g16135), .A1(g12187), .A2(g10980) );
  AND2_X1 AND2_1283( .ZN(g16136), .A1(g5640), .A2(g11819) );
  AND2_X1 AND2_1284( .ZN(g16137), .A1(g12275), .A2(g10983) );
  AND2_X1 AND2_1285( .ZN(g16138), .A1(g5641), .A2(g11820) );
  AND2_X1 AND2_1286( .ZN(g16139), .A1(g5704), .A2(g11824) );
  AND2_X1 AND2_1287( .ZN(g16140), .A1(g5705), .A2(g11825) );
  AND2_X1 AND2_1288( .ZN(g16141), .A1(g5706), .A2(g11826) );
  AND2_X1 AND2_1289( .ZN(g16152), .A1(g517), .A2(g11829) );
  AND2_X1 AND2_1290( .ZN(g16153), .A1(g5592), .A2(g13229) );
  AND2_X1 AND2_1291( .ZN(g16158), .A1(g5718), .A2(g11834) );
  AND2_X1 AND2_1292( .ZN(g16159), .A1(g5719), .A2(g11835) );
  AND2_X1 AND2_1293( .ZN(g16160), .A1(g8286), .A2(g11836) );
  AND2_X1 AND2_1294( .ZN(g16161), .A1(g1202), .A2(g11837) );
  AND2_X1 AND2_1295( .ZN(g16162), .A1(g5597), .A2(g13234) );
  AND2_X1 AND2_1296( .ZN(g16163), .A1(g5736), .A2(g11841) );
  AND2_X1 AND2_1297( .ZN(g16170), .A1(g3616), .A2(g11842) );
  AND2_X1 AND2_1298( .ZN(g16178), .A1(g2372), .A2(g11846) );
  AND2_X1 AND2_1299( .ZN(g16182), .A1(g7149), .A2(g11852) );
  AND2_X1 AND2_1300( .ZN(g16183), .A1(g12235), .A2(g11014) );
  AND2_X1 AND2_1301( .ZN(g16184), .A1(g5663), .A2(g11853) );
  AND2_X1 AND2_1302( .ZN(g16185), .A1(g12308), .A2(g11017) );
  AND2_X1 AND2_1303( .ZN(g16186), .A1(g5753), .A2(g11856) );
  AND2_X1 AND2_1304( .ZN(g16187), .A1(g5754), .A2(g11857) );
  AND2_X1 AND2_1305( .ZN(g16188), .A1(g5755), .A2(g11858) );
  AND2_X1 AND2_1306( .ZN(g16197), .A1(g518), .A2(g11862) );
  AND2_X1 AND2_1307( .ZN(g16198), .A1(g5762), .A2(g11866) );
  AND2_X1 AND2_1308( .ZN(g16199), .A1(g5763), .A2(g11867) );
  AND2_X1 AND2_1309( .ZN(g16200), .A1(g5764), .A2(g11868) );
  AND2_X1 AND2_1310( .ZN(g16211), .A1(g1203), .A2(g11871) );
  AND2_X1 AND2_1311( .ZN(g16212), .A1(g5609), .A2(g13252) );
  AND2_X1 AND2_1312( .ZN(g16217), .A1(g5776), .A2(g11876) );
  AND2_X1 AND2_1313( .ZN(g16218), .A1(g5777), .A2(g11877) );
  AND2_X1 AND2_1314( .ZN(g16219), .A1(g8295), .A2(g11878) );
  AND2_X1 AND2_1315( .ZN(g16220), .A1(g1896), .A2(g11879) );
  AND2_X1 AND2_1316( .ZN(g16221), .A1(g5614), .A2(g13257) );
  AND2_X1 AND2_1317( .ZN(g16222), .A1(g5794), .A2(g11883) );
  AND2_X1 AND2_1318( .ZN(g16229), .A1(g3772), .A2(g11884) );
  AND2_X1 AND2_1319( .ZN(g16237), .A1(g5379), .A2(g11886) );
  AND2_X2 AND2_1320( .ZN(g16238), .A1(g12275), .A2(g11066) );
  AND2_X2 AND2_1321( .ZN(g16239), .A1(g5700), .A2(g11887) );
  AND2_X2 AND2_1322( .ZN(g16240), .A1(g5804), .A2(g11891) );
  AND2_X1 AND2_1323( .ZN(g16241), .A1(g5805), .A2(g11892) );
  AND2_X1 AND2_1324( .ZN(g16242), .A1(g5806), .A2(g11893) );
  AND2_X1 AND2_1325( .ZN(g16250), .A1(g519), .A2(g11895) );
  AND2_X1 AND2_1326( .ZN(g16251), .A1(g5812), .A2(g11898) );
  AND2_X1 AND2_1327( .ZN(g16252), .A1(g5813), .A2(g11899) );
  AND2_X1 AND2_1328( .ZN(g16253), .A1(g5814), .A2(g11900) );
  AND2_X1 AND2_1329( .ZN(g16262), .A1(g1204), .A2(g11904) );
  AND2_X1 AND2_1330( .ZN(g16263), .A1(g5821), .A2(g11908) );
  AND2_X1 AND2_1331( .ZN(g16264), .A1(g5822), .A2(g11909) );
  AND2_X1 AND2_1332( .ZN(g16265), .A1(g5823), .A2(g11910) );
  AND2_X1 AND2_1333( .ZN(g16276), .A1(g1897), .A2(g11913) );
  AND2_X1 AND2_1334( .ZN(g16277), .A1(g5634), .A2(g13275) );
  AND2_X1 AND2_1335( .ZN(g16282), .A1(g5835), .A2(g11918) );
  AND2_X1 AND2_1336( .ZN(g16283), .A1(g5836), .A2(g11919) );
  AND2_X1 AND2_1337( .ZN(g16284), .A1(g8304), .A2(g11920) );
  AND2_X1 AND2_1338( .ZN(g16285), .A1(g2590), .A2(g11921) );
  AND2_X1 AND2_1339( .ZN(g16286), .A1(g5639), .A2(g13280) );
  AND2_X1 AND2_1340( .ZN(g16288), .A1(g12308), .A2(g11129) );
  AND2_X1 AND2_1341( .ZN(g16289), .A1(g5853), .A2(g11929) );
  AND2_X1 AND2_1342( .ZN(g16290), .A1(g5854), .A2(g11930) );
  AND2_X1 AND2_1343( .ZN(g16291), .A1(g5855), .A2(g11931) );
  AND2_X1 AND2_1344( .ZN(g16292), .A1(g294), .A2(g11932) );
  AND2_X1 AND2_1345( .ZN(g16298), .A1(g520), .A2(g11936) );
  AND2_X1 AND2_1346( .ZN(g16299), .A1(g5860), .A2(g11941) );
  AND2_X1 AND2_1347( .ZN(g16300), .A1(g5861), .A2(g11942) );
  AND2_X1 AND2_1348( .ZN(g16301), .A1(g5862), .A2(g11943) );
  AND2_X1 AND2_1349( .ZN(g16309), .A1(g1205), .A2(g11945) );
  AND2_X1 AND2_1350( .ZN(g16310), .A1(g5868), .A2(g11948) );
  AND2_X1 AND2_1351( .ZN(g16311), .A1(g5869), .A2(g11949) );
  AND2_X1 AND2_1352( .ZN(g16312), .A1(g5870), .A2(g11950) );
  AND2_X1 AND2_1353( .ZN(g16321), .A1(g1898), .A2(g11954) );
  AND2_X1 AND2_1354( .ZN(g16322), .A1(g5877), .A2(g11958) );
  AND2_X1 AND2_1355( .ZN(g16323), .A1(g5878), .A2(g11959) );
  AND2_X1 AND2_1356( .ZN(g16324), .A1(g5879), .A2(g11960) );
  AND2_X1 AND2_1357( .ZN(g16335), .A1(g2591), .A2(g11963) );
  AND2_X1 AND2_1358( .ZN(g16336), .A1(g5662), .A2(g13300) );
  AND2_X1 AND2_1359( .ZN(g16342), .A1(g5894), .A2(g11968) );
  AND2_X1 AND2_1360( .ZN(g16343), .A1(g5895), .A2(g11969) );
  AND2_X1 AND2_1361( .ZN(g16344), .A1(g5896), .A2(g11970) );
  AND2_X1 AND2_1362( .ZN(g16345), .A1(g5897), .A2(g11971) );
  AND2_X1 AND2_1363( .ZN(g16346), .A1(g295), .A2(g11972) );
  AND2_X1 AND2_1364( .ZN(g16347), .A1(g5900), .A2(g11982) );
  AND2_X1 AND2_1365( .ZN(g16348), .A1(g5901), .A2(g11983) );
  AND2_X1 AND2_1366( .ZN(g16349), .A1(g5902), .A2(g11984) );
  AND2_X1 AND2_1367( .ZN(g16350), .A1(g981), .A2(g11985) );
  AND2_X1 AND2_1368( .ZN(g16356), .A1(g1206), .A2(g11989) );
  AND2_X1 AND2_1369( .ZN(g16357), .A1(g5907), .A2(g11994) );
  AND2_X1 AND2_1370( .ZN(g16358), .A1(g5908), .A2(g11995) );
  AND2_X1 AND2_1371( .ZN(g16359), .A1(g5909), .A2(g11996) );
  AND2_X1 AND2_1372( .ZN(g16367), .A1(g1899), .A2(g11998) );
  AND2_X1 AND2_1373( .ZN(g16368), .A1(g5915), .A2(g12001) );
  AND2_X1 AND2_1374( .ZN(g16369), .A1(g5916), .A2(g12002) );
  AND2_X1 AND2_1375( .ZN(g16370), .A1(g5917), .A2(g12003) );
  AND2_X1 AND2_1376( .ZN(g16379), .A1(g2592), .A2(g12007) );
  AND2_X1 AND2_1377( .ZN(g16380), .A1(g5925), .A2(g12020) );
  AND2_X1 AND2_1378( .ZN(g16381), .A1(g5926), .A2(g12021) );
  AND2_X1 AND2_1379( .ZN(g16382), .A1(g5927), .A2(g12022) );
  AND2_X2 AND2_1380( .ZN(g16383), .A1(g5928), .A2(g12023) );
  AND2_X2 AND2_1381( .ZN(g16384), .A1(g296), .A2(g12024) );
  AND2_X1 AND2_1382( .ZN(g16385), .A1(g5714), .A2(g13336) );
  AND2_X1 AND2_1383( .ZN(g16386), .A1(g5933), .A2(g12037) );
  AND2_X1 AND2_1384( .ZN(g16387), .A1(g5934), .A2(g12038) );
  AND2_X1 AND2_1385( .ZN(g16388), .A1(g5935), .A2(g12039) );
  AND2_X1 AND2_1386( .ZN(g16389), .A1(g5936), .A2(g12040) );
  AND2_X1 AND2_1387( .ZN(g16390), .A1(g982), .A2(g12041) );
  AND2_X1 AND2_1388( .ZN(g16391), .A1(g5939), .A2(g12051) );
  AND2_X1 AND2_1389( .ZN(g16392), .A1(g5940), .A2(g12052) );
  AND2_X1 AND2_1390( .ZN(g16393), .A1(g5941), .A2(g12053) );
  AND2_X1 AND2_1391( .ZN(g16394), .A1(g1675), .A2(g12054) );
  AND2_X1 AND2_1392( .ZN(g16400), .A1(g1900), .A2(g12058) );
  AND2_X1 AND2_1393( .ZN(g16401), .A1(g5946), .A2(g12063) );
  AND2_X1 AND2_1394( .ZN(g16402), .A1(g5947), .A2(g12064) );
  AND2_X1 AND2_1395( .ZN(g16403), .A1(g5948), .A2(g12065) );
  AND2_X1 AND2_1396( .ZN(g16411), .A1(g2593), .A2(g12067) );
  AND2_X1 AND2_1397( .ZN(g16413), .A1(g5954), .A2(g12075) );
  AND2_X1 AND2_1398( .ZN(g16414), .A1(g5955), .A2(g12076) );
  AND2_X1 AND2_1399( .ZN(g16415), .A1(g5956), .A2(g12077) );
  AND2_X1 AND2_1400( .ZN(g16416), .A1(g5957), .A2(g12078) );
  AND2_X1 AND2_1401( .ZN(g16417), .A1(g5759), .A2(g13356) );
  AND2_X1 AND2_1402( .ZN(g16418), .A1(g5959), .A2(g12084) );
  AND2_X1 AND2_1403( .ZN(g16419), .A1(g5960), .A2(g12085) );
  AND2_X1 AND2_1404( .ZN(g16420), .A1(g5961), .A2(g12086) );
  AND2_X1 AND2_1405( .ZN(g16421), .A1(g5962), .A2(g12087) );
  AND2_X1 AND2_1406( .ZN(g16422), .A1(g983), .A2(g12088) );
  AND2_X1 AND2_1407( .ZN(g16423), .A1(g5772), .A2(g13361) );
  AND2_X1 AND2_1408( .ZN(g16424), .A1(g5967), .A2(g12101) );
  AND2_X1 AND2_1409( .ZN(g16425), .A1(g5968), .A2(g12102) );
  AND2_X1 AND2_1410( .ZN(g16426), .A1(g5969), .A2(g12103) );
  AND2_X1 AND2_1411( .ZN(g16427), .A1(g5970), .A2(g12104) );
  AND2_X1 AND2_1412( .ZN(g16428), .A1(g1676), .A2(g12105) );
  AND2_X1 AND2_1413( .ZN(g16429), .A1(g5973), .A2(g12115) );
  AND2_X1 AND2_1414( .ZN(g16430), .A1(g5974), .A2(g12116) );
  AND2_X1 AND2_1415( .ZN(g16431), .A1(g5975), .A2(g12117) );
  AND2_X1 AND2_1416( .ZN(g16432), .A1(g2369), .A2(g12118) );
  AND2_X1 AND2_1417( .ZN(g16438), .A1(g2594), .A2(g12122) );
  AND2_X1 AND2_1418( .ZN(g16443), .A1(g5980), .A2(g12134) );
  AND2_X1 AND2_1419( .ZN(g16444), .A1(g5981), .A2(g12135) );
  AND2_X1 AND2_1420( .ZN(g16445), .A1(g5808), .A2(g13381) );
  AND2_X1 AND2_1421( .ZN(g16447), .A1(g5983), .A2(g12147) );
  AND2_X1 AND2_1422( .ZN(g16448), .A1(g5984), .A2(g12148) );
  AND2_X1 AND2_1423( .ZN(g16449), .A1(g5985), .A2(g12149) );
  AND2_X1 AND2_1424( .ZN(g16450), .A1(g5986), .A2(g12150) );
  AND2_X1 AND2_1425( .ZN(g16451), .A1(g5818), .A2(g13386) );
  AND2_X1 AND2_1426( .ZN(g16452), .A1(g5988), .A2(g12156) );
  AND2_X1 AND2_1427( .ZN(g16453), .A1(g5989), .A2(g12157) );
  AND2_X1 AND2_1428( .ZN(g16454), .A1(g5990), .A2(g12158) );
  AND2_X1 AND2_1429( .ZN(g16455), .A1(g5991), .A2(g12159) );
  AND2_X1 AND2_1430( .ZN(g16456), .A1(g1677), .A2(g12160) );
  AND2_X1 AND2_1431( .ZN(g16457), .A1(g5831), .A2(g13391) );
  AND2_X1 AND2_1432( .ZN(g16458), .A1(g5996), .A2(g12173) );
  AND2_X1 AND2_1433( .ZN(g16459), .A1(g5997), .A2(g12174) );
  AND2_X1 AND2_1434( .ZN(g16460), .A1(g5998), .A2(g12175) );
  AND2_X1 AND2_1435( .ZN(g16461), .A1(g5999), .A2(g12176) );
  AND2_X1 AND2_1436( .ZN(g16462), .A1(g2370), .A2(g12177) );
  AND4_X1 AND4_22( .ZN(g16505), .A1(g14776), .A2(g14797), .A3(g16142), .A4(g16243) );
  AND4_X1 AND4_23( .ZN(g16513), .A1(g15065), .A2(g13724), .A3(g13764), .A4(g13797) );
  AND4_X1 AND4_24( .ZN(g16527), .A1(g14811), .A2(g14849), .A3(g16201), .A4(g16302) );
  AND4_X1 AND4_25( .ZN(g16535), .A1(g15161), .A2(g13774), .A3(g13805), .A4(g13825) );
  AND4_X1 AND4_26( .ZN(g16558), .A1(g14863), .A2(g14922), .A3(g16266), .A4(g16360) );
  AND4_X1 AND4_27( .ZN(g16590), .A1(g14936), .A2(g15003), .A3(g16325), .A4(g16404) );
  AND2_X1 AND2_1437( .ZN(g16607), .A1(g15022), .A2(g15096) );
  AND2_X1 AND2_1438( .ZN(g16625), .A1(g15118), .A2(g15188) );
  AND2_X1 AND2_1439( .ZN(g16639), .A1(g15210), .A2(g15274) );
  AND2_X1 AND2_1440( .ZN(g16650), .A1(g15296), .A2(g15366) );
  AND2_X1 AND2_1441( .ZN(g16850), .A1(g6226), .A2(g14764) );
  AND2_X1 AND2_1442( .ZN(g16855), .A1(g15722), .A2(g8646) );
  AND2_X1 AND2_1443( .ZN(g16856), .A1(g6443), .A2(g14794) );
  AND2_X1 AND2_1444( .ZN(g16859), .A1(g15762), .A2(g8662) );
  AND2_X1 AND2_1445( .ZN(g16864), .A1(g15790), .A2(g8681) );
  AND2_X1 AND2_1446( .ZN(g16865), .A1(g6896), .A2(g14881) );
  AND2_X1 AND2_1447( .ZN(g16879), .A1(g15813), .A2(g8693) );
  AND2_X1 AND2_1448( .ZN(g16894), .A1(g7156), .A2(g14959) );
  AND2_X1 AND2_1449( .ZN(g16907), .A1(g7335), .A2(g15017) );
  AND2_X1 AND2_1450( .ZN(g16908), .A1(g7838), .A2(g15032) );
  AND2_X1 AND2_1451( .ZN(g16909), .A1(g6908), .A2(g15033) );
  AND2_X1 AND2_1452( .ZN(g16923), .A1(g7352), .A2(g15048) );
  AND2_X1 AND2_1453( .ZN(g16938), .A1(g7858), .A2(g15128) );
  AND2_X1 AND2_1454( .ZN(g16939), .A1(g7158), .A2(g15129) );
  AND2_X1 AND2_1455( .ZN(g16953), .A1(g7482), .A2(g15144) );
  AND2_X1 AND2_1456( .ZN(g16964), .A1(g7520), .A2(g15170) );
  AND2_X1 AND2_1457( .ZN(g16966), .A1(g7529), .A2(g15174) );
  AND2_X1 AND2_1458( .ZN(g16967), .A1(g7827), .A2(g15175) );
  AND2_X1 AND2_1459( .ZN(g16968), .A1(g6672), .A2(g15176) );
  AND2_X1 AND2_1460( .ZN(g16969), .A1(g7888), .A2(g15220) );
  AND2_X1 AND2_1461( .ZN(g16970), .A1(g7354), .A2(g15221) );
  AND2_X1 AND2_1462( .ZN(g16984), .A1(g7538), .A2(g15236) );
  AND2_X1 AND2_1463( .ZN(g16987), .A1(g7555), .A2(g15260) );
  AND2_X1 AND2_1464( .ZN(g16988), .A1(g7842), .A2(g15261) );
  AND2_X1 AND2_1465( .ZN(g16989), .A1(g6974), .A2(g15262) );
  AND2_X1 AND2_1466( .ZN(g16990), .A1(g7912), .A2(g15306) );
  AND2_X1 AND2_1467( .ZN(g16991), .A1(g7484), .A2(g15307) );
  AND2_X1 AND2_1468( .ZN(g16993), .A1(g7576), .A2(g15322) );
  AND2_X1 AND2_1469( .ZN(g16994), .A1(g7819), .A2(g15323) );
  AND2_X1 AND2_1470( .ZN(g16997), .A1(g7578), .A2(g15352) );
  AND2_X1 AND2_1471( .ZN(g16998), .A1(g7862), .A2(g15353) );
  AND2_X1 AND2_1472( .ZN(g16999), .A1(g7224), .A2(g15354) );
  AND3_X1 AND3_14( .ZN(g17001), .A1(g3254), .A2(g10694), .A3(g14144) );
  AND2_X1 AND2_1473( .ZN(g17015), .A1(g7996), .A2(g15390) );
  AND2_X1 AND2_1474( .ZN(g17017), .A1(g7590), .A2(g15408) );
  AND2_X1 AND2_1475( .ZN(g17018), .A1(g7830), .A2(g15409) );
  AND2_X1 AND2_1476( .ZN(g17021), .A1(g7592), .A2(g15438) );
  AND2_X1 AND2_1477( .ZN(g17022), .A1(g7892), .A2(g15439) );
  AND2_X1 AND2_1478( .ZN(g17023), .A1(g7420), .A2(g15440) );
  AND2_X1 AND2_1479( .ZN(g17028), .A1(g7604), .A2(g15458) );
  AND3_X1 AND3_15( .ZN(g17031), .A1(g3410), .A2(g10714), .A3(g14259) );
  AND2_X1 AND2_1480( .ZN(g17045), .A1(g8071), .A2(g15474) );
  AND2_X1 AND2_1481( .ZN(g17047), .A1(g7605), .A2(g15492) );
  AND2_X1 AND2_1482( .ZN(g17048), .A1(g7845), .A2(g15493) );
  AND2_X1 AND2_1483( .ZN(g17055), .A1(g7153), .A2(g15524) );
  AND2_X1 AND2_1484( .ZN(g17056), .A1(g7953), .A2(g15525) );
  AND2_X1 AND2_1485( .ZN(g17062), .A1(g7613), .A2(g15544) );
  AND3_X1 AND3_16( .ZN(g17065), .A1(g3566), .A2(g10735), .A3(g14381) );
  AND2_X1 AND2_1486( .ZN(g17079), .A1(g8156), .A2(g15560) );
  AND2_X1 AND2_1487( .ZN(g17081), .A1(g7614), .A2(g15578) );
  AND2_X1 AND2_1488( .ZN(g17082), .A1(g7865), .A2(g15579) );
  AND2_X1 AND2_1489( .ZN(g17084), .A1(g7629), .A2(g13954) );
  AND2_X1 AND2_1490( .ZN(g17090), .A1(g7349), .A2(g15602) );
  AND2_X1 AND2_1491( .ZN(g17091), .A1(g8004), .A2(g15603) );
  AND2_X1 AND2_1492( .ZN(g17097), .A1(g7622), .A2(g15622) );
  AND3_X1 AND3_17( .ZN(g17100), .A1(g3722), .A2(g10754), .A3(g14493) );
  AND2_X1 AND2_1493( .ZN(g17114), .A1(g8242), .A2(g15638) );
  AND2_X1 AND2_1494( .ZN(g17116), .A1(g7649), .A2(g14008) );
  AND2_X1 AND2_1495( .ZN(g17117), .A1(g7906), .A2(g15665) );
  AND2_X1 AND2_1496( .ZN(g17122), .A1(g7658), .A2(g14024) );
  AND2_X1 AND2_1497( .ZN(g17128), .A1(g7479), .A2(g15678) );
  AND2_X1 AND2_1498( .ZN(g17129), .A1(g8079), .A2(g15679) );
  AND2_X1 AND2_1499( .ZN(g17135), .A1(g7638), .A2(g15698) );
  AND2_X1 AND2_1500( .ZN(g17138), .A1(g7676), .A2(g14068) );
  AND2_X1 AND2_1501( .ZN(g17143), .A1(g7685), .A2(g14099) );
  AND2_X1 AND2_1502( .ZN(g17144), .A1(g7958), .A2(g15724) );
  AND2_X1 AND2_1503( .ZN(g17149), .A1(g7694), .A2(g14115) );
  AND2_X1 AND2_1504( .ZN(g17155), .A1(g7535), .A2(g15737) );
  AND2_X1 AND2_1505( .ZN(g17156), .A1(g8164), .A2(g15738) );
  AND2_X1 AND2_1506( .ZN(g17161), .A1(g7712), .A2(g14183) );
  AND2_X1 AND2_1507( .ZN(g17166), .A1(g7721), .A2(g14214) );
  AND2_X1 AND2_1508( .ZN(g17167), .A1(g8009), .A2(g15764) );
  AND2_X1 AND2_1509( .ZN(g17172), .A1(g7730), .A2(g14230) );
  AND2_X1 AND2_1510( .ZN(g17176), .A1(g7742), .A2(g14298) );
  AND2_X1 AND2_1511( .ZN(g17181), .A1(g7751), .A2(g14329) );
  AND2_X1 AND2_1512( .ZN(g17182), .A1(g8084), .A2(g15792) );
  AND2_X1 AND2_1513( .ZN(g17193), .A1(g7766), .A2(g14420) );
  AND2_X1 AND2_1514( .ZN(g17268), .A1(g8024), .A2(g15991) );
  AND2_X1 AND2_1515( .ZN(g17301), .A1(g8097), .A2(g15994) );
  AND2_X1 AND2_1516( .ZN(g17339), .A1(g8176), .A2(g15997) );
  AND2_X1 AND2_1517( .ZN(g17352), .A1(g3942), .A2(g14960) );
  AND2_X1 AND2_1518( .ZN(g17353), .A1(g3945), .A2(g14963) );
  AND2_X1 AND2_1519( .ZN(g17381), .A1(g8250), .A2(g16001) );
  AND2_X1 AND2_1520( .ZN(g17382), .A1(g8252), .A2(g16002) );
  AND2_X1 AND2_1521( .ZN(g17393), .A1(g3941), .A2(g16005) );
  AND2_X1 AND2_1522( .ZN(g17395), .A1(g6177), .A2(g15034) );
  AND2_X1 AND2_1523( .ZN(g17396), .A1(g4020), .A2(g15037) );
  AND2_X1 AND2_1524( .ZN(g17397), .A1(g4023), .A2(g15040) );
  AND2_X1 AND2_1525( .ZN(g17398), .A1(g4026), .A2(g15043) );
  AND2_X1 AND2_1526( .ZN(g17408), .A1(g4049), .A2(g15049) );
  AND2_X1 AND2_1527( .ZN(g17409), .A1(g4052), .A2(g15052) );
  AND2_X1 AND2_1528( .ZN(g17428), .A1(g3994), .A2(g16007) );
  AND2_X1 AND2_1529( .ZN(g17446), .A1(g6284), .A2(g16011) );
  AND2_X1 AND2_1530( .ZN(g17447), .A1(g4115), .A2(g15106) );
  AND2_X1 AND2_1531( .ZN(g17448), .A1(g4118), .A2(g15109) );
  AND2_X1 AND2_1532( .ZN(g17449), .A1(g4121), .A2(g15112) );
  AND2_X1 AND2_1533( .ZN(g17450), .A1(g4124), .A2(g15115) );
  AND2_X1 AND2_1534( .ZN(g17460), .A1(g4048), .A2(g16012) );
  AND2_X1 AND2_1535( .ZN(g17461), .A1(g6209), .A2(g15130) );
  AND2_X1 AND2_1536( .ZN(g17462), .A1(g4147), .A2(g15133) );
  AND2_X1 AND2_1537( .ZN(g17463), .A1(g4150), .A2(g15136) );
  AND2_X1 AND2_1538( .ZN(g17464), .A1(g4153), .A2(g15139) );
  AND2_X1 AND2_1539( .ZN(g17474), .A1(g4176), .A2(g15145) );
  AND2_X1 AND2_1540( .ZN(g17475), .A1(g4179), .A2(g15148) );
  AND2_X1 AND2_1541( .ZN(g17485), .A1(g4089), .A2(g16013) );
  AND2_X1 AND2_1542( .ZN(g17486), .A1(g4091), .A2(g16014) );
  AND2_X1 AND2_1543( .ZN(g17506), .A1(g6675), .A2(g16023) );
  AND2_X1 AND2_1544( .ZN(g17508), .A1(g4225), .A2(g15179) );
  AND2_X1 AND2_1545( .ZN(g17509), .A1(g4228), .A2(g15182) );
  AND2_X1 AND2_1546( .ZN(g17510), .A1(g4231), .A2(g15185) );
  AND2_X1 AND2_1547( .ZN(g17526), .A1(g6421), .A2(g16025) );
  AND2_X1 AND2_1548( .ZN(g17527), .A1(g4254), .A2(g15198) );
  AND2_X1 AND2_1549( .ZN(g17528), .A1(g4257), .A2(g15201) );
  AND2_X1 AND2_1550( .ZN(g17529), .A1(g4260), .A2(g15204) );
  AND2_X1 AND2_1551( .ZN(g17530), .A1(g4263), .A2(g15207) );
  AND2_X1 AND2_1552( .ZN(g17540), .A1(g4175), .A2(g16026) );
  AND2_X1 AND2_1553( .ZN(g17541), .A1(g6298), .A2(g15222) );
  AND2_X1 AND2_1554( .ZN(g17542), .A1(g4286), .A2(g15225) );
  AND2_X1 AND2_1555( .ZN(g17543), .A1(g4289), .A2(g15228) );
  AND2_X1 AND2_1556( .ZN(g17544), .A1(g4292), .A2(g15231) );
  AND2_X1 AND2_1557( .ZN(g17554), .A1(g4315), .A2(g15237) );
  AND2_X1 AND2_1558( .ZN(g17555), .A1(g4318), .A2(g15240) );
  AND2_X1 AND2_1559( .ZN(g17556), .A1(g4201), .A2(g16027) );
  AND2_X1 AND2_1560( .ZN(g17576), .A1(g4348), .A2(g15248) );
  AND2_X1 AND2_1561( .ZN(g17577), .A1(g4351), .A2(g15251) );
  AND2_X1 AND2_1562( .ZN(g17578), .A1(g4354), .A2(g15254) );
  AND2_X1 AND2_1563( .ZN(g17597), .A1(g6977), .A2(g16039) );
  AND2_X1 AND2_1564( .ZN(g17598), .A1(g4380), .A2(g15265) );
  AND2_X1 AND2_1565( .ZN(g17599), .A1(g4383), .A2(g15268) );
  AND2_X1 AND2_1566( .ZN(g17600), .A1(g4386), .A2(g15271) );
  AND2_X1 AND2_1567( .ZN(g17616), .A1(g6626), .A2(g16041) );
  AND2_X1 AND2_1568( .ZN(g17617), .A1(g4409), .A2(g15284) );
  AND2_X1 AND2_1569( .ZN(g17618), .A1(g4412), .A2(g15287) );
  AND2_X1 AND2_1570( .ZN(g17619), .A1(g4415), .A2(g15290) );
  AND2_X1 AND2_1571( .ZN(g17620), .A1(g4418), .A2(g15293) );
  AND2_X1 AND2_1572( .ZN(g17630), .A1(g4314), .A2(g16042) );
  AND2_X1 AND2_1573( .ZN(g17631), .A1(g6435), .A2(g15308) );
  AND2_X1 AND2_1574( .ZN(g17632), .A1(g4441), .A2(g15311) );
  AND2_X1 AND2_1575( .ZN(g17633), .A1(g4444), .A2(g15314) );
  AND2_X1 AND2_1576( .ZN(g17634), .A1(g4447), .A2(g15317) );
  AND2_X1 AND2_1577( .ZN(g17635), .A1(g4322), .A2(g16043) );
  AND2_X1 AND2_1578( .ZN(g17636), .A1(g4324), .A2(g16044) );
  AND2_X1 AND2_1579( .ZN(g17652), .A1(g4480), .A2(g15326) );
  AND2_X1 AND2_1580( .ZN(g17653), .A1(g4483), .A2(g15329) );
  AND2_X1 AND2_1581( .ZN(g17654), .A1(g4486), .A2(g15332) );
  AND2_X1 AND2_1582( .ZN(g17673), .A1(g4517), .A2(g15340) );
  AND2_X1 AND2_1583( .ZN(g17674), .A1(g4520), .A2(g15343) );
  AND2_X1 AND2_1584( .ZN(g17675), .A1(g4523), .A2(g15346) );
  AND2_X1 AND2_1585( .ZN(g17694), .A1(g7227), .A2(g16061) );
  AND2_X1 AND2_1586( .ZN(g17695), .A1(g4549), .A2(g15357) );
  AND2_X1 AND2_1587( .ZN(g17696), .A1(g4552), .A2(g15360) );
  AND2_X1 AND2_1588( .ZN(g17697), .A1(g4555), .A2(g15363) );
  AND2_X1 AND2_1589( .ZN(g17713), .A1(g6890), .A2(g16063) );
  AND2_X1 AND2_1590( .ZN(g17714), .A1(g4578), .A2(g15376) );
  AND2_X1 AND2_1591( .ZN(g17715), .A1(g4581), .A2(g15379) );
  AND2_X1 AND2_1592( .ZN(g17716), .A1(g4584), .A2(g15382) );
  AND2_X1 AND2_1593( .ZN(g17717), .A1(g4587), .A2(g15385) );
  AND2_X1 AND2_1594( .ZN(g17718), .A1(g4451), .A2(g16064) );
  AND2_X1 AND2_1595( .ZN(g17719), .A1(g2993), .A2(g16065) );
  AND2_X1 AND2_1596( .ZN(g17734), .A1(g4611), .A2(g15393) );
  AND2_X1 AND2_1597( .ZN(g17735), .A1(g4614), .A2(g15396) );
  AND2_X1 AND2_1598( .ZN(g17736), .A1(g4617), .A2(g15399) );
  AND2_X1 AND2_1599( .ZN(g17737), .A1(g4626), .A2(g15404) );
  AND2_X2 AND2_1600( .ZN(g17752), .A1(g4656), .A2(g15412) );
  AND2_X2 AND2_1601( .ZN(g17753), .A1(g4659), .A2(g15415) );
  AND2_X2 AND2_1602( .ZN(g17754), .A1(g4662), .A2(g15418) );
  AND2_X2 AND2_1603( .ZN(g17773), .A1(g4693), .A2(g15426) );
  AND2_X2 AND2_1604( .ZN(g17774), .A1(g4696), .A2(g15429) );
  AND2_X2 AND2_1605( .ZN(g17775), .A1(g4699), .A2(g15432) );
  AND2_X1 AND2_1606( .ZN(g17794), .A1(g7423), .A2(g16097) );
  AND2_X1 AND2_1607( .ZN(g17795), .A1(g4725), .A2(g15443) );
  AND2_X1 AND2_1608( .ZN(g17796), .A1(g4728), .A2(g15446) );
  AND2_X1 AND2_1609( .ZN(g17797), .A1(g4731), .A2(g15449) );
  AND2_X1 AND2_1610( .ZN(g17798), .A1(g4591), .A2(g16099) );
  AND2_X1 AND2_1611( .ZN(g17812), .A1(g4754), .A2(g15461) );
  AND2_X1 AND2_1612( .ZN(g17813), .A1(g4757), .A2(g15464) );
  AND2_X1 AND2_1613( .ZN(g17814), .A1(g4760), .A2(g15467) );
  AND2_X1 AND2_1614( .ZN(g17824), .A1(g4766), .A2(g15471) );
  AND2_X1 AND2_1615( .ZN(g17835), .A1(g4788), .A2(g15477) );
  AND2_X1 AND2_1616( .ZN(g17836), .A1(g4791), .A2(g15480) );
  AND2_X1 AND2_1617( .ZN(g17837), .A1(g4794), .A2(g15483) );
  AND2_X1 AND2_1618( .ZN(g17838), .A1(g4803), .A2(g15488) );
  AND2_X1 AND2_1619( .ZN(g17853), .A1(g4833), .A2(g15496) );
  AND2_X1 AND2_1620( .ZN(g17854), .A1(g4836), .A2(g15499) );
  AND2_X1 AND2_1621( .ZN(g17855), .A1(g4839), .A2(g15502) );
  AND2_X1 AND2_1622( .ZN(g17874), .A1(g4870), .A2(g15510) );
  AND2_X1 AND2_1623( .ZN(g17875), .A1(g4873), .A2(g15513) );
  AND2_X1 AND2_1624( .ZN(g17876), .A1(g4876), .A2(g15516) );
  AND2_X1 AND2_1625( .ZN(g17877), .A1(g2998), .A2(g15521) );
  AND2_X1 AND2_1626( .ZN(g17900), .A1(g4899), .A2(g15528) );
  AND2_X1 AND2_1627( .ZN(g17901), .A1(g4902), .A2(g15531) );
  AND2_X1 AND2_1628( .ZN(g17902), .A1(g4905), .A2(g15534) );
  AND2_X1 AND2_1629( .ZN(g17912), .A1(g4908), .A2(g15537) );
  AND2_X1 AND2_1630( .ZN(g17924), .A1(g4930), .A2(g15547) );
  AND2_X1 AND2_1631( .ZN(g17925), .A1(g4933), .A2(g15550) );
  AND2_X1 AND2_1632( .ZN(g17926), .A1(g4936), .A2(g15553) );
  AND2_X1 AND2_1633( .ZN(g17936), .A1(g4942), .A2(g15557) );
  AND2_X1 AND2_1634( .ZN(g17947), .A1(g4964), .A2(g15563) );
  AND2_X1 AND2_1635( .ZN(g17948), .A1(g4967), .A2(g15566) );
  AND2_X1 AND2_1636( .ZN(g17949), .A1(g4970), .A2(g15569) );
  AND2_X1 AND2_1637( .ZN(g17950), .A1(g4979), .A2(g15574) );
  AND2_X1 AND2_1638( .ZN(g17965), .A1(g5009), .A2(g15582) );
  AND2_X1 AND2_1639( .ZN(g17966), .A1(g5012), .A2(g15585) );
  AND2_X1 AND2_1640( .ZN(g17967), .A1(g5015), .A2(g15588) );
  AND2_X1 AND2_1641( .ZN(g17989), .A1(g5035), .A2(g15596) );
  AND2_X1 AND2_1642( .ZN(g17990), .A1(g5038), .A2(g15599) );
  AND2_X1 AND2_1643( .ZN(g18011), .A1(g5058), .A2(g15606) );
  AND2_X1 AND2_1644( .ZN(g18012), .A1(g5061), .A2(g15609) );
  AND2_X1 AND2_1645( .ZN(g18013), .A1(g5064), .A2(g15612) );
  AND2_X1 AND2_1646( .ZN(g18023), .A1(g5067), .A2(g15615) );
  AND2_X1 AND2_1647( .ZN(g18035), .A1(g5089), .A2(g15625) );
  AND2_X1 AND2_1648( .ZN(g18036), .A1(g5092), .A2(g15628) );
  AND2_X1 AND2_1649( .ZN(g18037), .A1(g5095), .A2(g15631) );
  AND2_X1 AND2_1650( .ZN(g18047), .A1(g5101), .A2(g15635) );
  AND2_X1 AND2_1651( .ZN(g18058), .A1(g5123), .A2(g15641) );
  AND2_X1 AND2_1652( .ZN(g18059), .A1(g5126), .A2(g15644) );
  AND2_X1 AND2_1653( .ZN(g18060), .A1(g5129), .A2(g15647) );
  AND2_X1 AND2_1654( .ZN(g18061), .A1(g5138), .A2(g15652) );
  AND2_X1 AND2_1655( .ZN(g18062), .A1(g7462), .A2(g15655) );
  AND2_X1 AND2_1656( .ZN(g18088), .A1(g5150), .A2(g15667) );
  AND2_X1 AND2_1657( .ZN(g18106), .A1(g5164), .A2(g15672) );
  AND2_X1 AND2_1658( .ZN(g18107), .A1(g5167), .A2(g15675) );
  AND2_X1 AND2_1659( .ZN(g18128), .A1(g5187), .A2(g15682) );
  AND2_X1 AND2_1660( .ZN(g18129), .A1(g5190), .A2(g15685) );
  AND2_X1 AND2_1661( .ZN(g18130), .A1(g5193), .A2(g15688) );
  AND2_X1 AND2_1662( .ZN(g18140), .A1(g5196), .A2(g15691) );
  AND2_X1 AND2_1663( .ZN(g18152), .A1(g5218), .A2(g15701) );
  AND2_X1 AND2_1664( .ZN(g18153), .A1(g5221), .A2(g15704) );
  AND2_X1 AND2_1665( .ZN(g18154), .A1(g5224), .A2(g15707) );
  AND2_X1 AND2_1666( .ZN(g18164), .A1(g5230), .A2(g15711) );
  AND2_X1 AND2_1667( .ZN(g18165), .A1(g2883), .A2(g16287) );
  AND2_X1 AND2_1668( .ZN(g18169), .A1(g7527), .A2(g15714) );
  AND2_X1 AND2_1669( .ZN(g18204), .A1(g5243), .A2(g15726) );
  AND2_X1 AND2_1670( .ZN(g18222), .A1(g5257), .A2(g15731) );
  AND2_X1 AND2_1671( .ZN(g18223), .A1(g5260), .A2(g15734) );
  AND2_X1 AND2_1672( .ZN(g18244), .A1(g5280), .A2(g15741) );
  AND2_X1 AND2_1673( .ZN(g18245), .A1(g5283), .A2(g15744) );
  AND2_X1 AND2_1674( .ZN(g18246), .A1(g5286), .A2(g15747) );
  AND2_X1 AND2_1675( .ZN(g18256), .A1(g5289), .A2(g15750) );
  AND2_X1 AND2_1676( .ZN(g18311), .A1(g5306), .A2(g15766) );
  AND2_X1 AND2_1677( .ZN(g18329), .A1(g5320), .A2(g15771) );
  AND2_X1 AND2_1678( .ZN(g18330), .A1(g5323), .A2(g15774) );
  AND2_X1 AND2_1679( .ZN(g18333), .A1(g2888), .A2(g15777) );
  AND2_X1 AND2_1680( .ZN(g18404), .A1(g5343), .A2(g15794) );
  AND3_X1 AND3_18( .ZN(II24619), .A1(g14776), .A2(g14837), .A3(g16142) );
  AND3_X1 AND3_19( .ZN(g18547), .A1(g13677), .A2(g13750), .A3(II24619) );
  AND3_X1 AND3_20( .ZN(II24689), .A1(g14811), .A2(g14910), .A3(g16201) );
  AND3_X1 AND3_21( .ZN(g18597), .A1(g13714), .A2(g13791), .A3(II24689) );
  AND3_X1 AND3_22( .ZN(II24738), .A1(g14863), .A2(g14991), .A3(g16266) );
  AND3_X1 AND3_23( .ZN(g18629), .A1(g13764), .A2(g13819), .A3(II24738) );
  AND3_X1 AND3_24( .ZN(II24758), .A1(g14936), .A2(g15080), .A3(g16325) );
  AND3_X1 AND3_25( .ZN(g18638), .A1(g13805), .A2(g13840), .A3(II24758) );
  AND4_X1 AND4_28( .ZN(g18645), .A1(g14776), .A2(g14895), .A3(g16142), .A4(g13750) );
  AND3_X1 AND3_26( .ZN(g18647), .A1(g14895), .A2(g16142), .A3(g16243) );
  AND4_X1 AND4_29( .ZN(g18648), .A1(g14811), .A2(g14976), .A3(g16201), .A4(g13791) );
  AND4_X2 AND4_30( .ZN(g18649), .A1(g14776), .A2(g14837), .A3(g13657), .A4(g16189) );
  AND3_X1 AND3_27( .ZN(g18650), .A1(g14976), .A2(g16201), .A3(g16302) );
  AND4_X1 AND4_31( .ZN(g18651), .A1(g14863), .A2(g15065), .A3(g16266), .A4(g13819) );
  AND4_X1 AND4_32( .ZN(g18652), .A1(g14797), .A2(g13657), .A3(g13677), .A4(g16243) );
  AND4_X1 AND4_33( .ZN(g18653), .A1(g14811), .A2(g14910), .A3(g13687), .A4(g16254) );
  AND3_X1 AND3_28( .ZN(g18654), .A1(g15065), .A2(g16266), .A3(g16360) );
  AND4_X1 AND4_34( .ZN(g18655), .A1(g14936), .A2(g15161), .A3(g16325), .A4(g13840) );
  AND4_X1 AND4_35( .ZN(g18665), .A1(g14776), .A2(g14837), .A3(g16189), .A4(g13706) );
  AND4_X1 AND4_36( .ZN(g18666), .A1(g14849), .A2(g13687), .A3(g13714), .A4(g16302) );
  AND4_X2 AND4_37( .ZN(g18667), .A1(g14863), .A2(g14991), .A3(g13724), .A4(g16313) );
  AND3_X1 AND3_29( .ZN(g18668), .A1(g15161), .A2(g16325), .A3(g16404) );
  AND4_X1 AND4_38( .ZN(g18688), .A1(g14811), .A2(g14910), .A3(g16254), .A4(g13756) );
  AND4_X1 AND4_39( .ZN(g18689), .A1(g14922), .A2(g13724), .A3(g13764), .A4(g16360) );
  AND4_X1 AND4_40( .ZN(g18690), .A1(g14936), .A2(g15080), .A3(g13774), .A4(g16371) );
  AND4_X1 AND4_41( .ZN(g18717), .A1(g14863), .A2(g14991), .A3(g16313), .A4(g13797) );
  AND4_X1 AND4_42( .ZN(g18718), .A1(g15003), .A2(g13774), .A3(g13805), .A4(g16404) );
  AND4_X1 AND4_43( .ZN(g18753), .A1(g14936), .A2(g15080), .A3(g16371), .A4(g13825) );
  AND2_X1 AND2_1681( .ZN(g18982), .A1(g13519), .A2(g16154) );
  AND2_X1 AND2_1682( .ZN(g18990), .A1(g13530), .A2(g16213) );
  AND4_X1 AND4_44( .ZN(g18994), .A1(g14895), .A2(g13657), .A3(g13677), .A4(g13706) );
  AND2_X1 AND2_1683( .ZN(g18997), .A1(g13541), .A2(g16278) );
  AND4_X1 AND4_45( .ZN(g19007), .A1(g14976), .A2(g13687), .A3(g13714), .A4(g13756) );
  AND2_X2 AND2_1684( .ZN(g19010), .A1(g13552), .A2(g16337) );
  AND4_X1 AND4_46( .ZN(g19063), .A1(g18679), .A2(g14910), .A3(g13687), .A4(g16254) );
  AND4_X1 AND4_47( .ZN(g19079), .A1(g14797), .A2(g18692), .A3(g16142), .A4(g16189) );
  AND4_X1 AND4_48( .ZN(g19080), .A1(g18708), .A2(g14991), .A3(g13724), .A4(g16313) );
  AND2_X1 AND2_1685( .ZN(g19087), .A1(g17215), .A2(g16540) );
  AND4_X1 AND4_49( .ZN(g19088), .A1(g18656), .A2(g14797), .A3(g16189), .A4(g13706) );
  AND4_X1 AND4_50( .ZN(g19089), .A1(g14849), .A2(g18728), .A3(g16201), .A4(g16254) );
  AND4_X1 AND4_51( .ZN(g19090), .A1(g18744), .A2(g15080), .A3(g13774), .A4(g16371) );
  AND4_X1 AND4_52( .ZN(g19092), .A1(g14776), .A2(g18670), .A3(g18692), .A4(g16293) );
  AND2_X1 AND2_1686( .ZN(g19093), .A1(g17218), .A2(g16572) );
  AND4_X1 AND4_53( .ZN(g19094), .A1(g18679), .A2(g14849), .A3(g16254), .A4(g13756) );
  AND4_X1 AND4_54( .ZN(g19095), .A1(g14922), .A2(g18765), .A3(g16266), .A4(g16313) );
  AND3_X1 AND3_30( .ZN(II25280), .A1(g18656), .A2(g18670), .A3(g18720) );
  AND3_X1 AND3_31( .ZN(g19097), .A1(g13657), .A2(g16243), .A3(II25280) );
  AND4_X1 AND4_55( .ZN(g19099), .A1(g14811), .A2(g18699), .A3(g18728), .A4(g16351) );
  AND2_X2 AND2_1687( .ZN(g19100), .A1(g17220), .A2(g16596) );
  AND4_X1 AND4_56( .ZN(g19101), .A1(g18708), .A2(g14922), .A3(g16313), .A4(g13797) );
  AND4_X1 AND4_57( .ZN(g19102), .A1(g15003), .A2(g18796), .A3(g16325), .A4(g16371) );
  AND3_X1 AND3_32( .ZN(II25291), .A1(g18679), .A2(g18699), .A3(g18758) );
  AND3_X1 AND3_33( .ZN(g19104), .A1(g13687), .A2(g16302), .A3(II25291) );
  AND4_X1 AND4_58( .ZN(g19106), .A1(g14863), .A2(g18735), .A3(g18765), .A4(g16395) );
  AND2_X2 AND2_1688( .ZN(g19107), .A1(g17223), .A2(g16616) );
  AND4_X1 AND4_59( .ZN(g19108), .A1(g18744), .A2(g15003), .A3(g16371), .A4(g13825) );
  AND3_X1 AND3_34( .ZN(II25300), .A1(g18708), .A2(g18735), .A3(g18789) );
  AND3_X4 AND3_35( .ZN(g19109), .A1(g13724), .A2(g16360), .A3(II25300) );
  AND4_X1 AND4_60( .ZN(g19111), .A1(g14936), .A2(g18772), .A3(g18796), .A4(g16433) );
  AND2_X1 AND2_1689( .ZN(g19112), .A1(g14657), .A2(g16633) );
  AND3_X1 AND3_36( .ZN(II25311), .A1(g18744), .A2(g18772), .A3(g18815) );
  AND3_X1 AND3_37( .ZN(g19116), .A1(g13774), .A2(g16404), .A3(II25311) );
  AND2_X1 AND2_1690( .ZN(g19117), .A1(g14691), .A2(g16644) );
  AND2_X1 AND2_1691( .ZN(g19124), .A1(g14725), .A2(g16656) );
  AND2_X1 AND2_1692( .ZN(g19131), .A1(g14753), .A2(g16673) );
  AND2_X1 AND2_1693( .ZN(g19142), .A1(g17159), .A2(g16719) );
  AND2_X1 AND2_1694( .ZN(g19143), .A1(g17174), .A2(g16761) );
  AND2_X1 AND2_1695( .ZN(g19146), .A1(g17191), .A2(g16788) );
  AND2_X1 AND2_1696( .ZN(g19148), .A1(g17202), .A2(g16817) );
  AND2_X1 AND2_1697( .ZN(g19150), .A1(g17189), .A2(g8602) );
  AND2_X1 AND2_1698( .ZN(g19155), .A1(g17200), .A2(g8614) );
  AND2_X1 AND2_1699( .ZN(g19161), .A1(g17207), .A2(g8627) );
  AND2_X1 AND2_1700( .ZN(g19166), .A1(g17212), .A2(g8637) );
  AND2_X1 AND2_1701( .ZN(g19228), .A1(g16662), .A2(g12125) );
  AND2_X1 AND2_1702( .ZN(g19236), .A1(g16935), .A2(g8802) );
  AND3_X1 AND3_38( .ZN(g19241), .A1(g16867), .A2(g14158), .A3(g14071) );
  AND2_X1 AND2_1703( .ZN(g19248), .A1(g16662), .A2(g8817) );
  AND2_X1 AND2_1704( .ZN(g19252), .A1(g18725), .A2(g9527) );
  AND3_X1 AND3_39( .ZN(g19254), .A1(g16895), .A2(g14273), .A3(g14186) );
  AND2_X1 AND2_1705( .ZN(g19260), .A1(g16749), .A2(g3124) );
  AND3_X1 AND3_40( .ZN(g19267), .A1(g16924), .A2(g14395), .A3(g14301) );
  AND3_X1 AND3_41( .ZN(g19282), .A1(g16954), .A2(g14507), .A3(g14423) );
  AND2_X1 AND2_1706( .ZN(g19284), .A1(g18063), .A2(g3111) );
  AND2_X1 AND2_1707( .ZN(g19285), .A1(g16749), .A2(g7642) );
  AND2_X1 AND2_1708( .ZN(g19289), .A1(g17029), .A2(g8580) );
  AND3_X1 AND3_42( .ZN(g19303), .A1(g16867), .A2(g16543), .A3(g14071) );
  AND2_X1 AND2_1709( .ZN(g19307), .A1(g17063), .A2(g8587) );
  AND2_X1 AND2_1710( .ZN(g19316), .A1(g18063), .A2(g3110) );
  AND2_X1 AND2_1711( .ZN(g19317), .A1(g16749), .A2(g3126) );
  AND3_X1 AND3_43( .ZN(g19320), .A1(g16867), .A2(g16515), .A3(g14158) );
  AND3_X1 AND3_44( .ZN(g19324), .A1(g16895), .A2(g16575), .A3(g14186) );
  AND2_X1 AND2_1712( .ZN(g19328), .A1(g17098), .A2(g8594) );
  AND3_X1 AND3_45( .ZN(g19347), .A1(g16895), .A2(g16546), .A3(g14273) );
  AND3_X1 AND3_46( .ZN(g19351), .A1(g16924), .A2(g16599), .A3(g14301) );
  AND2_X1 AND2_1713( .ZN(g19355), .A1(g17136), .A2(g8605) );
  AND2_X1 AND2_1714( .ZN(g19356), .A1(g18063), .A2(g3112) );
  AND3_X1 AND3_47( .ZN(g19381), .A1(g16924), .A2(g16578), .A3(g14395) );
  AND3_X1 AND3_48( .ZN(g19385), .A1(g16954), .A2(g16619), .A3(g14423) );
  AND3_X1 AND3_49( .ZN(g19413), .A1(g16954), .A2(g16602), .A3(g14507) );
  AND3_X1 AND3_50( .ZN(g19449), .A1(g16884), .A2(g14797), .A3(g14776) );
  AND3_X1 AND3_51( .ZN(g19476), .A1(g16913), .A2(g14849), .A3(g14811) );
  AND3_X1 AND3_52( .ZN(g19499), .A1(g16943), .A2(g14922), .A3(g14863) );
  AND3_X1 AND3_53( .ZN(g19520), .A1(g16974), .A2(g15003), .A3(g14936) );
  AND3_X1 AND3_54( .ZN(g19531), .A1(g16884), .A2(g16722), .A3(g14776) );
  AND3_X1 AND3_55( .ZN(g19540), .A1(g16884), .A2(g16697), .A3(g14797) );
  AND3_X1 AND3_56( .ZN(g19541), .A1(g16913), .A2(g16764), .A3(g14811) );
  AND3_X1 AND3_57( .ZN(g19544), .A1(g16913), .A2(g16728), .A3(g14849) );
  AND3_X1 AND3_58( .ZN(g19545), .A1(g16943), .A2(g16791), .A3(g14863) );
  AND3_X1 AND3_59( .ZN(g19547), .A1(g16943), .A2(g16770), .A3(g14922) );
  AND3_X1 AND3_60( .ZN(g19548), .A1(g16974), .A2(g16820), .A3(g14936) );
  AND2_X1 AND2_1715( .ZN(g19549), .A1(g7950), .A2(g17230) );
  AND3_X1 AND3_61( .ZN(g19551), .A1(g16974), .A2(g16797), .A3(g15003) );
  AND2_X1 AND2_1716( .ZN(g19552), .A1(g16829), .A2(g6048) );
  AND2_X1 AND2_1717( .ZN(g19553), .A1(g7990), .A2(g17237) );
  AND2_X1 AND2_1718( .ZN(g19554), .A1(g7993), .A2(g17240) );
  AND2_X1 AND2_1719( .ZN(g19555), .A1(g8001), .A2(g17243) );
  AND2_X1 AND2_1720( .ZN(g19557), .A1(g8053), .A2(g17249) );
  AND2_X1 AND2_1721( .ZN(g19558), .A1(g8056), .A2(g17252) );
  AND2_X1 AND2_1722( .ZN(g19559), .A1(g8059), .A2(g17255) );
  AND2_X1 AND2_1723( .ZN(g19560), .A1(g8065), .A2(g17259) );
  AND2_X1 AND2_1724( .ZN(g19561), .A1(g8068), .A2(g17262) );
  AND2_X2 AND2_1725( .ZN(g19562), .A1(g8076), .A2(g17265) );
  AND2_X2 AND2_1726( .ZN(g19564), .A1(g8123), .A2(g17272) );
  AND2_X2 AND2_1727( .ZN(g19565), .A1(g8126), .A2(g17275) );
  AND2_X1 AND2_1728( .ZN(g19566), .A1(g8129), .A2(g17278) );
  AND2_X1 AND2_1729( .ZN(g19567), .A1(g8138), .A2(g17282) );
  AND2_X1 AND2_1730( .ZN(g19568), .A1(g8141), .A2(g17285) );
  AND2_X1 AND2_1731( .ZN(g19569), .A1(g8144), .A2(g17288) );
  AND2_X1 AND2_1732( .ZN(g19570), .A1(g8150), .A2(g17291) );
  AND2_X1 AND2_1733( .ZN(g19571), .A1(g8153), .A2(g17294) );
  AND2_X1 AND2_1734( .ZN(g19572), .A1(g8161), .A2(g17297) );
  AND2_X1 AND2_1735( .ZN(g19574), .A1(g8191), .A2(g17304) );
  AND2_X1 AND2_1736( .ZN(g19575), .A1(g8194), .A2(g17307) );
  AND2_X1 AND2_1737( .ZN(g19576), .A1(g8197), .A2(g17310) );
  AND2_X1 AND2_1738( .ZN(g19584), .A1(g640), .A2(g18756) );
  AND2_X1 AND2_1739( .ZN(g19585), .A1(g692), .A2(g18757) );
  AND2_X1 AND2_1740( .ZN(g19586), .A1(g8209), .A2(g17315) );
  AND2_X1 AND2_1741( .ZN(g19587), .A1(g8212), .A2(g17318) );
  AND2_X1 AND2_1742( .ZN(g19588), .A1(g8215), .A2(g17321) );
  AND2_X1 AND2_1743( .ZN(g19589), .A1(g8224), .A2(g17324) );
  AND2_X1 AND2_1744( .ZN(g19590), .A1(g8227), .A2(g17327) );
  AND2_X1 AND2_1745( .ZN(g19591), .A1(g8230), .A2(g17330) );
  AND2_X1 AND2_1746( .ZN(g19592), .A1(g8236), .A2(g17333) );
  AND2_X1 AND2_1747( .ZN(g19593), .A1(g8239), .A2(g17336) );
  AND2_X1 AND2_1748( .ZN(g19594), .A1(g16935), .A2(g12555) );
  AND2_X1 AND2_1749( .ZN(g19597), .A1(g3922), .A2(g17342) );
  AND2_X1 AND2_1750( .ZN(g19598), .A1(g3925), .A2(g17345) );
  AND2_X1 AND2_1751( .ZN(g19599), .A1(g3928), .A2(g17348) );
  AND2_X1 AND2_1752( .ZN(g19600), .A1(g633), .A2(g18783) );
  AND2_X1 AND2_1753( .ZN(g19601), .A1(g640), .A2(g18784) );
  AND2_X1 AND2_1754( .ZN(g19602), .A1(g633), .A2(g18785) );
  AND2_X1 AND2_1755( .ZN(g19603), .A1(g692), .A2(g18786) );
  AND2_X1 AND2_1756( .ZN(g19604), .A1(g3948), .A2(g17354) );
  AND2_X1 AND2_1757( .ZN(g19605), .A1(g3951), .A2(g17357) );
  AND2_X1 AND2_1758( .ZN(g19606), .A1(g3954), .A2(g17360) );
  AND2_X1 AND2_1759( .ZN(g19614), .A1(g1326), .A2(g18787) );
  AND2_X1 AND2_1760( .ZN(g19615), .A1(g1378), .A2(g18788) );
  AND2_X1 AND2_1761( .ZN(g19616), .A1(g3966), .A2(g17363) );
  AND2_X1 AND2_1762( .ZN(g19617), .A1(g3969), .A2(g17366) );
  AND2_X1 AND2_1763( .ZN(g19618), .A1(g3972), .A2(g17369) );
  AND2_X1 AND2_1764( .ZN(g19619), .A1(g3981), .A2(g17372) );
  AND2_X1 AND2_1765( .ZN(g19620), .A1(g3984), .A2(g17375) );
  AND2_X1 AND2_1766( .ZN(g19621), .A1(g3987), .A2(g17378) );
  AND2_X1 AND2_1767( .ZN(g19623), .A1(g4000), .A2(g17384) );
  AND2_X1 AND2_1768( .ZN(g19624), .A1(g4003), .A2(g17387) );
  AND2_X1 AND2_1769( .ZN(g19625), .A1(g4006), .A2(g17390) );
  AND2_X1 AND2_1770( .ZN(g19626), .A1(g640), .A2(g18805) );
  AND2_X1 AND2_1771( .ZN(g19627), .A1(g633), .A2(g18806) );
  AND2_X1 AND2_1772( .ZN(g19628), .A1(g653), .A2(g18807) );
  AND2_X1 AND2_1773( .ZN(g19629), .A1(g692), .A2(g18808) );
  AND2_X1 AND2_1774( .ZN(g19630), .A1(g4029), .A2(g17399) );
  AND2_X1 AND2_1775( .ZN(g19631), .A1(g4032), .A2(g17402) );
  AND2_X1 AND2_1776( .ZN(g19632), .A1(g4035), .A2(g17405) );
  AND2_X1 AND2_1777( .ZN(g19633), .A1(g1319), .A2(g18809) );
  AND2_X1 AND2_1778( .ZN(g19634), .A1(g1326), .A2(g18810) );
  AND2_X1 AND2_1779( .ZN(g19635), .A1(g1319), .A2(g18811) );
  AND2_X1 AND2_1780( .ZN(g19636), .A1(g1378), .A2(g18812) );
  AND2_X1 AND2_1781( .ZN(g19637), .A1(g4055), .A2(g17410) );
  AND2_X1 AND2_1782( .ZN(g19638), .A1(g4058), .A2(g17413) );
  AND2_X1 AND2_1783( .ZN(g19639), .A1(g4061), .A2(g17416) );
  AND2_X1 AND2_1784( .ZN(g19647), .A1(g2020), .A2(g18813) );
  AND2_X1 AND2_1785( .ZN(g19648), .A1(g2072), .A2(g18814) );
  AND2_X1 AND2_1786( .ZN(g19649), .A1(g4073), .A2(g17419) );
  AND2_X1 AND2_1787( .ZN(g19650), .A1(g4076), .A2(g17422) );
  AND2_X1 AND2_1788( .ZN(g19651), .A1(g4079), .A2(g17425) );
  AND2_X1 AND2_1789( .ZN(g19653), .A1(g4095), .A2(g17430) );
  AND2_X1 AND2_1790( .ZN(g19654), .A1(g4098), .A2(g17433) );
  AND2_X1 AND2_1791( .ZN(g19655), .A1(g4101), .A2(g17436) );
  AND2_X1 AND2_1792( .ZN(g19656), .A1(g4104), .A2(g17439) );
  AND2_X1 AND2_1793( .ZN(g19660), .A1(g633), .A2(g18822) );
  AND2_X1 AND2_1794( .ZN(g19661), .A1(g653), .A2(g18823) );
  AND2_X1 AND2_1795( .ZN(g19662), .A1(g646), .A2(g18824) );
  AND2_X1 AND2_1796( .ZN(g19663), .A1(g4127), .A2(g17451) );
  AND2_X2 AND2_1797( .ZN(g19664), .A1(g4130), .A2(g17454) );
  AND2_X2 AND2_1798( .ZN(g19665), .A1(g4133), .A2(g17457) );
  AND2_X2 AND2_1799( .ZN(g19666), .A1(g1326), .A2(g18825) );
  AND2_X1 AND2_1800( .ZN(g19667), .A1(g1319), .A2(g18826) );
  AND2_X1 AND2_1801( .ZN(g19668), .A1(g1339), .A2(g18827) );
  AND2_X1 AND2_1802( .ZN(g19669), .A1(g1378), .A2(g18828) );
  AND2_X1 AND2_1803( .ZN(g19670), .A1(g4156), .A2(g17465) );
  AND2_X1 AND2_1804( .ZN(g19671), .A1(g4159), .A2(g17468) );
  AND2_X1 AND2_1805( .ZN(g19672), .A1(g4162), .A2(g17471) );
  AND2_X1 AND2_1806( .ZN(g19673), .A1(g2013), .A2(g18829) );
  AND2_X1 AND2_1807( .ZN(g19674), .A1(g2020), .A2(g18830) );
  AND2_X1 AND2_1808( .ZN(g19675), .A1(g2013), .A2(g18831) );
  AND2_X1 AND2_1809( .ZN(g19676), .A1(g2072), .A2(g18832) );
  AND2_X1 AND2_1810( .ZN(g19677), .A1(g4182), .A2(g17476) );
  AND2_X1 AND2_1811( .ZN(g19678), .A1(g4185), .A2(g17479) );
  AND2_X1 AND2_1812( .ZN(g19679), .A1(g4188), .A2(g17482) );
  AND2_X1 AND2_1813( .ZN(g19687), .A1(g2714), .A2(g18833) );
  AND2_X1 AND2_1814( .ZN(g19688), .A1(g2766), .A2(g18834) );
  AND2_X1 AND2_1815( .ZN(g19691), .A1(g16841), .A2(g10865) );
  AND2_X1 AND2_1816( .ZN(g19692), .A1(g4205), .A2(g17487) );
  AND2_X1 AND2_1817( .ZN(g19693), .A1(g4208), .A2(g17490) );
  AND2_X1 AND2_1818( .ZN(g19694), .A1(g4211), .A2(g17493) );
  AND2_X1 AND2_1819( .ZN(g19695), .A1(g4214), .A2(g17496) );
  AND2_X1 AND2_1820( .ZN(g19697), .A1(g653), .A2(g18838) );
  AND2_X1 AND2_1821( .ZN(g19698), .A1(g646), .A2(g18839) );
  AND2_X1 AND2_1822( .ZN(g19699), .A1(g660), .A2(g18840) );
  AND2_X1 AND2_1823( .ZN(g19700), .A1(g17815), .A2(g16024) );
  AND2_X1 AND2_1824( .ZN(g19701), .A1(g4234), .A2(g17511) );
  AND2_X1 AND2_1825( .ZN(g19702), .A1(g4237), .A2(g17514) );
  AND2_X1 AND2_1826( .ZN(g19703), .A1(g4240), .A2(g17517) );
  AND2_X1 AND2_1827( .ZN(g19704), .A1(g4243), .A2(g17520) );
  AND2_X1 AND2_1828( .ZN(g19708), .A1(g1319), .A2(g18841) );
  AND2_X1 AND2_1829( .ZN(g19709), .A1(g1339), .A2(g18842) );
  AND2_X1 AND2_1830( .ZN(g19710), .A1(g1332), .A2(g18843) );
  AND2_X1 AND2_1831( .ZN(g19711), .A1(g4266), .A2(g17531) );
  AND2_X1 AND2_1832( .ZN(g19712), .A1(g4269), .A2(g17534) );
  AND2_X1 AND2_1833( .ZN(g19713), .A1(g4272), .A2(g17537) );
  AND2_X1 AND2_1834( .ZN(g19714), .A1(g2020), .A2(g18844) );
  AND2_X1 AND2_1835( .ZN(g19715), .A1(g2013), .A2(g18845) );
  AND2_X1 AND2_1836( .ZN(g19716), .A1(g2033), .A2(g18846) );
  AND2_X1 AND2_1837( .ZN(g19717), .A1(g2072), .A2(g18847) );
  AND2_X1 AND2_1838( .ZN(g19718), .A1(g4295), .A2(g17545) );
  AND2_X1 AND2_1839( .ZN(g19719), .A1(g4298), .A2(g17548) );
  AND2_X1 AND2_1840( .ZN(g19720), .A1(g4301), .A2(g17551) );
  AND2_X1 AND2_1841( .ZN(g19721), .A1(g2707), .A2(g18848) );
  AND2_X1 AND2_1842( .ZN(g19722), .A1(g2714), .A2(g18849) );
  AND2_X1 AND2_1843( .ZN(g19723), .A1(g2707), .A2(g18850) );
  AND2_X1 AND2_1844( .ZN(g19724), .A1(g2766), .A2(g18851) );
  AND2_X1 AND2_1845( .ZN(g19726), .A1(g16847), .A2(g6131) );
  AND2_X1 AND2_1846( .ZN(g19727), .A1(g4329), .A2(g17557) );
  AND2_X1 AND2_1847( .ZN(g19728), .A1(g4332), .A2(g17560) );
  AND2_X1 AND2_1848( .ZN(g19729), .A1(g4335), .A2(g17563) );
  AND2_X1 AND2_1849( .ZN(g19730), .A1(g653), .A2(g17573) );
  AND2_X1 AND2_1850( .ZN(g19731), .A1(g646), .A2(g18853) );
  AND2_X1 AND2_1851( .ZN(g19732), .A1(g660), .A2(g18854) );
  AND2_X1 AND2_1852( .ZN(g19733), .A1(g672), .A2(g18855) );
  AND2_X1 AND2_1853( .ZN(g19734), .A1(g17815), .A2(g16034) );
  AND2_X1 AND2_1854( .ZN(g19735), .A1(g17903), .A2(g16035) );
  AND2_X1 AND2_1855( .ZN(g19736), .A1(g4360), .A2(g17579) );
  AND2_X1 AND2_1856( .ZN(g19737), .A1(g4363), .A2(g17582) );
  AND2_X1 AND2_1857( .ZN(g19738), .A1(g4366), .A2(g17585) );
  AND2_X1 AND2_1858( .ZN(g19739), .A1(g4369), .A2(g17588) );
  AND2_X1 AND2_1859( .ZN(g19741), .A1(g1339), .A2(g18856) );
  AND2_X1 AND2_1860( .ZN(g19742), .A1(g1332), .A2(g18857) );
  AND2_X1 AND2_1861( .ZN(g19743), .A1(g1346), .A2(g18858) );
  AND2_X1 AND2_1862( .ZN(g19744), .A1(g17927), .A2(g16040) );
  AND2_X1 AND2_1863( .ZN(g19745), .A1(g4389), .A2(g17601) );
  AND2_X1 AND2_1864( .ZN(g19746), .A1(g4392), .A2(g17604) );
  AND2_X1 AND2_1865( .ZN(g19747), .A1(g4395), .A2(g17607) );
  AND2_X1 AND2_1866( .ZN(g19748), .A1(g4398), .A2(g17610) );
  AND2_X1 AND2_1867( .ZN(g19752), .A1(g2013), .A2(g18859) );
  AND2_X1 AND2_1868( .ZN(g19753), .A1(g2033), .A2(g18860) );
  AND2_X1 AND2_1869( .ZN(g19754), .A1(g2026), .A2(g18861) );
  AND2_X1 AND2_1870( .ZN(g19755), .A1(g4421), .A2(g17621) );
  AND2_X1 AND2_1871( .ZN(g19756), .A1(g4424), .A2(g17624) );
  AND2_X1 AND2_1872( .ZN(g19757), .A1(g4427), .A2(g17627) );
  AND2_X1 AND2_1873( .ZN(g19758), .A1(g2714), .A2(g18862) );
  AND2_X1 AND2_1874( .ZN(g19759), .A1(g2707), .A2(g18863) );
  AND2_X1 AND2_1875( .ZN(g19760), .A1(g2727), .A2(g18864) );
  AND2_X1 AND2_1876( .ZN(g19761), .A1(g2766), .A2(g18865) );
  AND2_X1 AND2_1877( .ZN(g19764), .A1(g4453), .A2(g17637) );
  AND2_X1 AND2_1878( .ZN(g19765), .A1(g660), .A2(g18870) );
  AND2_X1 AND2_1879( .ZN(g19766), .A1(g672), .A2(g18871) );
  AND2_X1 AND2_1880( .ZN(g19767), .A1(g666), .A2(g18872) );
  AND2_X1 AND2_1881( .ZN(g19768), .A1(g17815), .A2(g16054) );
  AND2_X1 AND2_1882( .ZN(g19769), .A1(g17903), .A2(g16055) );
  AND2_X1 AND2_1883( .ZN(g19770), .A1(g4498), .A2(g17655) );
  AND2_X1 AND2_1884( .ZN(g19771), .A1(g4501), .A2(g17658) );
  AND2_X1 AND2_1885( .ZN(g19772), .A1(g4504), .A2(g17661) );
  AND2_X1 AND2_1886( .ZN(g19773), .A1(g1339), .A2(g17670) );
  AND2_X1 AND2_1887( .ZN(g19774), .A1(g1332), .A2(g18874) );
  AND2_X1 AND2_1888( .ZN(g19775), .A1(g1346), .A2(g18875) );
  AND2_X1 AND2_1889( .ZN(g19776), .A1(g1358), .A2(g18876) );
  AND2_X1 AND2_1890( .ZN(g19777), .A1(g17927), .A2(g16056) );
  AND2_X1 AND2_1891( .ZN(g19778), .A1(g18014), .A2(g16057) );
  AND2_X1 AND2_1892( .ZN(g19779), .A1(g4529), .A2(g17676) );
  AND2_X1 AND2_1893( .ZN(g19780), .A1(g4532), .A2(g17679) );
  AND2_X1 AND2_1894( .ZN(g19781), .A1(g4535), .A2(g17682) );
  AND2_X1 AND2_1895( .ZN(g19782), .A1(g4538), .A2(g17685) );
  AND2_X1 AND2_1896( .ZN(g19784), .A1(g2033), .A2(g18877) );
  AND2_X1 AND2_1897( .ZN(g19785), .A1(g2026), .A2(g18878) );
  AND2_X1 AND2_1898( .ZN(g19786), .A1(g2040), .A2(g18879) );
  AND2_X1 AND2_1899( .ZN(g19787), .A1(g18038), .A2(g16062) );
  AND2_X1 AND2_1900( .ZN(g19788), .A1(g4558), .A2(g17698) );
  AND2_X1 AND2_1901( .ZN(g19789), .A1(g4561), .A2(g17701) );
  AND2_X1 AND2_1902( .ZN(g19790), .A1(g4564), .A2(g17704) );
  AND2_X1 AND2_1903( .ZN(g19791), .A1(g4567), .A2(g17707) );
  AND2_X1 AND2_1904( .ZN(g19795), .A1(g2707), .A2(g18880) );
  AND2_X1 AND2_1905( .ZN(g19796), .A1(g2727), .A2(g18881) );
  AND2_X1 AND2_1906( .ZN(g19797), .A1(g2720), .A2(g18882) );
  AND3_X1 AND3_62( .ZN(II26240), .A1(g18174), .A2(g18341), .A3(g17974) );
  AND3_X1 AND3_63( .ZN(g19799), .A1(g17640), .A2(g18074), .A3(II26240) );
  AND2_X1 AND2_1907( .ZN(g19802), .A1(g672), .A2(g18891) );
  AND2_X1 AND2_1908( .ZN(g19803), .A1(g666), .A2(g18892) );
  AND2_X1 AND2_1909( .ZN(g19804), .A1(g679), .A2(g18893) );
  AND2_X1 AND2_1910( .ZN(g19805), .A1(g17903), .A2(g16088) );
  AND2_X2 AND2_1911( .ZN(g19806), .A1(g4629), .A2(g17738) );
  AND2_X2 AND2_1912( .ZN(g19807), .A1(g1346), .A2(g18896) );
  AND2_X2 AND2_1913( .ZN(g19808), .A1(g1358), .A2(g18897) );
  AND2_X1 AND2_1914( .ZN(g19809), .A1(g1352), .A2(g18898) );
  AND2_X1 AND2_1915( .ZN(g19810), .A1(g17927), .A2(g16090) );
  AND2_X1 AND2_1916( .ZN(g19811), .A1(g18014), .A2(g16091) );
  AND2_X1 AND2_1917( .ZN(g19812), .A1(g4674), .A2(g17755) );
  AND2_X1 AND2_1918( .ZN(g19813), .A1(g4677), .A2(g17758) );
  AND2_X1 AND2_1919( .ZN(g19814), .A1(g4680), .A2(g17761) );
  AND2_X1 AND2_1920( .ZN(g19815), .A1(g2033), .A2(g17770) );
  AND2_X1 AND2_1921( .ZN(g19816), .A1(g2026), .A2(g18900) );
  AND2_X1 AND2_1922( .ZN(g19817), .A1(g2040), .A2(g18901) );
  AND2_X1 AND2_1923( .ZN(g19818), .A1(g2052), .A2(g18902) );
  AND2_X1 AND2_1924( .ZN(g19819), .A1(g18038), .A2(g16092) );
  AND2_X1 AND2_1925( .ZN(g19820), .A1(g18131), .A2(g16093) );
  AND2_X1 AND2_1926( .ZN(g19821), .A1(g4705), .A2(g17776) );
  AND2_X1 AND2_1927( .ZN(g19822), .A1(g4708), .A2(g17779) );
  AND2_X1 AND2_1928( .ZN(g19823), .A1(g4711), .A2(g17782) );
  AND2_X1 AND2_1929( .ZN(g19824), .A1(g4714), .A2(g17785) );
  AND2_X1 AND2_1930( .ZN(g19826), .A1(g2727), .A2(g18903) );
  AND2_X1 AND2_1931( .ZN(g19827), .A1(g2720), .A2(g18904) );
  AND2_X1 AND2_1932( .ZN(g19828), .A1(g2734), .A2(g18905) );
  AND2_X1 AND2_1933( .ZN(g19829), .A1(g18155), .A2(g16098) );
  AND2_X1 AND2_1934( .ZN(g19836), .A1(g7143), .A2(g18908) );
  AND2_X1 AND2_1935( .ZN(g19837), .A1(g6901), .A2(g17799) );
  AND2_X1 AND2_1936( .ZN(g19839), .A1(g666), .A2(g18909) );
  AND2_X1 AND2_1937( .ZN(g19840), .A1(g679), .A2(g18910) );
  AND2_X1 AND2_1938( .ZN(g19841), .A1(g686), .A2(g18911) );
  AND3_X1 AND3_64( .ZN(II26282), .A1(g18188), .A2(g18089), .A3(g17991) );
  AND3_X1 AND3_65( .ZN(g19842), .A1(g14525), .A2(g13922), .A3(II26282) );
  AND3_X1 AND3_66( .ZN(II26285), .A1(g18281), .A2(g18436), .A3(g18091) );
  AND3_X1 AND3_67( .ZN(g19843), .A1(g17741), .A2(g18190), .A3(II26285) );
  AND2_X1 AND2_1939( .ZN(g19846), .A1(g1358), .A2(g18914) );
  AND2_X1 AND2_1940( .ZN(g19847), .A1(g1352), .A2(g18915) );
  AND2_X1 AND2_1941( .ZN(g19848), .A1(g1365), .A2(g18916) );
  AND2_X1 AND2_1942( .ZN(g19849), .A1(g18014), .A2(g16126) );
  AND2_X1 AND2_1943( .ZN(g19850), .A1(g4806), .A2(g17839) );
  AND2_X1 AND2_1944( .ZN(g19851), .A1(g2040), .A2(g18919) );
  AND2_X1 AND2_1945( .ZN(g19852), .A1(g2052), .A2(g18920) );
  AND2_X1 AND2_1946( .ZN(g19853), .A1(g2046), .A2(g18921) );
  AND2_X1 AND2_1947( .ZN(g19854), .A1(g18038), .A2(g16128) );
  AND2_X1 AND2_1948( .ZN(g19855), .A1(g18131), .A2(g16129) );
  AND2_X1 AND2_1949( .ZN(g19856), .A1(g4851), .A2(g17856) );
  AND2_X1 AND2_1950( .ZN(g19857), .A1(g4854), .A2(g17859) );
  AND2_X1 AND2_1951( .ZN(g19858), .A1(g4857), .A2(g17862) );
  AND2_X1 AND2_1952( .ZN(g19859), .A1(g2727), .A2(g17871) );
  AND2_X1 AND2_1953( .ZN(g19860), .A1(g2720), .A2(g18923) );
  AND2_X1 AND2_1954( .ZN(g19861), .A1(g2734), .A2(g18924) );
  AND2_X1 AND2_1955( .ZN(g19862), .A1(g2746), .A2(g18925) );
  AND2_X1 AND2_1956( .ZN(g19863), .A1(g18155), .A2(g16130) );
  AND2_X1 AND2_1957( .ZN(g19864), .A1(g18247), .A2(g16131) );
  AND3_X1 AND3_68( .ZN(g19868), .A1(g16498), .A2(g16867), .A3(g19001) );
  AND2_X1 AND2_1958( .ZN(g19869), .A1(g679), .A2(g18926) );
  AND2_X1 AND2_1959( .ZN(g19870), .A1(g686), .A2(g18927) );
  AND3_X1 AND3_69( .ZN(II26311), .A1(g18353), .A2(g13958), .A3(g14011) );
  AND3_X1 AND3_70( .ZN(g19871), .A1(g14086), .A2(g18275), .A3(II26311) );
  AND2_X1 AND2_1960( .ZN(g19872), .A1(g1352), .A2(g18928) );
  AND2_X1 AND2_1961( .ZN(g19873), .A1(g1365), .A2(g18929) );
  AND2_X1 AND2_1962( .ZN(g19874), .A1(g1372), .A2(g18930) );
  AND3_X1 AND3_71( .ZN(II26317), .A1(g18295), .A2(g18205), .A3(g18108) );
  AND3_X1 AND3_72( .ZN(g19875), .A1(g14580), .A2(g13978), .A3(II26317) );
  AND3_X1 AND3_73( .ZN(II26320), .A1(g18374), .A2(g18509), .A3(g18207) );
  AND3_X1 AND3_74( .ZN(g19876), .A1(g17842), .A2(g18297), .A3(II26320) );
  AND2_X2 AND2_1963( .ZN(g19879), .A1(g2052), .A2(g18933) );
  AND2_X2 AND2_1964( .ZN(g19880), .A1(g2046), .A2(g18934) );
  AND2_X2 AND2_1965( .ZN(g19881), .A1(g2059), .A2(g18935) );
  AND2_X2 AND2_1966( .ZN(g19882), .A1(g18131), .A2(g16177) );
  AND2_X1 AND2_1967( .ZN(g19883), .A1(g4982), .A2(g17951) );
  AND2_X1 AND2_1968( .ZN(g19884), .A1(g2734), .A2(g18938) );
  AND2_X1 AND2_1969( .ZN(g19885), .A1(g2746), .A2(g18939) );
  AND2_X1 AND2_1970( .ZN(g19886), .A1(g2740), .A2(g18940) );
  AND2_X1 AND2_1971( .ZN(g19887), .A1(g18155), .A2(g16179) );
  AND2_X1 AND2_1972( .ZN(g19888), .A1(g18247), .A2(g16180) );
  AND2_X1 AND2_1973( .ZN(g19889), .A1(g2912), .A2(g18943) );
  AND2_X1 AND2_1974( .ZN(g19895), .A1(g686), .A2(g18945) );
  AND3_X1 AND3_75( .ZN(g19899), .A1(g16520), .A2(g16895), .A3(g16507) );
  AND2_X1 AND2_1975( .ZN(g19900), .A1(g1365), .A2(g18946) );
  AND2_X1 AND2_1976( .ZN(g19901), .A1(g1372), .A2(g18947) );
  AND3_X1 AND3_76( .ZN(II26348), .A1(g18448), .A2(g14028), .A3(g14102) );
  AND3_X1 AND3_77( .ZN(g19902), .A1(g14201), .A2(g18368), .A3(II26348) );
  AND2_X1 AND2_1977( .ZN(g19903), .A1(g2046), .A2(g18948) );
  AND2_X1 AND2_1978( .ZN(g19904), .A1(g2059), .A2(g18949) );
  AND2_X1 AND2_1979( .ZN(g19905), .A1(g2066), .A2(g18950) );
  AND3_X1 AND3_78( .ZN(II26354), .A1(g18388), .A2(g18312), .A3(g18224) );
  AND3_X1 AND3_79( .ZN(g19906), .A1(g14614), .A2(g14048), .A3(II26354) );
  AND3_X1 AND3_80( .ZN(II26357), .A1(g18469), .A2(g18573), .A3(g18314) );
  AND3_X1 AND3_81( .ZN(g19907), .A1(g17954), .A2(g18390), .A3(II26357) );
  AND2_X1 AND2_1980( .ZN(g19910), .A1(g2746), .A2(g18953) );
  AND2_X1 AND2_1981( .ZN(g19911), .A1(g2740), .A2(g18954) );
  AND2_X1 AND2_1982( .ZN(g19912), .A1(g2753), .A2(g18955) );
  AND2_X1 AND2_1983( .ZN(g19913), .A1(g18247), .A2(g16236) );
  AND2_X1 AND2_1984( .ZN(g19914), .A1(g3018), .A2(g18958) );
  AND2_X1 AND2_1985( .ZN(g19920), .A1(g1372), .A2(g18961) );
  AND3_X1 AND3_82( .ZN(g19924), .A1(g16551), .A2(g16924), .A3(g16529) );
  AND2_X1 AND2_1986( .ZN(g19925), .A1(g2059), .A2(g18962) );
  AND2_X1 AND2_1987( .ZN(g19926), .A1(g2066), .A2(g18963) );
  AND3_X1 AND3_83( .ZN(II26377), .A1(g18521), .A2(g14119), .A3(g14217) );
  AND3_X1 AND3_84( .ZN(g19927), .A1(g14316), .A2(g18463), .A3(II26377) );
  AND2_X1 AND2_1988( .ZN(g19928), .A1(g2740), .A2(g18964) );
  AND2_X1 AND2_1989( .ZN(g19929), .A1(g2753), .A2(g18965) );
  AND2_X1 AND2_1990( .ZN(g19930), .A1(g2760), .A2(g18966) );
  AND3_X1 AND3_85( .ZN(II26383), .A1(g18483), .A2(g18405), .A3(g18331) );
  AND3_X1 AND3_86( .ZN(g19931), .A1(g14637), .A2(g14139), .A3(II26383) );
  AND2_X1 AND2_1991( .ZN(g19932), .A1(g2917), .A2(g18166) );
  AND2_X1 AND2_1992( .ZN(g19935), .A1(g2066), .A2(g18972) );
  AND3_X1 AND3_87( .ZN(g19939), .A1(g16583), .A2(g16954), .A3(g16560) );
  AND2_X1 AND2_1993( .ZN(g19940), .A1(g2753), .A2(g18973) );
  AND2_X1 AND2_1994( .ZN(g19941), .A1(g2760), .A2(g18974) );
  AND3_X1 AND3_88( .ZN(II26396), .A1(g18585), .A2(g14234), .A3(g14332) );
  AND3_X1 AND3_89( .ZN(g19942), .A1(g14438), .A2(g18536), .A3(II26396) );
  AND2_X1 AND2_1995( .ZN(g19943), .A1(g7562), .A2(g18976) );
  AND2_X1 AND2_1996( .ZN(g19944), .A1(g3028), .A2(g18258) );
  AND2_X1 AND2_1997( .ZN(g19949), .A1(g5293), .A2(g18278) );
  AND2_X1 AND2_1998( .ZN(g19952), .A1(g2760), .A2(g18987) );
  AND2_X1 AND2_1999( .ZN(g19953), .A1(g7566), .A2(g18334) );
  AND3_X1 AND3_90( .ZN(II26416), .A1(g18553), .A2(g18491), .A3(g18431) );
  AND3_X1 AND3_91( .ZN(g19970), .A1(g18354), .A2(g18276), .A3(II26416) );
  AND2_X1 AND2_2000( .ZN(g19971), .A1(g5327), .A2(g18355) );
  AND2_X1 AND2_2001( .ZN(g19976), .A1(g5330), .A2(g18371) );
  AND3_X1 AND3_92( .ZN(II26432), .A1(g18277), .A2(g18189), .A3(g18090) );
  AND3_X1 AND3_93( .ZN(g19982), .A1(g17992), .A2(g17913), .A3(II26432) );
  AND2_X1 AND2_2002( .ZN(g19983), .A1(g5352), .A2(g18432) );
  AND3_X1 AND3_94( .ZN(II26440), .A1(g18603), .A2(g18555), .A3(g18504) );
  AND3_X1 AND3_95( .ZN(g20000), .A1(g18449), .A2(g18369), .A3(II26440) );
  AND2_X1 AND2_2003( .ZN(g20001), .A1(g5355), .A2(g18450) );
  AND2_X1 AND2_2004( .ZN(g20006), .A1(g5358), .A2(g18466) );
  AND2_X1 AND2_2005( .ZN(g20011), .A1(g18063), .A2(g3113) );
  AND2_X1 AND2_2006( .ZN(g20012), .A1(g16804), .A2(g3135) );
  AND2_X1 AND2_2007( .ZN(g20013), .A1(g17720), .A2(g12848) );
  AND2_X1 AND2_2008( .ZN(g20014), .A1(g7615), .A2(g16749) );
  AND3_X1 AND3_96( .ZN(II26464), .A1(g18370), .A2(g18296), .A3(g18206) );
  AND3_X1 AND3_97( .ZN(g20020), .A1(g18109), .A2(g18024), .A3(II26464) );
  AND2_X1 AND2_2009( .ZN(g20021), .A1(g5369), .A2(g18505) );
  AND3_X1 AND3_98( .ZN(II26472), .A1(g18635), .A2(g18605), .A3(g18568) );
  AND3_X1 AND3_99( .ZN(g20038), .A1(g18522), .A2(g18464), .A3(II26472) );
  AND2_X1 AND2_2010( .ZN(g20039), .A1(g5372), .A2(g18523) );
  AND2_X1 AND2_2011( .ZN(g20044), .A1(g5375), .A2(g18539) );
  AND2_X1 AND2_2012( .ZN(g20048), .A1(g16749), .A2(g3127) );
  AND2_X1 AND2_2013( .ZN(g20049), .A1(g17878), .A2(g3155) );
  AND2_X1 AND2_2014( .ZN(g20050), .A1(g18070), .A2(g3161) );
  AND2_X1 AND2_2015( .ZN(g20051), .A1(g18063), .A2(g3114) );
  AND2_X1 AND2_2016( .ZN(g20052), .A1(g16804), .A2(g3134) );
  AND2_X1 AND2_2017( .ZN(g20053), .A1(g17720), .A2(g12875) );
  AND3_X1 AND3_100( .ZN(II26500), .A1(g18465), .A2(g18389), .A3(g18313) );
  AND3_X1 AND3_101( .ZN(g20062), .A1(g18225), .A2(g18141), .A3(II26500) );
  AND2_X1 AND2_2018( .ZN(g20063), .A1(g5382), .A2(g18569) );
  AND3_X1 AND3_102( .ZN(II26508), .A1(g18644), .A2(g18637), .A3(g18618) );
  AND3_X1 AND3_103( .ZN(g20080), .A1(g18586), .A2(g18537), .A3(II26508) );
  AND2_X1 AND2_2019( .ZN(g20081), .A1(g5385), .A2(g18587) );
  AND2_X1 AND2_2020( .ZN(g20084), .A1(g17969), .A2(g3158) );
  AND2_X1 AND2_2021( .ZN(g20085), .A1(g18170), .A2(g3164) );
  AND2_X1 AND2_2022( .ZN(g20086), .A1(g18337), .A2(g3170) );
  AND2_X1 AND2_2023( .ZN(g20087), .A1(g16749), .A2(g7574) );
  AND2_X1 AND2_2024( .ZN(g20088), .A1(g16836), .A2(g3147) );
  AND2_X1 AND2_2025( .ZN(g20089), .A1(g17969), .A2(g9160) );
  AND2_X1 AND2_2026( .ZN(g20090), .A1(g18063), .A2(g3120) );
  AND2_X1 AND2_2027( .ZN(g20091), .A1(g16804), .A2(g3136) );
  AND2_X1 AND2_2028( .ZN(g20092), .A1(g16749), .A2(g7603) );
  AND3_X1 AND3_104( .ZN(II26525), .A1(g18656), .A2(g18670), .A3(g18692) );
  AND4_X1 AND4_61( .ZN(g20093), .A1(g13657), .A2(g13677), .A3(g13750), .A4(II26525) );
  AND3_X1 AND3_105( .ZN(II26528), .A1(g18656), .A2(g14837), .A3(g13657) );
  AND3_X1 AND3_106( .ZN(g20094), .A1(g13677), .A2(g13706), .A3(II26528) );
  AND3_X1 AND3_107( .ZN(II26541), .A1(g18538), .A2(g18484), .A3(g18406) );
  AND3_X1 AND3_108( .ZN(g20103), .A1(g18332), .A2(g18257), .A3(II26541) );
  AND2_X1 AND2_2029( .ZN(g20104), .A1(g5391), .A2(g18619) );
  AND2_X1 AND2_2030( .ZN(g20106), .A1(g18261), .A2(g3167) );
  AND2_X1 AND2_2031( .ZN(g20107), .A1(g18415), .A2(g3173) );
  AND2_X1 AND2_2032( .ZN(g20108), .A1(g18543), .A2(g3179) );
  AND2_X1 AND2_2033( .ZN(g20109), .A1(g17878), .A2(g9504) );
  AND2_X1 AND2_2034( .ZN(g20110), .A1(g18070), .A2(g9286) );
  AND2_X1 AND2_2035( .ZN(g20111), .A1(g18261), .A2(g9884) );
  AND2_X1 AND2_2036( .ZN(g20112), .A1(g16749), .A2(g3132) );
  AND2_X1 AND2_2037( .ZN(g20113), .A1(g16836), .A2(g3142) );
  AND2_X1 AND2_2038( .ZN(g20114), .A1(g17969), .A2(g9755) );
  AND2_X1 AND2_2039( .ZN(g20115), .A1(g16804), .A2(g3139) );
  AND3_X1 AND3_109( .ZN(II26558), .A1(g14776), .A2(g18670), .A3(g18720) );
  AND4_X1 AND4_62( .ZN(g20116), .A1(g16142), .A2(g13677), .A3(g13706), .A4(II26558) );
  AND3_X1 AND3_110( .ZN(II26561), .A1(g14776), .A2(g18720), .A3(g13657) );
  AND3_X1 AND3_111( .ZN(g20117), .A1(g16189), .A2(g13706), .A3(II26561) );
  AND3_X1 AND3_112( .ZN(II26564), .A1(g18679), .A2(g18699), .A3(g18728) );
  AND4_X1 AND4_63( .ZN(g20118), .A1(g13687), .A2(g13714), .A3(g13791), .A4(II26564) );
  AND3_X1 AND3_113( .ZN(II26567), .A1(g18679), .A2(g14910), .A3(g13687) );
  AND3_X1 AND3_114( .ZN(g20119), .A1(g13714), .A2(g13756), .A3(II26567) );
  AND2_X1 AND2_2040( .ZN(g20131), .A1(g18486), .A2(g3176) );
  AND2_X1 AND2_2041( .ZN(g20132), .A1(g18593), .A2(g3182) );
  AND2_X1 AND2_2042( .ZN(g20133), .A1(g18170), .A2(g9505) );
  AND2_X1 AND2_2043( .ZN(g20134), .A1(g18337), .A2(g9506) );
  AND2_X1 AND2_2044( .ZN(g20135), .A1(g18486), .A2(g9885) );
  AND2_X1 AND2_2045( .ZN(g20136), .A1(g17878), .A2(g9423) );
  AND2_X1 AND2_2046( .ZN(g20137), .A1(g18070), .A2(g9226) );
  AND2_X1 AND2_2047( .ZN(g20138), .A1(g18261), .A2(g9756) );
  AND2_X1 AND2_2048( .ZN(g20139), .A1(g16836), .A2(g3151) );
  AND3_X1 AND3_115( .ZN(g20144), .A1(g16679), .A2(g16884), .A3(g16665) );
  AND4_X1 AND4_64( .ZN(g20145), .A1(g14776), .A2(g18670), .A3(g16142), .A4(g16189) );
  AND3_X1 AND3_116( .ZN(II26590), .A1(g14811), .A2(g18699), .A3(g18758) );
  AND4_X1 AND4_65( .ZN(g20146), .A1(g16201), .A2(g13714), .A3(g13756), .A4(II26590) );
  AND3_X1 AND3_117( .ZN(II26593), .A1(g14811), .A2(g18758), .A3(g13687) );
  AND3_X1 AND3_118( .ZN(g20147), .A1(g16254), .A2(g13756), .A3(II26593) );
  AND3_X1 AND3_119( .ZN(II26596), .A1(g18708), .A2(g18735), .A3(g18765) );
  AND4_X1 AND4_66( .ZN(g20148), .A1(g13724), .A2(g13764), .A3(g13819), .A4(II26596) );
  AND3_X1 AND3_120( .ZN(II26599), .A1(g18708), .A2(g14991), .A3(g13724) );
  AND3_X1 AND3_121( .ZN(g20149), .A1(g13764), .A2(g13797), .A3(II26599) );
  AND2_X1 AND2_2049( .ZN(g20156), .A1(g16809), .A2(g3185) );
  AND2_X1 AND2_2050( .ZN(g20157), .A1(g18415), .A2(g9287) );
  AND2_X1 AND2_2051( .ZN(g20158), .A1(g18543), .A2(g9886) );
  AND2_X1 AND2_2052( .ZN(g20159), .A1(g16809), .A2(g9288) );
  AND2_X1 AND2_2053( .ZN(g20160), .A1(g18170), .A2(g9424) );
  AND2_X1 AND2_2054( .ZN(g20161), .A1(g18337), .A2(g9426) );
  AND2_X1 AND2_2055( .ZN(g20162), .A1(g18486), .A2(g9757) );
  AND3_X1 AND3_122( .ZN(II26615), .A1(g14797), .A2(g18692), .A3(g13657) );
  AND3_X1 AND3_123( .ZN(g20177), .A1(g13677), .A2(g13750), .A3(II26615) );
  AND3_X1 AND3_124( .ZN(g20182), .A1(g16705), .A2(g16913), .A3(g16686) );
  AND4_X1 AND4_67( .ZN(g20183), .A1(g14811), .A2(g18699), .A3(g16201), .A4(g16254) );
  AND3_X1 AND3_125( .ZN(II26621), .A1(g14863), .A2(g18735), .A3(g18789) );
  AND4_X1 AND4_68( .ZN(g20184), .A1(g16266), .A2(g13764), .A3(g13797), .A4(II26621) );
  AND3_X1 AND3_126( .ZN(II26624), .A1(g14863), .A2(g18789), .A3(g13724) );
  AND3_X1 AND3_127( .ZN(g20185), .A1(g16313), .A2(g13797), .A3(II26624) );
  AND3_X1 AND3_128( .ZN(II26627), .A1(g18744), .A2(g18772), .A3(g18796) );
  AND4_X1 AND4_69( .ZN(g20186), .A1(g13774), .A2(g13805), .A3(g13840), .A4(II26627) );
  AND3_X1 AND3_129( .ZN(II26630), .A1(g18744), .A2(g15080), .A3(g13774) );
  AND3_X1 AND3_130( .ZN(g20187), .A1(g13805), .A2(g13825), .A3(II26630) );
  AND2_X1 AND2_2056( .ZN(g20188), .A1(g18593), .A2(g9425) );
  AND2_X1 AND2_2057( .ZN(g20189), .A1(g16825), .A2(g9289) );
  AND2_X1 AND2_2058( .ZN(g20190), .A1(g18415), .A2(g9227) );
  AND2_X1 AND2_2059( .ZN(g20191), .A1(g18543), .A2(g9758) );
  AND2_X1 AND2_2060( .ZN(g20192), .A1(g16809), .A2(g9228) );
  AND3_X1 AND3_131( .ZN(II26639), .A1(g18656), .A2(g18670), .A3(g16142) );
  AND3_X1 AND3_132( .ZN(g20197), .A1(g13677), .A2(g13706), .A3(II26639) );
  AND3_X1 AND3_133( .ZN(II26645), .A1(g14849), .A2(g18728), .A3(g13687) );
  AND3_X1 AND3_134( .ZN(g20211), .A1(g13714), .A2(g13791), .A3(II26645) );
  AND3_X1 AND3_135( .ZN(g20216), .A1(g16736), .A2(g16943), .A3(g16712) );
  AND4_X1 AND4_70( .ZN(g20217), .A1(g14863), .A2(g18735), .A3(g16266), .A4(g16313) );
  AND3_X1 AND3_136( .ZN(II26651), .A1(g14936), .A2(g18772), .A3(g18815) );
  AND4_X1 AND4_71( .ZN(g20218), .A1(g16325), .A2(g13805), .A3(g13825), .A4(II26651) );
  AND3_X1 AND3_137( .ZN(II26654), .A1(g14936), .A2(g18815), .A3(g13774) );
  AND3_X1 AND3_138( .ZN(g20219), .A1(g16371), .A2(g13825), .A3(II26654) );
  AND2_X1 AND2_2061( .ZN(g20220), .A1(g18593), .A2(g9355) );
  AND2_X1 AND2_2062( .ZN(g20221), .A1(g16825), .A2(g10099) );
  AND4_X1 AND4_72( .ZN(g20222), .A1(g18656), .A2(g18720), .A3(g13657), .A4(g16293) );
  AND3_X1 AND3_139( .ZN(II26661), .A1(g18679), .A2(g18699), .A3(g16201) );
  AND3_X1 AND3_140( .ZN(g20227), .A1(g13714), .A2(g13756), .A3(II26661) );
  AND3_X1 AND3_141( .ZN(II26667), .A1(g14922), .A2(g18765), .A3(g13724) );
  AND3_X1 AND3_142( .ZN(g20241), .A1(g13764), .A2(g13819), .A3(II26667) );
  AND3_X1 AND3_143( .ZN(g20246), .A1(g16778), .A2(g16974), .A3(g16743) );
  AND4_X1 AND4_73( .ZN(g20247), .A1(g14936), .A2(g18772), .A3(g16325), .A4(g16371) );
  AND3_X1 AND3_144( .ZN(g20248), .A1(g18656), .A2(g14837), .A3(g16293) );
  AND4_X1 AND4_74( .ZN(g20249), .A1(g18679), .A2(g18758), .A3(g13687), .A4(g16351) );
  AND3_X1 AND3_145( .ZN(II26676), .A1(g18708), .A2(g18735), .A3(g16266) );
  AND3_X1 AND3_146( .ZN(g20254), .A1(g13764), .A2(g13797), .A3(II26676) );
  AND3_X1 AND3_147( .ZN(II26682), .A1(g15003), .A2(g18796), .A3(g13774) );
  AND3_X1 AND3_148( .ZN(g20268), .A1(g13805), .A2(g13840), .A3(II26682) );
  AND4_X1 AND4_75( .ZN(g20270), .A1(g14797), .A2(g18692), .A3(g13657), .A4(g16243) );
  AND3_X1 AND3_149( .ZN(g20271), .A1(g18679), .A2(g14910), .A3(g16351) );
  AND4_X1 AND4_76( .ZN(g20272), .A1(g18708), .A2(g18789), .A3(g13724), .A4(g16395) );
  AND3_X1 AND3_150( .ZN(II26690), .A1(g18744), .A2(g18772), .A3(g16325) );
  AND3_X1 AND3_151( .ZN(g20277), .A1(g13805), .A2(g13825), .A3(II26690) );
  AND3_X1 AND3_152( .ZN(II26695), .A1(g18670), .A2(g18692), .A3(g16142) );
  AND3_X1 AND3_153( .ZN(g20280), .A1(g13677), .A2(g16243), .A3(II26695) );
  AND4_X1 AND4_77( .ZN(g20282), .A1(g14849), .A2(g18728), .A3(g13687), .A4(g16302) );
  AND3_X1 AND3_154( .ZN(g20283), .A1(g18708), .A2(g14991), .A3(g16395) );
  AND4_X1 AND4_78( .ZN(g20284), .A1(g18744), .A2(g18815), .A3(g13774), .A4(g16433) );
  AND2_X1 AND2_2063( .ZN(g20285), .A1(g16846), .A2(g8103) );
  AND3_X1 AND3_155( .ZN(II26708), .A1(g18699), .A2(g18728), .A3(g16201) );
  AND3_X1 AND3_156( .ZN(g20291), .A1(g13714), .A2(g16302), .A3(II26708) );
  AND4_X1 AND4_79( .ZN(g20293), .A1(g14922), .A2(g18765), .A3(g13724), .A4(g16360) );
  AND3_X1 AND3_157( .ZN(g20294), .A1(g18744), .A2(g15080), .A3(g16433) );
  AND3_X1 AND3_158( .ZN(II26726), .A1(g18735), .A2(g18765), .A3(g16266) );
  AND3_X1 AND3_159( .ZN(g20307), .A1(g13764), .A2(g16360), .A3(II26726) );
  AND4_X1 AND4_80( .ZN(g20309), .A1(g15003), .A2(g18796), .A3(g13774), .A4(g16404) );
  AND3_X1 AND3_160( .ZN(II26745), .A1(g18772), .A2(g18796), .A3(g16325) );
  AND3_X1 AND3_161( .ZN(g20326), .A1(g13805), .A2(g16404), .A3(II26745) );
  AND2_X1 AND2_2064( .ZN(g20460), .A1(g17351), .A2(g13644) );
  AND2_X1 AND2_2065( .ZN(g20472), .A1(g17314), .A2(g13669) );
  AND2_X1 AND2_2066( .ZN(g20480), .A1(g17313), .A2(g11827) );
  AND2_X1 AND2_2067( .ZN(g20486), .A1(g17281), .A2(g11859) );
  AND2_X1 AND2_2068( .ZN(g20492), .A1(g17258), .A2(g11894) );
  AND2_X1 AND2_2069( .ZN(g20499), .A1(g17648), .A2(g11933) );
  AND2_X1 AND2_2070( .ZN(g20502), .A1(g17566), .A2(g11973) );
  AND2_X1 AND2_2071( .ZN(g20503), .A1(g17507), .A2(g13817) );
  AND2_X1 AND2_2072( .ZN(g20506), .A1(g17499), .A2(g12025) );
  AND2_X1 AND2_2073( .ZN(g20512), .A1(g17445), .A2(g13836) );
  AND2_X1 AND2_2074( .ZN(g20525), .A1(g17394), .A2(g13849) );
  AND4_X1 AND4_81( .ZN(g20538), .A1(g18656), .A2(g14837), .A3(g13657), .A4(g16189) );
  AND2_X1 AND2_2075( .ZN(g20640), .A1(g4809), .A2(g19064) );
  AND2_X1 AND2_2076( .ZN(g20647), .A1(g5888), .A2(g19075) );
  AND2_X1 AND2_2077( .ZN(g20665), .A1(g4985), .A2(g19081) );
  AND2_X1 AND2_2078( .ZN(g20809), .A1(g5712), .A2(g19113) );
  AND2_X1 AND2_2079( .ZN(g20826), .A1(g5770), .A2(g19118) );
  AND2_X1 AND2_2080( .ZN(g20836), .A1(g5829), .A2(g19125) );
  AND2_X1 AND2_2081( .ZN(g20840), .A1(g5885), .A2(g19132) );
  AND3_X1 AND3_162( .ZN(g21049), .A1(g20016), .A2(g14079), .A3(g14165) );
  AND2_X1 AND2_2082( .ZN(g21067), .A1(g20193), .A2(g12030) );
  AND3_X4 AND3_163( .ZN(g21068), .A1(g20058), .A2(g14194), .A3(g14280) );
  AND2_X1 AND2_2083( .ZN(g21077), .A1(g20223), .A2(g12094) );
  AND3_X2 AND3_164( .ZN(g21078), .A1(g20099), .A2(g14309), .A3(g14402) );
  AND3_X1 AND3_165( .ZN(g21085), .A1(g19484), .A2(g14158), .A3(g19001) );
  AND2_X1 AND2_2084( .ZN(g21086), .A1(g20193), .A2(g12142) );
  AND2_X1 AND2_2085( .ZN(g21091), .A1(g20250), .A2(g12166) );
  AND3_X1 AND3_166( .ZN(g21092), .A1(g20124), .A2(g14431), .A3(g14514) );
  AND3_X1 AND3_167( .ZN(g21097), .A1(g19505), .A2(g14273), .A3(g16507) );
  AND2_X1 AND2_2086( .ZN(g21098), .A1(g20223), .A2(g12204) );
  AND2_X1 AND2_2087( .ZN(g21103), .A1(g20273), .A2(g12228) );
  AND3_X1 AND3_168( .ZN(g21107), .A1(g19444), .A2(g17893), .A3(g14079) );
  AND3_X1 AND3_169( .ZN(g21111), .A1(g19524), .A2(g14395), .A3(g16529) );
  AND2_X2 AND2_2088( .ZN(g21112), .A1(g20250), .A2(g12259) );
  AND2_X2 AND2_2089( .ZN(g21121), .A1(g20054), .A2(g14244) );
  AND2_X1 AND2_2090( .ZN(g21122), .A1(g20140), .A2(g12279) );
  AND2_X1 AND2_2091( .ZN(g21123), .A1(g19970), .A2(g19982) );
  AND3_X1 AND3_170( .ZN(g21124), .A1(g19471), .A2(g18004), .A3(g14194) );
  AND3_X1 AND3_171( .ZN(g21128), .A1(g19534), .A2(g14507), .A3(g16560) );
  AND2_X1 AND2_2092( .ZN(g21129), .A1(g20273), .A2(g12302) );
  AND3_X1 AND3_172( .ZN(II27695), .A1(g19318), .A2(g19300), .A3(g19286) );
  AND3_X1 AND3_173( .ZN(g21136), .A1(g19271), .A2(g19261), .A3(II27695) );
  AND2_X1 AND2_2093( .ZN(g21137), .A1(g5750), .A2(g19272) );
  AND2_X1 AND2_2094( .ZN(g21138), .A1(g19484), .A2(g14347) );
  AND2_X1 AND2_2095( .ZN(g21140), .A1(g20095), .A2(g14366) );
  AND2_X1 AND2_2096( .ZN(g21141), .A1(g20178), .A2(g12315) );
  AND2_X1 AND2_2097( .ZN(g21142), .A1(g20000), .A2(g20020) );
  AND3_X1 AND3_174( .ZN(g21143), .A1(g19494), .A2(g18121), .A3(g14309) );
  AND3_X1 AND3_175( .ZN(II27711), .A1(g19262), .A2(g19414), .A3(g19386) );
  AND3_X1 AND3_176( .ZN(g21152), .A1(g19357), .A2(g19334), .A3(II27711) );
  AND3_X1 AND3_177( .ZN(g21153), .A1(g20054), .A2(g16543), .A3(g16501) );
  AND2_X1 AND2_2098( .ZN(g21154), .A1(g20193), .A2(g12333) );
  AND2_X1 AND2_2099( .ZN(g21155), .A1(g20140), .A2(g12336) );
  AND3_X1 AND3_178( .ZN(II27717), .A1(g19345), .A2(g19321), .A3(g19304) );
  AND3_X1 AND3_179( .ZN(g21156), .A1(g19290), .A2(g19276), .A3(II27717) );
  AND2_X1 AND2_2100( .ZN(g21157), .A1(g5809), .A2(g19291) );
  AND2_X1 AND2_2101( .ZN(g21158), .A1(g19505), .A2(g14459) );
  AND2_X1 AND2_2102( .ZN(g21160), .A1(g20120), .A2(g14478) );
  AND2_X1 AND2_2103( .ZN(g21161), .A1(g20212), .A2(g12343) );
  AND2_X1 AND2_2104( .ZN(g21162), .A1(g20038), .A2(g20062) );
  AND3_X1 AND3_180( .ZN(g21163), .A1(g19515), .A2(g18237), .A3(g14431) );
  AND3_X1 AND3_181( .ZN(II27733), .A1(g19277), .A2(g19451), .A3(g19416) );
  AND3_X1 AND3_182( .ZN(g21172), .A1(g19389), .A2(g19368), .A3(II27733) );
  AND3_X1 AND3_183( .ZN(g21173), .A1(g20095), .A2(g16575), .A3(g16523) );
  AND2_X1 AND2_2105( .ZN(g21174), .A1(g20223), .A2(g12363) );
  AND2_X1 AND2_2106( .ZN(g21175), .A1(g20178), .A2(g12366) );
  AND3_X1 AND3_184( .ZN(II27739), .A1(g19379), .A2(g19348), .A3(g19325) );
  AND3_X1 AND3_185( .ZN(g21176), .A1(g19308), .A2(g19295), .A3(II27739) );
  AND2_X1 AND2_2107( .ZN(g21177), .A1(g5865), .A2(g19309) );
  AND2_X1 AND2_2108( .ZN(g21178), .A1(g19524), .A2(g14546) );
  AND2_X1 AND2_2109( .ZN(g21180), .A1(g20150), .A2(g14565) );
  AND2_X1 AND2_2110( .ZN(g21181), .A1(g20242), .A2(g12373) );
  AND2_X1 AND2_2111( .ZN(g21182), .A1(g20080), .A2(g20103) );
  AND2_X1 AND2_2112( .ZN(g21188), .A1(g20140), .A2(g12379) );
  AND3_X1 AND3_186( .ZN(II27755), .A1(g19296), .A2(g19478), .A3(g19453) );
  AND3_X1 AND3_187( .ZN(g21192), .A1(g19419), .A2(g19400), .A3(II27755) );
  AND3_X1 AND3_188( .ZN(g21193), .A1(g20120), .A2(g16599), .A3(g16554) );
  AND2_X1 AND2_2113( .ZN(g21194), .A1(g20250), .A2(g12382) );
  AND2_X1 AND2_2114( .ZN(g21195), .A1(g20212), .A2(g12385) );
  AND3_X1 AND3_189( .ZN(II27761), .A1(g19411), .A2(g19382), .A3(g19352) );
  AND3_X1 AND3_190( .ZN(g21196), .A1(g19329), .A2(g19313), .A3(II27761) );
  AND2_X1 AND2_2115( .ZN(g21197), .A1(g5912), .A2(g19330) );
  AND2_X1 AND2_2116( .ZN(g21198), .A1(g19534), .A2(g14601) );
  AND2_X1 AND2_2117( .ZN(g21203), .A1(g20178), .A2(g12409) );
  AND3_X1 AND3_191( .ZN(II27772), .A1(g19314), .A2(g19501), .A3(g19480) );
  AND3_X1 AND3_192( .ZN(g21207), .A1(g19456), .A2(g19430), .A3(II27772) );
  AND3_X1 AND3_193( .ZN(g21208), .A1(g20150), .A2(g16619), .A3(g16586) );
  AND2_X1 AND2_2118( .ZN(g21209), .A1(g20273), .A2(g12412) );
  AND2_X1 AND2_2119( .ZN(g21210), .A1(g20242), .A2(g12415) );
  AND2_X1 AND2_2120( .ZN(g21218), .A1(g20212), .A2(g12421) );
  AND2_X1 AND2_2121( .ZN(g21226), .A1(g20242), .A2(g12426) );
  AND3_X1 AND3_194( .ZN(g21229), .A1(g19578), .A2(g14797), .A3(g16665) );
  AND3_X1 AND3_195( .ZN(g21234), .A1(g19608), .A2(g14849), .A3(g16686) );
  AND3_X1 AND3_196( .ZN(g21243), .A1(g19641), .A2(g14922), .A3(g16712) );
  AND2_X1 AND2_2122( .ZN(g21245), .A1(g20299), .A2(g14837) );
  AND3_X1 AND3_197( .ZN(g21251), .A1(g19681), .A2(g15003), .A3(g16743) );
  AND2_X1 AND2_2123( .ZN(g21252), .A1(g19578), .A2(g14895) );
  AND2_X1 AND2_2124( .ZN(g21254), .A1(g20318), .A2(g14910) );
  AND3_X1 AND3_198( .ZN(g21259), .A1(g20299), .A2(g16722), .A3(g16682) );
  AND2_X1 AND2_2125( .ZN(g21260), .A1(g19608), .A2(g14976) );
  AND2_X1 AND2_2126( .ZN(g21262), .A1(g20337), .A2(g14991) );
  AND3_X1 AND3_199( .ZN(g21267), .A1(g20318), .A2(g16764), .A3(g16708) );
  AND2_X1 AND2_2127( .ZN(g21268), .A1(g19641), .A2(g15065) );
  AND2_X1 AND2_2128( .ZN(g21270), .A1(g20357), .A2(g15080) );
  AND3_X1 AND3_200( .ZN(g21276), .A1(g20337), .A2(g16791), .A3(g16739) );
  AND2_X1 AND2_2129( .ZN(g21277), .A1(g19681), .A2(g15161) );
  AND3_X1 AND3_201( .ZN(g21283), .A1(g20357), .A2(g16820), .A3(g16781) );
  AND2_X1 AND2_2130( .ZN(g21284), .A1(g9356), .A2(g20269) );
  AND2_X1 AND2_2131( .ZN(g21290), .A1(g9356), .A2(g20278) );
  AND2_X1 AND2_2132( .ZN(g21291), .A1(g9293), .A2(g20279) );
  AND2_X1 AND2_2133( .ZN(g21292), .A1(g9453), .A2(g20281) );
  AND2_X1 AND2_2134( .ZN(g21298), .A1(g9356), .A2(g20286) );
  AND2_X1 AND2_2135( .ZN(g21299), .A1(g9293), .A2(g20287) );
  AND2_X1 AND2_2136( .ZN(g21300), .A1(g9232), .A2(g20288) );
  AND2_X1 AND2_2137( .ZN(g21301), .A1(g9453), .A2(g20289) );
  AND2_X1 AND2_2138( .ZN(g21302), .A1(g9374), .A2(g20290) );
  AND2_X1 AND2_2139( .ZN(g21303), .A1(g9595), .A2(g20292) );
  AND2_X1 AND2_2140( .ZN(g21304), .A1(g9293), .A2(g20296) );
  AND2_X1 AND2_2141( .ZN(g21305), .A1(g9232), .A2(g20297) );
  AND2_X2 AND2_2142( .ZN(g21306), .A1(g9187), .A2(g20298) );
  AND2_X2 AND2_2143( .ZN(g21307), .A1(g9453), .A2(g20302) );
  AND2_X2 AND2_2144( .ZN(g21308), .A1(g9374), .A2(g20303) );
  AND2_X2 AND2_2145( .ZN(g21309), .A1(g9310), .A2(g20304) );
  AND2_X1 AND2_2146( .ZN(g21310), .A1(g9595), .A2(g20305) );
  AND2_X1 AND2_2147( .ZN(g21311), .A1(g9471), .A2(g20306) );
  AND2_X1 AND2_2148( .ZN(g21312), .A1(g9737), .A2(g20308) );
  AND2_X1 AND2_2149( .ZN(g21313), .A1(g9232), .A2(g20311) );
  AND2_X1 AND2_2150( .ZN(g21314), .A1(g9187), .A2(g20312) );
  AND2_X1 AND2_2151( .ZN(g21315), .A1(g9161), .A2(g20313) );
  AND2_X1 AND2_2152( .ZN(g21319), .A1(g9374), .A2(g20315) );
  AND2_X1 AND2_2153( .ZN(g21320), .A1(g9310), .A2(g20316) );
  AND2_X1 AND2_2154( .ZN(g21321), .A1(g9248), .A2(g20317) );
  AND2_X1 AND2_2155( .ZN(g21322), .A1(g9595), .A2(g20321) );
  AND2_X1 AND2_2156( .ZN(g21323), .A1(g9471), .A2(g20322) );
  AND2_X1 AND2_2157( .ZN(g21324), .A1(g9391), .A2(g20323) );
  AND2_X1 AND2_2158( .ZN(g21325), .A1(g9737), .A2(g20324) );
  AND2_X1 AND2_2159( .ZN(g21326), .A1(g9613), .A2(g20325) );
  AND2_X1 AND2_2160( .ZN(g21328), .A1(g9187), .A2(g20327) );
  AND2_X1 AND2_2161( .ZN(g21329), .A1(g9161), .A2(g20328) );
  AND2_X1 AND2_2162( .ZN(g21330), .A1(g9150), .A2(g20329) );
  AND2_X1 AND2_2163( .ZN(g21334), .A1(g9310), .A2(g20330) );
  AND2_X1 AND2_2164( .ZN(g21335), .A1(g9248), .A2(g20331) );
  AND2_X1 AND2_2165( .ZN(g21336), .A1(g9203), .A2(g20332) );
  AND2_X1 AND2_2166( .ZN(g21337), .A1(g9471), .A2(g20334) );
  AND2_X1 AND2_2167( .ZN(g21338), .A1(g9391), .A2(g20335) );
  AND2_X1 AND2_2168( .ZN(g21339), .A1(g9326), .A2(g20336) );
  AND2_X1 AND2_2169( .ZN(g21340), .A1(g9737), .A2(g20340) );
  AND2_X1 AND2_2170( .ZN(g21341), .A1(g9613), .A2(g20341) );
  AND2_X1 AND2_2171( .ZN(g21342), .A1(g9488), .A2(g20342) );
  AND2_X1 AND2_2172( .ZN(g21343), .A1(g9161), .A2(g20344) );
  AND2_X1 AND2_2173( .ZN(g21344), .A1(g9150), .A2(g20345) );
  AND2_X1 AND2_2174( .ZN(g21345), .A1(g15096), .A2(g20346) );
  AND2_X1 AND2_2175( .ZN(g21349), .A1(g9248), .A2(g20347) );
  AND2_X1 AND2_2176( .ZN(g21350), .A1(g9203), .A2(g20348) );
  AND2_X1 AND2_2177( .ZN(g21351), .A1(g9174), .A2(g20349) );
  AND2_X1 AND2_2178( .ZN(g21352), .A1(g9391), .A2(g20350) );
  AND2_X1 AND2_2179( .ZN(g21353), .A1(g9326), .A2(g20351) );
  AND2_X1 AND2_2180( .ZN(g21354), .A1(g9264), .A2(g20352) );
  AND2_X1 AND2_2181( .ZN(g21355), .A1(g9613), .A2(g20354) );
  AND2_X1 AND2_2182( .ZN(g21356), .A1(g9488), .A2(g20355) );
  AND2_X1 AND2_2183( .ZN(g21357), .A1(g9407), .A2(g20356) );
  AND2_X1 AND2_2184( .ZN(g21360), .A1(g9507), .A2(g20361) );
  AND2_X1 AND2_2185( .ZN(g21361), .A1(g9150), .A2(g20362) );
  AND2_X1 AND2_2186( .ZN(g21362), .A1(g15096), .A2(g20363) );
  AND2_X1 AND2_2187( .ZN(g21363), .A1(g15022), .A2(g20364) );
  AND2_X1 AND2_2188( .ZN(g21367), .A1(g9203), .A2(g20366) );
  AND2_X1 AND2_2189( .ZN(g21368), .A1(g9174), .A2(g20367) );
  AND2_X1 AND2_2190( .ZN(g21369), .A1(g15188), .A2(g20368) );
  AND2_X1 AND2_2191( .ZN(g21370), .A1(g9326), .A2(g20369) );
  AND2_X1 AND2_2192( .ZN(g21371), .A1(g9264), .A2(g20370) );
  AND2_X1 AND2_2193( .ZN(g21372), .A1(g9216), .A2(g20371) );
  AND2_X1 AND2_2194( .ZN(g21373), .A1(g9488), .A2(g20372) );
  AND2_X1 AND2_2195( .ZN(g21374), .A1(g9407), .A2(g20373) );
  AND2_X1 AND2_2196( .ZN(g21375), .A1(g9342), .A2(g20374) );
  AND2_X1 AND2_2197( .ZN(g21378), .A1(g9507), .A2(g20378) );
  AND2_X1 AND2_2198( .ZN(g21379), .A1(g9427), .A2(g20379) );
  AND2_X1 AND2_2199( .ZN(g21380), .A1(g15096), .A2(g20380) );
  AND2_X1 AND2_2200( .ZN(g21381), .A1(g15022), .A2(g20381) );
  AND2_X1 AND2_2201( .ZN(g21388), .A1(g6201), .A2(g19657) );
  AND2_X1 AND2_2202( .ZN(g21389), .A1(g9649), .A2(g20384) );
  AND2_X1 AND2_2203( .ZN(g21390), .A1(g9174), .A2(g20385) );
  AND2_X1 AND2_2204( .ZN(g21391), .A1(g15188), .A2(g20386) );
  AND2_X1 AND2_2205( .ZN(g21392), .A1(g15118), .A2(g20387) );
  AND2_X1 AND2_2206( .ZN(g21393), .A1(g9264), .A2(g20389) );
  AND2_X1 AND2_2207( .ZN(g21394), .A1(g9216), .A2(g20390) );
  AND2_X1 AND2_2208( .ZN(g21395), .A1(g15274), .A2(g20391) );
  AND2_X1 AND2_2209( .ZN(g21396), .A1(g9407), .A2(g20392) );
  AND2_X1 AND2_2210( .ZN(g21397), .A1(g9342), .A2(g20393) );
  AND2_X1 AND2_2211( .ZN(g21398), .A1(g9277), .A2(g20394) );
  AND2_X1 AND2_2212( .ZN(g21401), .A1(g9507), .A2(g20397) );
  AND2_X1 AND2_2213( .ZN(g21402), .A1(g9427), .A2(g20398) );
  AND2_X1 AND2_2214( .ZN(g21403), .A1(g15022), .A2(g20399) );
  AND2_X1 AND2_2215( .ZN(g21410), .A1(g6363), .A2(g20402) );
  AND2_X1 AND2_2216( .ZN(g21411), .A1(g9649), .A2(g20403) );
  AND2_X1 AND2_2217( .ZN(g21412), .A1(g9569), .A2(g20404) );
  AND2_X1 AND2_2218( .ZN(g21413), .A1(g15188), .A2(g20405) );
  AND2_X1 AND2_2219( .ZN(g21414), .A1(g15118), .A2(g20406) );
  AND2_X1 AND2_2220( .ZN(g21418), .A1(g6290), .A2(g19705) );
  AND2_X1 AND2_2221( .ZN(g21419), .A1(g9795), .A2(g20409) );
  AND2_X1 AND2_2222( .ZN(g21420), .A1(g9216), .A2(g20410) );
  AND2_X1 AND2_2223( .ZN(g21421), .A1(g15274), .A2(g20411) );
  AND2_X1 AND2_2224( .ZN(g21422), .A1(g15210), .A2(g20412) );
  AND2_X1 AND2_2225( .ZN(g21423), .A1(g9342), .A2(g20414) );
  AND2_X1 AND2_2226( .ZN(g21424), .A1(g9277), .A2(g20415) );
  AND2_X1 AND2_2227( .ZN(g21425), .A1(g15366), .A2(g20416) );
  AND2_X1 AND2_2228( .ZN(g21428), .A1(g9427), .A2(g20420) );
  AND2_X1 AND2_2229( .ZN(g21438), .A1(g9649), .A2(g20422) );
  AND2_X1 AND2_2230( .ZN(g21439), .A1(g9569), .A2(g20423) );
  AND2_X1 AND2_2231( .ZN(g21440), .A1(g15118), .A2(g20424) );
  AND2_X1 AND2_2232( .ZN(g21444), .A1(g6568), .A2(g20427) );
  AND2_X1 AND2_2233( .ZN(g21445), .A1(g9795), .A2(g20428) );
  AND2_X1 AND2_2234( .ZN(g21446), .A1(g9711), .A2(g20429) );
  AND2_X1 AND2_2235( .ZN(g21447), .A1(g15274), .A2(g20430) );
  AND2_X1 AND2_2236( .ZN(g21448), .A1(g15210), .A2(g20431) );
  AND2_X1 AND2_2237( .ZN(g21452), .A1(g6427), .A2(g19749) );
  AND2_X1 AND2_2238( .ZN(g21453), .A1(g9941), .A2(g20434) );
  AND2_X1 AND2_2239( .ZN(g21454), .A1(g9277), .A2(g20435) );
  AND2_X1 AND2_2240( .ZN(g21455), .A1(g15366), .A2(g20436) );
  AND2_X1 AND2_2241( .ZN(g21456), .A1(g15296), .A2(g20437) );
  AND2_X1 AND2_2242( .ZN(g21476), .A1(g9569), .A2(g20442) );
  AND2_X1 AND2_2243( .ZN(g21480), .A1(g9795), .A2(g20444) );
  AND2_X1 AND2_2244( .ZN(g21481), .A1(g9711), .A2(g20445) );
  AND2_X1 AND2_2245( .ZN(g21482), .A1(g15210), .A2(g20446) );
  AND2_X1 AND2_2246( .ZN(g21486), .A1(g6832), .A2(g20449) );
  AND2_X1 AND2_2247( .ZN(g21487), .A1(g9941), .A2(g20450) );
  AND2_X1 AND2_2248( .ZN(g21488), .A1(g9857), .A2(g20451) );
  AND2_X1 AND2_2249( .ZN(g21489), .A1(g15366), .A2(g20452) );
  AND2_X1 AND2_2250( .ZN(g21490), .A1(g15296), .A2(g20453) );
  AND2_X1 AND2_2251( .ZN(g21494), .A1(g6632), .A2(g19792) );
  AND2_X1 AND2_2252( .ZN(g21497), .A1(g3006), .A2(g20456) );
  AND2_X1 AND2_2253( .ZN(g21517), .A1(g9711), .A2(g20461) );
  AND2_X1 AND2_2254( .ZN(g21521), .A1(g9941), .A2(g20463) );
  AND2_X1 AND2_2255( .ZN(g21522), .A1(g9857), .A2(g20464) );
  AND2_X1 AND2_2256( .ZN(g21523), .A1(g15296), .A2(g20465) );
  AND2_X1 AND2_2257( .ZN(g21527), .A1(g7134), .A2(g20468) );
  AND3_X1 AND3_202( .ZN(II28068), .A1(g17802), .A2(g18265), .A3(g17882) );
  AND4_X1 AND4_82( .ZN(g21533), .A1(g17724), .A2(g18179), .A3(g19799), .A4(II28068) );
  AND2_X1 AND2_2258( .ZN(g21553), .A1(g9857), .A2(g20476) );
  AND3_X1 AND3_203( .ZN(II28096), .A1(g13907), .A2(g14238), .A3(g13946) );
  AND4_X1 AND4_83( .ZN(g21564), .A1(g13886), .A2(g14153), .A3(g19799), .A4(II28096) );
  AND3_X1 AND3_204( .ZN(II28103), .A1(g17914), .A2(g18358), .A3(g17993) );
  AND4_X1 AND4_84( .ZN(g21569), .A1(g17825), .A2(g18286), .A3(g19843), .A4(II28103) );
  AND2_X1 AND2_2259( .ZN(g21589), .A1(g3002), .A2(g19890) );
  AND3_X1 AND3_205( .ZN(g21593), .A1(g16498), .A2(g19484), .A3(g14071) );
  AND3_X1 AND3_206( .ZN(II28126), .A1(g13963), .A2(g14360), .A3(g14016) );
  AND4_X1 AND4_85( .ZN(g21597), .A1(g13927), .A2(g14268), .A3(g19843), .A4(II28126) );
  AND3_X1 AND3_207( .ZN(II28133), .A1(g18025), .A2(g18453), .A3(g18110) );
  AND4_X1 AND4_86( .ZN(g21602), .A1(g17937), .A2(g18379), .A3(g19876), .A4(II28133) );
  AND2_X1 AND2_2260( .ZN(g21610), .A1(g7522), .A2(g20490) );
  AND2_X1 AND2_2261( .ZN(g21611), .A1(g7471), .A2(g19915) );
  AND3_X1 AND3_208( .ZN(g21622), .A1(g16520), .A2(g19505), .A3(g14186) );
  AND3_X1 AND3_209( .ZN(II28155), .A1(g14033), .A2(g14472), .A3(g14107) );
  AND4_X1 AND4_87( .ZN(g21626), .A1(g13983), .A2(g14390), .A3(g19876), .A4(II28155) );
  AND3_X1 AND3_210( .ZN(II28162), .A1(g18142), .A2(g18526), .A3(g18226) );
  AND4_X1 AND4_88( .ZN(g21631), .A1(g18048), .A2(g18474), .A3(g19907), .A4(II28162) );
  AND2_X1 AND2_2262( .ZN(g21635), .A1(g7549), .A2(g20496) );
  AND2_X1 AND2_2263( .ZN(g21639), .A1(g3398), .A2(g20500) );
  AND3_X1 AND3_211( .ZN(g21650), .A1(g16551), .A2(g19524), .A3(g14301) );
  AND3_X1 AND3_212( .ZN(II28181), .A1(g14124), .A2(g14559), .A3(g14222) );
  AND4_X1 AND4_89( .ZN(g21654), .A1(g14053), .A2(g14502), .A3(g19907), .A4(II28181) );
  AND2_X1 AND2_2264( .ZN(g21658), .A1(g2896), .A2(g20501) );
  AND2_X1 AND2_2265( .ZN(g21666), .A1(g3398), .A2(g20504) );
  AND2_X1 AND2_2266( .ZN(g21670), .A1(g3554), .A2(g20505) );
  AND3_X1 AND3_213( .ZN(g21681), .A1(g16583), .A2(g19534), .A3(g14423) );
  AND2_X1 AND2_2267( .ZN(g21687), .A1(g3398), .A2(g20516) );
  AND2_X1 AND2_2268( .ZN(g21695), .A1(g3554), .A2(g20517) );
  AND2_X1 AND2_2269( .ZN(g21699), .A1(g3710), .A2(g20518) );
  AND2_X1 AND2_2270( .ZN(g21707), .A1(g2892), .A2(g19978) );
  AND2_X1 AND2_2271( .ZN(g21723), .A1(g3554), .A2(g20534) );
  AND2_X1 AND2_2272( .ZN(g21731), .A1(g3710), .A2(g20535) );
  AND2_X1 AND2_2273( .ZN(g21735), .A1(g3866), .A2(g20536) );
  AND2_X1 AND2_2274( .ZN(g21749), .A1(g3710), .A2(g20553) );
  AND2_X1 AND2_2275( .ZN(g21757), .A1(g3866), .A2(g20554) );
  AND2_X1 AND2_2276( .ZN(g21758), .A1(g7607), .A2(g20045) );
  AND2_X1 AND2_2277( .ZN(g21773), .A1(g3866), .A2(g19078) );
  AND3_X1 AND3_214( .ZN(g21805), .A1(g16679), .A2(g19578), .A3(g14776) );
  AND3_X1 AND3_215( .ZN(g21812), .A1(g16705), .A2(g19608), .A3(g14811) );
  AND3_X1 AND3_216( .ZN(g21818), .A1(g16736), .A2(g19641), .A3(g14863) );
  AND3_X1 AND3_217( .ZN(g21822), .A1(g16778), .A2(g19681), .A3(g14936) );
  AND2_X1 AND2_2278( .ZN(g21891), .A1(g19302), .A2(g11749) );
  AND2_X1 AND2_2279( .ZN(g21892), .A1(g19288), .A2(g13011) );
  AND2_X1 AND2_2280( .ZN(g21899), .A1(g19323), .A2(g11749) );
  AND2_X1 AND2_2281( .ZN(g21900), .A1(g19306), .A2(g13011) );
  AND2_X1 AND2_2282( .ZN(g21906), .A1(g5715), .A2(g20513) );
  AND2_X1 AND2_2283( .ZN(g21911), .A1(g19350), .A2(g11749) );
  AND2_X1 AND2_2284( .ZN(g21912), .A1(g19327), .A2(g13011) );
  AND2_X1 AND2_2285( .ZN(g21913), .A1(g4456), .A2(g20519) );
  AND2_X1 AND2_2286( .ZN(g21920), .A1(g5773), .A2(g20531) );
  AND2_X1 AND2_2287( .ZN(g21925), .A1(g19384), .A2(g11749) );
  AND2_X1 AND2_2288( .ZN(g21926), .A1(g19354), .A2(g13011) );
  AND2_X1 AND2_2289( .ZN(g21931), .A1(g4632), .A2(g20539) );
  AND2_X1 AND2_2290( .ZN(g21938), .A1(g5832), .A2(g20550) );
  AND2_X1 AND2_2291( .ZN(g21990), .A1(g291), .A2(g21187) );
  AND2_X1 AND2_2292( .ZN(g22004), .A1(g978), .A2(g21202) );
  AND2_X1 AND2_2293( .ZN(g22015), .A1(g1672), .A2(g21217) );
  AND2_X1 AND2_2294( .ZN(g22020), .A1(g2366), .A2(g21225) );
  AND3_X1 AND3_218( .ZN(II28582), .A1(g19141), .A2(g21133), .A3(g21116) );
  AND4_X1 AND4_90( .ZN(g22036), .A1(g21104), .A2(g21095), .A3(g21084), .A4(II28582) );
  AND3_X1 AND3_219( .ZN(II28594), .A1(g21167), .A2(g21147), .A3(g21134) );
  AND4_X1 AND4_91( .ZN(g22046), .A1(g21117), .A2(g21105), .A3(g21096), .A4(II28594) );
  AND3_X1 AND3_220( .ZN(II28609), .A1(g21183), .A2(g21168), .A3(g21148) );
  AND4_X1 AND4_92( .ZN(g22062), .A1(g21135), .A2(g21118), .A3(g21106), .A4(II28609) );
  AND2_X1 AND2_2295( .ZN(g22187), .A1(g21564), .A2(g20986) );
  AND2_X1 AND2_2296( .ZN(g22196), .A1(g21597), .A2(g21012) );
  AND2_X1 AND2_2297( .ZN(g22201), .A1(g21271), .A2(g16881) );
  AND2_X1 AND2_2298( .ZN(g22202), .A1(g21626), .A2(g21036) );
  AND2_X1 AND2_2299( .ZN(g22206), .A1(g21895), .A2(g11976) );
  AND2_X1 AND2_2300( .ZN(g22207), .A1(g21278), .A2(g16910) );
  AND2_X1 AND2_2301( .ZN(g22208), .A1(g21654), .A2(g21057) );
  AND2_X1 AND2_2302( .ZN(g22211), .A1(g21661), .A2(g12027) );
  AND2_X1 AND2_2303( .ZN(g22214), .A1(g21907), .A2(g12045) );
  AND2_X1 AND2_2304( .ZN(g22215), .A1(g21285), .A2(g16940) );
  AND2_X1 AND2_2305( .ZN(g22220), .A1(g21690), .A2(g12091) );
  AND2_X1 AND2_2306( .ZN(g22223), .A1(g21921), .A2(g12109) );
  AND2_X1 AND2_2307( .ZN(g22224), .A1(g21293), .A2(g16971) );
  AND2_X1 AND2_2308( .ZN(g22228), .A1(g21716), .A2(g12136) );
  AND2_X1 AND2_2309( .ZN(g22229), .A1(g21661), .A2(g12139) );
  AND2_X1 AND2_2310( .ZN(g22235), .A1(g21726), .A2(g12163) );
  AND2_X1 AND2_2311( .ZN(g22238), .A1(g21939), .A2(g12181) );
  AND2_X1 AND2_2312( .ZN(g22244), .A1(g21742), .A2(g12198) );
  AND2_X1 AND2_2313( .ZN(g22245), .A1(g21690), .A2(g12201) );
  AND2_X1 AND2_2314( .ZN(g22250), .A1(g21752), .A2(g12225) );
  AND2_X1 AND2_2315( .ZN(g22254), .A1(g21716), .A2(g12239) );
  AND2_X1 AND2_2316( .ZN(g22255), .A1(g21661), .A2(g12242) );
  AND2_X1 AND2_2317( .ZN(g22264), .A1(g21766), .A2(g12253) );
  AND2_X1 AND2_2318( .ZN(g22265), .A1(g21726), .A2(g12256) );
  AND2_X1 AND2_2319( .ZN(g22270), .A1(g92), .A2(g21529) );
  AND2_X1 AND2_2320( .ZN(g22272), .A1(g21742), .A2(g12282) );
  AND2_X1 AND2_2321( .ZN(g22273), .A1(g21690), .A2(g12285) );
  AND2_X1 AND2_2322( .ZN(g22281), .A1(g21782), .A2(g12296) );
  AND2_X1 AND2_2323( .ZN(g22282), .A1(g21752), .A2(g12299) );
  AND2_X1 AND2_2324( .ZN(g22285), .A1(g21716), .A2(g12312) );
  AND2_X1 AND2_2325( .ZN(g22289), .A1(g780), .A2(g21565) );
  AND2_X1 AND2_2326( .ZN(g22291), .A1(g21766), .A2(g12318) );
  AND2_X1 AND2_2327( .ZN(g22292), .A1(g21726), .A2(g12321) );
  AND2_X1 AND2_2328( .ZN(g22305), .A1(g21742), .A2(g12340) );
  AND2_X1 AND2_2329( .ZN(g22309), .A1(g1466), .A2(g21598) );
  AND2_X1 AND2_2330( .ZN(g22311), .A1(g21782), .A2(g12346) );
  AND2_X1 AND2_2331( .ZN(g22312), .A1(g21752), .A2(g12349) );
  AND2_X1 AND2_2332( .ZN(g22333), .A1(g21766), .A2(g12370) );
  AND2_X1 AND2_2333( .ZN(g22337), .A1(g2160), .A2(g21627) );
  AND2_X1 AND2_2334( .ZN(g22340), .A1(g88), .A2(g21184) );
  AND2_X1 AND2_2335( .ZN(g22358), .A1(g21782), .A2(g12389) );
  AND2_X1 AND2_2336( .ZN(g22363), .A1(g776), .A2(g21199) );
  AND2_X1 AND2_2337( .ZN(g22383), .A1(g1462), .A2(g21214) );
  AND2_X1 AND2_2338( .ZN(g22398), .A1(g2156), .A2(g21222) );
  AND2_X1 AND2_2339( .ZN(g22483), .A1(g646), .A2(g21861) );
  AND2_X1 AND2_2340( .ZN(g22515), .A1(g13873), .A2(g21382) );
  AND2_X1 AND2_2341( .ZN(g22516), .A1(g20885), .A2(g17442) );
  AND2_X1 AND2_2342( .ZN(g22517), .A1(g21895), .A2(g12608) );
  AND2_X1 AND2_2343( .ZN(g22526), .A1(g1332), .A2(g21867) );
  AND2_X1 AND2_2344( .ZN(g22546), .A1(g13886), .A2(g21404) );
  AND2_X1 AND2_2345( .ZN(g22555), .A1(g13895), .A2(g21415) );
  AND2_X1 AND2_2346( .ZN(g22556), .A1(g20904), .A2(g17523) );
  AND2_X1 AND2_2347( .ZN(g22557), .A1(g21907), .A2(g12654) );
  AND2_X1 AND2_2348( .ZN(g22566), .A1(g2026), .A2(g21872) );
  AND2_X1 AND2_2349( .ZN(g22577), .A1(g13907), .A2(g21429) );
  AND2_X1 AND2_2350( .ZN(g22581), .A1(g21895), .A2(g12699) );
  AND2_X1 AND2_2351( .ZN(g22587), .A1(g13927), .A2(g21441) );
  AND2_X1 AND2_2352( .ZN(g22595), .A1(g13936), .A2(g21449) );
  AND2_X1 AND2_2353( .ZN(g22596), .A1(g20928), .A2(g17613) );
  AND2_X1 AND2_2354( .ZN(g22597), .A1(g21921), .A2(g12708) );
  AND2_X1 AND2_2355( .ZN(g22606), .A1(g2720), .A2(g21876) );
  AND2_X1 AND2_2356( .ZN(g22607), .A1(g13946), .A2(g21458) );
  AND2_X1 AND2_2357( .ZN(g22610), .A1(g660), .A2(g21473) );
  AND2_X1 AND2_2358( .ZN(g22614), .A1(g13963), .A2(g21477) );
  AND2_X2 AND2_2359( .ZN(g22618), .A1(g21907), .A2(g12756) );
  AND2_X2 AND2_2360( .ZN(g22624), .A1(g13983), .A2(g21483) );
  AND2_X2 AND2_2361( .ZN(g22632), .A1(g13992), .A2(g21491) );
  AND2_X2 AND2_2362( .ZN(g22633), .A1(g20956), .A2(g17710) );
  AND2_X1 AND2_2363( .ZN(g22634), .A1(g21939), .A2(g12765) );
  AND2_X1 AND2_2364( .ZN(g22637), .A1(g20841), .A2(g10927) );
  AND2_X1 AND2_2365( .ZN(g22638), .A1(g14001), .A2(g21498) );
  AND2_X1 AND2_2366( .ZN(g22643), .A1(g14016), .A2(g21505) );
  AND2_X1 AND2_2367( .ZN(g22646), .A1(g1346), .A2(g21514) );
  AND2_X1 AND2_2368( .ZN(g22650), .A1(g14033), .A2(g21518) );
  AND2_X1 AND2_2369( .ZN(g22654), .A1(g21921), .A2(g12798) );
  AND2_X1 AND2_2370( .ZN(g22660), .A1(g14053), .A2(g21524) );
  AND2_X1 AND2_2371( .ZN(g22665), .A1(g20920), .A2(g6153) );
  AND2_X1 AND2_2372( .ZN(g22666), .A1(g21825), .A2(g20014) );
  AND2_X1 AND2_2373( .ZN(g22667), .A1(g14062), .A2(g21530) );
  AND2_X1 AND2_2374( .ZN(g22674), .A1(g14092), .A2(g21537) );
  AND2_X1 AND2_2375( .ZN(g22679), .A1(g14107), .A2(g21541) );
  AND2_X1 AND2_2376( .ZN(g22682), .A1(g2040), .A2(g21550) );
  AND2_X1 AND2_2377( .ZN(g22686), .A1(g14124), .A2(g21554) );
  AND2_X1 AND2_2378( .ZN(g22690), .A1(g21939), .A2(g12837) );
  AND2_X1 AND2_2379( .ZN(g22699), .A1(g7338), .A2(g21883) );
  AND2_X1 AND2_2380( .ZN(g22700), .A1(g7146), .A2(g21558) );
  AND2_X1 AND2_2381( .ZN(g22701), .A1(g18174), .A2(g21561) );
  AND2_X1 AND2_2382( .ZN(g22707), .A1(g14177), .A2(g21566) );
  AND2_X1 AND2_2383( .ZN(g22714), .A1(g14207), .A2(g21573) );
  AND2_X1 AND2_2384( .ZN(g22719), .A1(g14222), .A2(g21577) );
  AND2_X1 AND2_2385( .ZN(g22722), .A1(g2734), .A2(g21586) );
  AND2_X1 AND2_2386( .ZN(g22726), .A1(g3036), .A2(g21886) );
  AND2_X1 AND2_2387( .ZN(g22727), .A1(g14238), .A2(g21590) );
  AND2_X1 AND2_2388( .ZN(g22732), .A1(g18281), .A2(g21594) );
  AND2_X1 AND2_2389( .ZN(g22738), .A1(g14292), .A2(g21599) );
  AND2_X1 AND2_2390( .ZN(g22745), .A1(g14322), .A2(g21606) );
  AND2_X1 AND2_2391( .ZN(g22754), .A1(g14342), .A2(g21612) );
  AND2_X1 AND2_2392( .ZN(g22759), .A1(g14360), .A2(g21619) );
  AND2_X1 AND2_2393( .ZN(g22764), .A1(g18374), .A2(g21623) );
  AND2_X1 AND2_2394( .ZN(g22770), .A1(g14414), .A2(g21628) );
  AND2_X1 AND2_2395( .ZN(g22788), .A1(g14454), .A2(g21640) );
  AND2_X1 AND2_2396( .ZN(g22793), .A1(g14472), .A2(g21647) );
  AND2_X1 AND2_2397( .ZN(g22798), .A1(g18469), .A2(g21651) );
  AND2_X1 AND2_2398( .ZN(g22804), .A1(g2920), .A2(g21655) );
  AND2_X1 AND2_2399( .ZN(g22830), .A1(g14541), .A2(g21671) );
  AND2_X1 AND2_2400( .ZN(g22835), .A1(g14559), .A2(g21678) );
  AND2_X1 AND2_2401( .ZN(g22841), .A1(g7583), .A2(g21902) );
  AND2_X1 AND2_2402( .ZN(g22842), .A1(g3032), .A2(g21682) );
  AND2_X1 AND2_2403( .ZN(g22869), .A1(g14596), .A2(g21700) );
  AND2_X1 AND2_2404( .ZN(g22874), .A1(g7587), .A2(g21708) );
  AND2_X1 AND2_2405( .ZN(g22906), .A1(g2924), .A2(g21927) );
  AND2_X1 AND2_2406( .ZN(g22984), .A1(g16840), .A2(g21400) );
  AND2_X1 AND2_2407( .ZN(g23104), .A1(g20842), .A2(g15859) );
  AND2_X1 AND2_2408( .ZN(g23106), .A1(g5857), .A2(g21050) );
  AND2_X1 AND2_2409( .ZN(g23118), .A1(g20850), .A2(g15890) );
  AND2_X1 AND2_2410( .ZN(g23119), .A1(g5904), .A2(g21069) );
  AND2_X1 AND2_2411( .ZN(g23127), .A1(g20858), .A2(g15923) );
  AND2_X1 AND2_2412( .ZN(g23128), .A1(g5943), .A2(g21079) );
  AND2_X1 AND2_2413( .ZN(g23138), .A1(g20866), .A2(g15952) );
  AND2_X1 AND2_2414( .ZN(g23139), .A1(g5977), .A2(g21093) );
  AND2_X1 AND2_2415( .ZN(g23409), .A1(g21533), .A2(g22408) );
  AND2_X1 AND2_2416( .ZN(g23414), .A1(g21569), .A2(g22421) );
  AND2_X1 AND2_2417( .ZN(g23419), .A1(g22755), .A2(g19577) );
  AND2_X1 AND2_2418( .ZN(g23423), .A1(g21602), .A2(g22443) );
  AND2_X1 AND2_2419( .ZN(g23428), .A1(g22789), .A2(g19607) );
  AND2_X1 AND2_2420( .ZN(g23432), .A1(g21631), .A2(g22476) );
  AND2_X1 AND2_2421( .ZN(g23434), .A1(g22831), .A2(g19640) );
  AND2_X1 AND2_2422( .ZN(g23440), .A1(g22870), .A2(g19680) );
  AND2_X1 AND2_2423( .ZN(g23451), .A1(g18552), .A2(g22547) );
  AND2_X1 AND2_2424( .ZN(g23458), .A1(g18602), .A2(g22588) );
  AND2_X1 AND2_2425( .ZN(g23462), .A1(g17988), .A2(g22609) );
  AND2_X1 AND2_2426( .ZN(g23467), .A1(g18634), .A2(g22625) );
  AND2_X1 AND2_2427( .ZN(g23471), .A1(g18105), .A2(g22645) );
  AND2_X1 AND2_2428( .ZN(g23476), .A1(g18643), .A2(g22661) );
  AND2_X1 AND2_2429( .ZN(g23483), .A1(g22945), .A2(g8847) );
  AND2_X1 AND2_2430( .ZN(g23484), .A1(g18221), .A2(g22681) );
  AND2_X1 AND2_2431( .ZN(g23494), .A1(g18328), .A2(g22721) );
  AND2_X1 AND2_2432( .ZN(g23496), .A1(g5802), .A2(g22300) );
  AND2_X1 AND2_2433( .ZN(g23510), .A1(g5890), .A2(g22753) );
  AND2_X1 AND2_2434( .ZN(g23512), .A1(g5858), .A2(g22328) );
  AND2_X1 AND2_2435( .ZN(g23525), .A1(g5929), .A2(g22787) );
  AND2_X1 AND2_2436( .ZN(g23527), .A1(g5905), .A2(g22353) );
  AND2_X1 AND2_2437( .ZN(g23536), .A1(g5963), .A2(g22829) );
  AND2_X1 AND2_2438( .ZN(g23538), .A1(g5944), .A2(g22376) );
  AND2_X1 AND2_2439( .ZN(g23544), .A1(g5992), .A2(g22868) );
  AND2_X1 AND2_2440( .ZN(g23547), .A1(g8062), .A2(g22405) );
  AND2_X1 AND2_2441( .ZN(g23550), .A1(g8132), .A2(g22409) );
  AND2_X1 AND2_2442( .ZN(g23551), .A1(g8135), .A2(g22412) );
  AND2_X1 AND2_2443( .ZN(g23552), .A1(g6136), .A2(g22415) );
  AND2_X1 AND2_2444( .ZN(g23554), .A1(g8147), .A2(g22418) );
  AND2_X1 AND2_2445( .ZN(g23558), .A1(g8200), .A2(g22422) );
  AND2_X1 AND2_2446( .ZN(g23559), .A1(g8203), .A2(g22425) );
  AND2_X1 AND2_2447( .ZN(g23560), .A1(g8206), .A2(g22428) );
  AND2_X1 AND2_2448( .ZN(g23563), .A1(g8218), .A2(g22431) );
  AND2_X1 AND2_2449( .ZN(g23564), .A1(g8221), .A2(g22434) );
  AND2_X1 AND2_2450( .ZN(g23565), .A1(g6146), .A2(g22437) );
  AND2_X1 AND2_2451( .ZN(g23567), .A1(g8233), .A2(g22440) );
  AND2_X1 AND2_2452( .ZN(g23571), .A1(g3931), .A2(g22445) );
  AND2_X1 AND2_2453( .ZN(g23572), .A1(g3934), .A2(g22448) );
  AND2_X1 AND2_2454( .ZN(g23573), .A1(g3937), .A2(g22451) );
  AND2_X1 AND2_2455( .ZN(g23577), .A1(g3957), .A2(g22455) );
  AND2_X1 AND2_2456( .ZN(g23578), .A1(g3960), .A2(g22458) );
  AND2_X1 AND2_2457( .ZN(g23579), .A1(g3963), .A2(g22461) );
  AND2_X1 AND2_2458( .ZN(g23582), .A1(g3975), .A2(g22464) );
  AND2_X1 AND2_2459( .ZN(g23583), .A1(g3978), .A2(g22467) );
  AND2_X1 AND2_2460( .ZN(g23584), .A1(g6167), .A2(g22470) );
  AND2_X1 AND2_2461( .ZN(g23586), .A1(g3990), .A2(g22473) );
  AND2_X1 AND2_2462( .ZN(g23590), .A1(g4009), .A2(g22477) );
  AND2_X1 AND2_2463( .ZN(g23591), .A1(g4012), .A2(g22480) );
  AND2_X1 AND2_2464( .ZN(g23592), .A1(g17640), .A2(g22986) );
  AND2_X1 AND2_2465( .ZN(g23593), .A1(g22845), .A2(g20365) );
  AND2_X1 AND2_2466( .ZN(g23598), .A1(g4038), .A2(g22484) );
  AND2_X1 AND2_2467( .ZN(g23599), .A1(g4041), .A2(g22487) );
  AND2_X1 AND2_2468( .ZN(g23600), .A1(g4044), .A2(g22490) );
  AND2_X1 AND2_2469( .ZN(g23604), .A1(g4064), .A2(g22494) );
  AND2_X1 AND2_2470( .ZN(g23605), .A1(g4067), .A2(g22497) );
  AND2_X1 AND2_2471( .ZN(g23606), .A1(g4070), .A2(g22500) );
  AND2_X1 AND2_2472( .ZN(g23609), .A1(g4082), .A2(g22503) );
  AND2_X1 AND2_2473( .ZN(g23610), .A1(g4085), .A2(g22506) );
  AND2_X1 AND2_2474( .ZN(g23611), .A1(g6194), .A2(g22509) );
  AND2_X1 AND2_2475( .ZN(g23615), .A1(g4107), .A2(g22512) );
  AND2_X1 AND2_2476( .ZN(g23616), .A1(g17724), .A2(g22988) );
  AND2_X1 AND2_2477( .ZN(g23617), .A1(g22810), .A2(g20382) );
  AND2_X1 AND2_2478( .ZN(g23618), .A1(g22608), .A2(g20383) );
  AND2_X1 AND2_2479( .ZN(g23622), .A1(g4136), .A2(g22520) );
  AND2_X1 AND2_2480( .ZN(g23623), .A1(g4139), .A2(g22523) );
  AND2_X1 AND2_2481( .ZN(g23624), .A1(g17741), .A2(g22989) );
  AND2_X1 AND2_2482( .ZN(g23625), .A1(g22880), .A2(g20388) );
  AND2_X1 AND2_2483( .ZN(g23630), .A1(g4165), .A2(g22527) );
  AND2_X1 AND2_2484( .ZN(g23631), .A1(g4168), .A2(g22530) );
  AND2_X1 AND2_2485( .ZN(g23632), .A1(g4171), .A2(g22533) );
  AND2_X1 AND2_2486( .ZN(g23636), .A1(g4191), .A2(g22537) );
  AND2_X1 AND2_2487( .ZN(g23637), .A1(g4194), .A2(g22540) );
  AND2_X1 AND2_2488( .ZN(g23638), .A1(g4197), .A2(g22543) );
  AND2_X1 AND2_2489( .ZN(g23639), .A1(g21825), .A2(g22805) );
  AND2_X1 AND2_2490( .ZN(g23643), .A1(g17802), .A2(g22991) );
  AND2_X1 AND2_2491( .ZN(g23659), .A1(g22784), .A2(g17500) );
  AND2_X1 AND2_2492( .ZN(g23664), .A1(g4246), .A2(g22552) );
  AND2_X1 AND2_2493( .ZN(g23665), .A1(g17825), .A2(g22995) );
  AND2_X1 AND2_2494( .ZN(g23666), .A1(g22851), .A2(g20407) );
  AND2_X1 AND2_2495( .ZN(g23667), .A1(g22644), .A2(g20408) );
  AND2_X1 AND2_2496( .ZN(g23671), .A1(g4275), .A2(g22560) );
  AND2_X1 AND2_2497( .ZN(g23672), .A1(g4278), .A2(g22563) );
  AND2_X1 AND2_2498( .ZN(g23673), .A1(g17842), .A2(g22996) );
  AND2_X1 AND2_2499( .ZN(g23674), .A1(g22915), .A2(g20413) );
  AND2_X1 AND2_2500( .ZN(g23679), .A1(g4304), .A2(g22567) );
  AND2_X1 AND2_2501( .ZN(g23680), .A1(g4307), .A2(g22570) );
  AND2_X1 AND2_2502( .ZN(g23681), .A1(g4310), .A2(g22573) );
  AND2_X1 AND2_2503( .ZN(g23686), .A1(g17882), .A2(g22998) );
  AND2_X1 AND2_2504( .ZN(g23687), .A1(g22668), .A2(g17570) );
  AND2_X1 AND2_2505( .ZN(g23689), .A1(g6513), .A2(g23001) );
  AND2_X1 AND2_2506( .ZN(g23693), .A1(g17914), .A2(g23002) );
  AND2_X1 AND2_2507( .ZN(g23709), .A1(g22826), .A2(g17591) );
  AND2_X1 AND2_2508( .ZN(g23714), .A1(g4401), .A2(g22592) );
  AND2_X1 AND2_2509( .ZN(g23715), .A1(g17937), .A2(g23006) );
  AND2_X1 AND2_2510( .ZN(g23716), .A1(g22886), .A2(g20432) );
  AND2_X1 AND2_2511( .ZN(g23717), .A1(g22680), .A2(g20433) );
  AND2_X1 AND2_2512( .ZN(g23721), .A1(g4430), .A2(g22600) );
  AND2_X1 AND2_2513( .ZN(g23722), .A1(g4433), .A2(g22603) );
  AND2_X1 AND2_2514( .ZN(g23723), .A1(g17954), .A2(g23007) );
  AND2_X1 AND2_2515( .ZN(g23724), .A1(g22940), .A2(g20438) );
  AND2_X1 AND2_2516( .ZN(g23726), .A1(g21825), .A2(g22843) );
  AND2_X1 AND2_2517( .ZN(g23734), .A1(g17974), .A2(g23008) );
  AND2_X1 AND2_2518( .ZN(g23735), .A1(g22949), .A2(g9450) );
  AND2_X1 AND2_2519( .ZN(g23740), .A1(g17993), .A2(g23012) );
  AND2_X1 AND2_2520( .ZN(g23741), .A1(g22708), .A2(g17667) );
  AND2_X1 AND2_2521( .ZN(g23743), .A1(g6777), .A2(g23015) );
  AND2_X1 AND2_2522( .ZN(g23747), .A1(g18025), .A2(g23016) );
  AND2_X1 AND2_2523( .ZN(g23763), .A1(g22865), .A2(g17688) );
  AND2_X1 AND2_2524( .ZN(g23768), .A1(g4570), .A2(g22629) );
  AND2_X1 AND2_2525( .ZN(g23769), .A1(g18048), .A2(g23020) );
  AND2_X1 AND2_2526( .ZN(g23770), .A1(g22921), .A2(g20454) );
  AND2_X1 AND2_2527( .ZN(g23771), .A1(g22720), .A2(g20455) );
  AND2_X1 AND2_2528( .ZN(g23772), .A1(g21825), .A2(g22875) );
  AND2_X1 AND2_2529( .ZN(g23776), .A1(g18074), .A2(g23021) );
  AND2_X1 AND2_2530( .ZN(g23777), .A1(g22949), .A2(g9528) );
  AND2_X1 AND2_2531( .ZN(g23778), .A1(g22954), .A2(g9531) );
  AND2_X1 AND2_2532( .ZN(g23789), .A1(g18091), .A2(g23024) );
  AND2_X2 AND2_2533( .ZN(g23790), .A1(g22958), .A2(g9592) );
  AND2_X2 AND2_2534( .ZN(g23795), .A1(g18110), .A2(g23028) );
  AND2_X2 AND2_2535( .ZN(g23796), .A1(g22739), .A2(g17767) );
  AND2_X1 AND2_2536( .ZN(g23798), .A1(g7079), .A2(g23031) );
  AND2_X1 AND2_2537( .ZN(g23802), .A1(g18142), .A2(g23032) );
  AND2_X1 AND2_2538( .ZN(g23818), .A1(g22900), .A2(g17788) );
  AND2_X1 AND2_2539( .ZN(g23820), .A1(g3013), .A2(g23036) );
  AND2_X1 AND2_2540( .ZN(g23822), .A1(g14148), .A2(g23037) );
  AND2_X1 AND2_2541( .ZN(g23824), .A1(g22949), .A2(g9641) );
  AND2_X1 AND2_2542( .ZN(g23825), .A1(g22954), .A2(g9644) );
  AND2_X1 AND2_2543( .ZN(g23829), .A1(g18190), .A2(g23038) );
  AND2_X1 AND2_2544( .ZN(g23830), .A1(g22958), .A2(g9670) );
  AND2_X1 AND2_2545( .ZN(g23831), .A1(g22962), .A2(g9673) );
  AND2_X1 AND2_2546( .ZN(g23842), .A1(g18207), .A2(g23041) );
  AND2_X1 AND2_2547( .ZN(g23843), .A1(g22966), .A2(g9734) );
  AND2_X1 AND2_2548( .ZN(g23848), .A1(g18226), .A2(g23045) );
  AND2_X1 AND2_2549( .ZN(g23849), .A1(g22771), .A2(g17868) );
  AND2_X1 AND2_2550( .ZN(g23851), .A1(g7329), .A2(g23048) );
  AND2_X1 AND2_2551( .ZN(g23852), .A1(g19179), .A2(g22696) );
  AND2_X1 AND2_2552( .ZN(g23854), .A1(g18265), .A2(g23049) );
  AND2_X1 AND2_2553( .ZN(g23855), .A1(g22954), .A2(g9767) );
  AND2_X1 AND2_2554( .ZN(g23857), .A1(g14263), .A2(g23056) );
  AND2_X1 AND2_2555( .ZN(g23859), .A1(g22958), .A2(g9787) );
  AND2_X1 AND2_2556( .ZN(g23860), .A1(g22962), .A2(g9790) );
  AND2_X1 AND2_2557( .ZN(g23864), .A1(g18297), .A2(g23057) );
  AND2_X1 AND2_2558( .ZN(g23865), .A1(g22966), .A2(g9816) );
  AND2_X1 AND2_2559( .ZN(g23866), .A1(g22971), .A2(g9819) );
  AND2_X1 AND2_2560( .ZN(g23877), .A1(g18314), .A2(g23060) );
  AND2_X1 AND2_2561( .ZN(g23878), .A1(g22975), .A2(g9880) );
  AND2_X1 AND2_2562( .ZN(g23886), .A1(g18341), .A2(g23064) );
  AND2_X1 AND2_2563( .ZN(g23888), .A1(g18358), .A2(g23069) );
  AND2_X1 AND2_2564( .ZN(g23889), .A1(g22962), .A2(g9913) );
  AND2_X1 AND2_2565( .ZN(g23891), .A1(g14385), .A2(g23074) );
  AND2_X1 AND2_2566( .ZN(g23893), .A1(g22966), .A2(g9933) );
  AND2_X1 AND2_2567( .ZN(g23894), .A1(g22971), .A2(g9936) );
  AND2_X1 AND2_2568( .ZN(g23898), .A1(g18390), .A2(g23075) );
  AND2_X1 AND2_2569( .ZN(g23899), .A1(g22975), .A2(g9962) );
  AND2_X1 AND2_2570( .ZN(g23900), .A1(g22980), .A2(g9965) );
  AND2_X1 AND2_2571( .ZN(g23904), .A1(g3010), .A2(g22750) );
  AND2_X1 AND2_2572( .ZN(g23907), .A1(g18436), .A2(g23079) );
  AND2_X1 AND2_2573( .ZN(g23909), .A1(g18453), .A2(g23082) );
  AND2_X1 AND2_2574( .ZN(g23910), .A1(g22971), .A2(g10067) );
  AND2_X1 AND2_2575( .ZN(g23912), .A1(g14497), .A2(g23087) );
  AND2_X1 AND2_2576( .ZN(g23914), .A1(g22975), .A2(g10087) );
  AND2_X1 AND2_2577( .ZN(g23915), .A1(g22980), .A2(g10090) );
  AND2_X1 AND2_2578( .ZN(g23917), .A1(g7545), .A2(g23088) );
  AND2_X1 AND2_2579( .ZN(g23939), .A1(g18509), .A2(g23095) );
  AND2_X1 AND2_2580( .ZN(g23941), .A1(g18526), .A2(g23098) );
  AND2_X1 AND2_2581( .ZN(g23942), .A1(g22980), .A2(g10176) );
  AND2_X1 AND2_2582( .ZN(g23944), .A1(g7570), .A2(g23103) );
  AND2_X1 AND2_2583( .ZN(g23971), .A1(g18573), .A2(g23112) );
  AND2_X1 AND2_2584( .ZN(g23972), .A1(g2903), .A2(g23115) );
  AND2_X1 AND2_2585( .ZN(g24029), .A1(g2900), .A2(g22903) );
  AND2_X1 AND2_2586( .ZN(g24211), .A1(g22014), .A2(g10969) );
  AND2_X1 AND2_2587( .ZN(g24217), .A1(g22825), .A2(g10999) );
  AND2_X1 AND2_2588( .ZN(g24221), .A1(g22979), .A2(g11042) );
  AND2_X1 AND2_2589( .ZN(g24224), .A1(g22219), .A2(g11045) );
  AND2_X1 AND2_2590( .ZN(g24229), .A1(g22232), .A2(g11105) );
  AND2_X1 AND2_2591( .ZN(g24236), .A1(g22243), .A2(g11157) );
  AND2_X1 AND2_2592( .ZN(g24241), .A1(g22259), .A2(g11228) );
  AND2_X1 AND2_2593( .ZN(g24246), .A1(g21982), .A2(g11291) );
  AND2_X1 AND2_2594( .ZN(g24247), .A1(g22551), .A2(g11297) );
  AND2_X1 AND2_2595( .ZN(g24253), .A1(g21995), .A2(g11370) );
  AND2_X1 AND2_2596( .ZN(g24256), .A1(g22003), .A2(g11438) );
  AND3_X1 AND3_221( .ZN(g24427), .A1(g17086), .A2(g24134), .A3(g13626) );
  AND2_X1 AND2_2597( .ZN(g24429), .A1(g24115), .A2(g13614) );
  AND3_X1 AND3_222( .ZN(g24431), .A1(g17124), .A2(g24153), .A3(g13637) );
  AND3_X1 AND3_223( .ZN(g24432), .A1(g14642), .A2(g15904), .A3(g24115) );
  AND2_X1 AND2_2598( .ZN(g24433), .A1(g24134), .A2(g13626) );
  AND3_X1 AND3_224( .ZN(g24435), .A1(g17151), .A2(g24168), .A3(g13649) );
  AND3_X1 AND3_225( .ZN(g24436), .A1(g14669), .A2(g15933), .A3(g24134) );
  AND2_X1 AND2_2599( .ZN(g24437), .A1(g24153), .A2(g13637) );
  AND3_X1 AND3_226( .ZN(g24439), .A1(g14703), .A2(g15962), .A3(g24153) );
  AND2_X1 AND2_2600( .ZN(g24440), .A1(g24168), .A2(g13649) );
  AND3_X1 AND3_227( .ZN(g24441), .A1(g14737), .A2(g15981), .A3(g24168) );
  AND3_X1 AND3_228( .ZN(g24478), .A1(g23545), .A2(g21119), .A3(g21227) );
  AND3_X1 AND3_229( .ZN(g24529), .A1(g19933), .A2(g17896), .A3(g23403) );
  AND3_X1 AND3_230( .ZN(g24540), .A1(g18548), .A2(g23089), .A3(g23403) );
  AND3_X1 AND3_231( .ZN(g24541), .A1(g23420), .A2(g17896), .A3(g23052) );
  AND3_X1 AND3_232( .ZN(g24542), .A1(g19950), .A2(g18007), .A3(g23410) );
  AND3_X1 AND3_233( .ZN(g24550), .A1(g18548), .A2(g23420), .A3(g19948) );
  AND3_X1 AND3_234( .ZN(g24552), .A1(g18598), .A2(g23107), .A3(g23410) );
  AND3_X1 AND3_235( .ZN(g24553), .A1(g23429), .A2(g18007), .A3(g23071) );
  AND3_X1 AND3_236( .ZN(g24554), .A1(g19977), .A2(g18124), .A3(g23415) );
  AND2_X1 AND2_2601( .ZN(g24559), .A1(g79), .A2(g23448) );
  AND3_X1 AND3_237( .ZN(g24561), .A1(g18598), .A2(g23429), .A3(g19975) );
  AND3_X1 AND3_238( .ZN(g24563), .A1(g18630), .A2(g23120), .A3(g23415) );
  AND3_X1 AND3_239( .ZN(g24564), .A1(g23435), .A2(g18124), .A3(g23084) );
  AND3_X1 AND3_240( .ZN(g24565), .A1(g20007), .A2(g18240), .A3(g23424) );
  AND2_X1 AND2_2602( .ZN(g24569), .A1(g767), .A2(g23455) );
  AND3_X1 AND3_241( .ZN(g24571), .A1(g18630), .A2(g23435), .A3(g20005) );
  AND3_X1 AND3_242( .ZN(g24573), .A1(g18639), .A2(g23129), .A3(g23424) );
  AND3_X1 AND3_243( .ZN(g24574), .A1(g23441), .A2(g18240), .A3(g23100) );
  AND2_X1 AND2_2603( .ZN(g24578), .A1(g1453), .A2(g23464) );
  AND3_X1 AND3_244( .ZN(g24580), .A1(g18639), .A2(g23441), .A3(g20043) );
  AND2_X1 AND2_2604( .ZN(g24585), .A1(g2147), .A2(g23473) );
  AND2_X1 AND2_2605( .ZN(g24590), .A1(g23486), .A2(g23478) );
  AND2_X1 AND2_2606( .ZN(g24591), .A1(g83), .A2(g23853) );
  AND2_X1 AND2_2607( .ZN(g24595), .A1(g23502), .A2(g23489) );
  AND2_X1 AND2_2608( .ZN(g24596), .A1(g771), .A2(g23887) );
  AND2_X1 AND2_2609( .ZN(g24603), .A1(g23518), .A2(g23505) );
  AND2_X1 AND2_2610( .ZN(g24604), .A1(g1457), .A2(g23908) );
  AND2_X1 AND2_2611( .ZN(g24610), .A1(g23533), .A2(g23521) );
  AND2_X1 AND2_2612( .ZN(g24611), .A1(g2151), .A2(g23940) );
  AND2_X1 AND2_2613( .ZN(g24644), .A1(g17203), .A2(g24115) );
  AND2_X1 AND2_2614( .ZN(g24664), .A1(g17208), .A2(g24134) );
  AND2_X1 AND2_2615( .ZN(g24676), .A1(g13568), .A2(g24115) );
  AND2_X1 AND2_2616( .ZN(g24683), .A1(g17214), .A2(g24153) );
  AND2_X1 AND2_2617( .ZN(g24695), .A1(g13576), .A2(g24134) );
  AND2_X1 AND2_2618( .ZN(g24700), .A1(g17217), .A2(g24168) );
  AND2_X1 AND2_2619( .ZN(g24712), .A1(g13585), .A2(g24153) );
  AND2_X1 AND2_2620( .ZN(g24723), .A1(g13605), .A2(g24168) );
  AND2_X1 AND2_2621( .ZN(g24745), .A1(g15454), .A2(g24096) );
  AND2_X1 AND2_2622( .ZN(g24746), .A1(g15454), .A2(g24098) );
  AND2_X1 AND2_2623( .ZN(g24747), .A1(g9427), .A2(g24099) );
  AND2_X1 AND2_2624( .ZN(g24748), .A1(g672), .A2(g24101) );
  AND2_X1 AND2_2625( .ZN(g24749), .A1(g15540), .A2(g24102) );
  AND2_X1 AND2_2626( .ZN(g24750), .A1(g15454), .A2(g24104) );
  AND2_X1 AND2_2627( .ZN(g24751), .A1(g9427), .A2(g24105) );
  AND2_X1 AND2_2628( .ZN(g24752), .A1(g9507), .A2(g24106) );
  AND2_X1 AND2_2629( .ZN(g24754), .A1(g15540), .A2(g24107) );
  AND2_X1 AND2_2630( .ZN(g24755), .A1(g9569), .A2(g24108) );
  AND2_X1 AND2_2631( .ZN(g24757), .A1(g1358), .A2(g24110) );
  AND2_X1 AND2_2632( .ZN(g24758), .A1(g15618), .A2(g24111) );
  AND2_X1 AND2_2633( .ZN(g24759), .A1(g21825), .A2(g23885) );
  AND2_X1 AND2_2634( .ZN(g24760), .A1(g9427), .A2(g24112) );
  AND2_X1 AND2_2635( .ZN(g24761), .A1(g9507), .A2(g24113) );
  AND2_X1 AND2_2636( .ZN(g24762), .A1(g12876), .A2(g24114) );
  AND2_X1 AND2_2637( .ZN(g24767), .A1(g15540), .A2(g24121) );
  AND2_X1 AND2_2638( .ZN(g24768), .A1(g9569), .A2(g24122) );
  AND2_X1 AND2_2639( .ZN(g24769), .A1(g9649), .A2(g24123) );
  AND2_X1 AND2_2640( .ZN(g24772), .A1(g15618), .A2(g24124) );
  AND2_X1 AND2_2641( .ZN(g24773), .A1(g9711), .A2(g24125) );
  AND2_X1 AND2_2642( .ZN(g24774), .A1(g2052), .A2(g24127) );
  AND2_X1 AND2_2643( .ZN(g24775), .A1(g15694), .A2(g24128) );
  AND2_X1 AND2_2644( .ZN(g24776), .A1(g9507), .A2(g24129) );
  AND2_X1 AND2_2645( .ZN(g24777), .A1(g12876), .A2(g24130) );
  AND2_X1 AND2_2646( .ZN(g24779), .A1(g9569), .A2(g24131) );
  AND2_X1 AND2_2647( .ZN(g24780), .A1(g9649), .A2(g24132) );
  AND2_X1 AND2_2648( .ZN(g24781), .A1(g12916), .A2(g24133) );
  AND2_X1 AND2_2649( .ZN(g24788), .A1(g15618), .A2(g24140) );
  AND2_X1 AND2_2650( .ZN(g24789), .A1(g9711), .A2(g24141) );
  AND2_X1 AND2_2651( .ZN(g24790), .A1(g9795), .A2(g24142) );
  AND2_X1 AND2_2652( .ZN(g24792), .A1(g15694), .A2(g24143) );
  AND2_X1 AND2_2653( .ZN(g24793), .A1(g9857), .A2(g24144) );
  AND2_X1 AND2_2654( .ZN(g24794), .A1(g2746), .A2(g24146) );
  AND2_X1 AND2_2655( .ZN(g24795), .A1(g12017), .A2(g24232) );
  AND2_X1 AND2_2656( .ZN(g24796), .A1(g12876), .A2(g24147) );
  AND2_X1 AND2_2657( .ZN(g24798), .A1(g9649), .A2(g24148) );
  AND2_X1 AND2_2658( .ZN(g24799), .A1(g12916), .A2(g24149) );
  AND2_X1 AND2_2659( .ZN(g24802), .A1(g9711), .A2(g24150) );
  AND2_X1 AND2_2660( .ZN(g24803), .A1(g9795), .A2(g24151) );
  AND2_X1 AND2_2661( .ZN(g24804), .A1(g12945), .A2(g24152) );
  AND2_X1 AND2_2662( .ZN(g24809), .A1(g15694), .A2(g24159) );
  AND2_X1 AND2_2663( .ZN(g24810), .A1(g9857), .A2(g24160) );
  AND2_X1 AND2_2664( .ZN(g24811), .A1(g9941), .A2(g24161) );
  AND2_X1 AND2_2665( .ZN(g24813), .A1(g21825), .A2(g23905) );
  AND2_X1 AND2_2666( .ZN(g24818), .A1(g12916), .A2(g24162) );
  AND2_X1 AND2_2667( .ZN(g24821), .A1(g9795), .A2(g24163) );
  AND2_X1 AND2_2668( .ZN(g24822), .A1(g12945), .A2(g24164) );
  AND2_X1 AND2_2669( .ZN(g24824), .A1(g9857), .A2(g24165) );
  AND2_X1 AND2_2670( .ZN(g24825), .A1(g9941), .A2(g24166) );
  AND2_X1 AND2_2671( .ZN(g24826), .A1(g12974), .A2(g24167) );
  AND2_X1 AND2_2672( .ZN(g24831), .A1(g24100), .A2(g20401) );
  AND2_X1 AND2_2673( .ZN(g24838), .A1(g12945), .A2(g24175) );
  AND2_X1 AND2_2674( .ZN(g24840), .A1(g9941), .A2(g24176) );
  AND2_X1 AND2_2675( .ZN(g24841), .A1(g12974), .A2(g24177) );
  AND2_X1 AND2_2676( .ZN(g24843), .A1(g21825), .A2(g23918) );
  AND2_X1 AND2_2677( .ZN(g24846), .A1(g24109), .A2(g20426) );
  AND2_X1 AND2_2678( .ZN(g24853), .A1(g12974), .A2(g24180) );
  AND2_X1 AND2_2679( .ZN(g24855), .A1(g18174), .A2(g23731) );
  AND2_X1 AND2_2680( .ZN(g24858), .A1(g24047), .A2(g18873) );
  AND2_X1 AND2_2681( .ZN(g24861), .A1(g24126), .A2(g20448) );
  AND2_X1 AND2_2682( .ZN(g24867), .A1(g666), .A2(g23779) );
  AND2_X1 AND2_2683( .ZN(g24869), .A1(g24047), .A2(g18894) );
  AND2_X1 AND2_2684( .ZN(g24870), .A1(g18281), .A2(g23786) );
  AND2_X1 AND2_2685( .ZN(g24874), .A1(g24060), .A2(g18899) );
  AND2_X2 AND2_2686( .ZN(g24876), .A1(g24145), .A2(g20467) );
  AND2_X2 AND2_2687( .ZN(g24878), .A1(g19830), .A2(g24210) );
  AND2_X2 AND2_2688( .ZN(g24881), .A1(g24047), .A2(g18912) );
  AND2_X1 AND2_2689( .ZN(g24882), .A1(g1352), .A2(g23832) );
  AND2_X1 AND2_2690( .ZN(g24884), .A1(g24060), .A2(g18917) );
  AND2_X1 AND2_2691( .ZN(g24885), .A1(g18374), .A2(g23839) );
  AND2_X1 AND2_2692( .ZN(g24888), .A1(g24073), .A2(g18922) );
  AND2_X1 AND2_2693( .ZN(g24898), .A1(g24060), .A2(g18931) );
  AND2_X1 AND2_2694( .ZN(g24899), .A1(g2046), .A2(g23867) );
  AND2_X1 AND2_2695( .ZN(g24901), .A1(g24073), .A2(g18936) );
  AND2_X1 AND2_2696( .ZN(g24902), .A1(g18469), .A2(g23874) );
  AND2_X1 AND2_2697( .ZN(g24905), .A1(g24084), .A2(g18941) );
  AND2_X1 AND2_2698( .ZN(g24906), .A1(g18886), .A2(g23879) );
  AND2_X1 AND2_2699( .ZN(g24907), .A1(g7466), .A2(g24220) );
  AND2_X1 AND2_2700( .ZN(g24908), .A1(g7342), .A2(g23882) );
  AND2_X1 AND2_2701( .ZN(g24921), .A1(g24073), .A2(g18951) );
  AND2_X1 AND2_2702( .ZN(g24922), .A1(g2740), .A2(g23901) );
  AND2_X1 AND2_2703( .ZN(g24924), .A1(g24084), .A2(g18956) );
  AND2_X1 AND2_2704( .ZN(g24938), .A1(g24084), .A2(g18967) );
  AND2_X1 AND2_2705( .ZN(g24964), .A1(g7595), .A2(g24251) );
  AND2_X1 AND2_2706( .ZN(g24974), .A1(g7600), .A2(g24030) );
  AND2_X1 AND2_2707( .ZN(g25086), .A1(g23444), .A2(g10880) );
  AND2_X1 AND2_2708( .ZN(g25102), .A1(g23444), .A2(g10915) );
  AND2_X1 AND2_2709( .ZN(g25117), .A1(g23444), .A2(g10974) );
  AND3_X1 AND3_245( .ZN(g25128), .A1(g17051), .A2(g24115), .A3(g13614) );
  AND2_X1 AND2_2710( .ZN(g25178), .A1(g24623), .A2(g20634) );
  AND2_X1 AND2_2711( .ZN(g25181), .A1(g24636), .A2(g20673) );
  AND2_X1 AND2_2712( .ZN(g25182), .A1(g24681), .A2(g20676) );
  AND2_X1 AND2_2713( .ZN(g25184), .A1(g24694), .A2(g20735) );
  AND2_X1 AND2_2714( .ZN(g25187), .A1(g24633), .A2(g16608) );
  AND2_X1 AND2_2715( .ZN(g25188), .A1(g24652), .A2(g20763) );
  AND2_X1 AND2_2716( .ZN(g25192), .A1(g24711), .A2(g20790) );
  AND2_X1 AND2_2717( .ZN(g25193), .A1(g24653), .A2(g16626) );
  AND2_X1 AND2_2718( .ZN(g25196), .A1(g24672), .A2(g16640) );
  AND2_X1 AND2_2719( .ZN(g25198), .A1(g24691), .A2(g16651) );
  AND2_X1 AND2_2720( .ZN(g25269), .A1(g24648), .A2(g8700) );
  AND2_X1 AND2_2721( .ZN(g25277), .A1(g24648), .A2(g8714) );
  AND2_X1 AND2_2722( .ZN(g25278), .A1(g24668), .A2(g8719) );
  AND2_X1 AND2_2723( .ZN(g25281), .A1(g5606), .A2(g24815) );
  AND2_X1 AND2_2724( .ZN(g25282), .A1(g24648), .A2(g8748) );
  AND2_X1 AND2_2725( .ZN(g25286), .A1(g24668), .A2(g8752) );
  AND2_X1 AND2_2726( .ZN(g25287), .A1(g24687), .A2(g8757) );
  AND2_X1 AND2_2727( .ZN(g25289), .A1(g5631), .A2(g24834) );
  AND2_X1 AND2_2728( .ZN(g25290), .A1(g24668), .A2(g8771) );
  AND2_X1 AND2_2729( .ZN(g25294), .A1(g24687), .A2(g8775) );
  AND2_X1 AND2_2730( .ZN(g25295), .A1(g24704), .A2(g8780) );
  AND2_X1 AND2_2731( .ZN(g25299), .A1(g5659), .A2(g24850) );
  AND2_X1 AND2_2732( .ZN(g25300), .A1(g24687), .A2(g8794) );
  AND2_X1 AND2_2733( .ZN(g25304), .A1(g24704), .A2(g8798) );
  AND2_X1 AND2_2734( .ZN(g25309), .A1(g5697), .A2(g24864) );
  AND2_X1 AND2_2735( .ZN(g25310), .A1(g24704), .A2(g8813) );
  AND3_X1 AND3_246( .ZN(g25318), .A1(g24682), .A2(g19358), .A3(g19335) );
  AND2_X1 AND2_2736( .ZN(g25321), .A1(g25075), .A2(g9669) );
  AND2_X1 AND2_2737( .ZN(g25328), .A1(g24644), .A2(g17892) );
  AND2_X1 AND2_2738( .ZN(g25334), .A1(g24644), .A2(g17984) );
  AND2_X1 AND2_2739( .ZN(g25337), .A1(g24664), .A2(g18003) );
  AND2_X1 AND2_2740( .ZN(g25342), .A1(g5851), .A2(g24600) );
  AND2_X1 AND2_2741( .ZN(g25346), .A1(g24644), .A2(g18084) );
  AND2_X1 AND2_2742( .ZN(g25348), .A1(g24664), .A2(g18101) );
  AND2_X1 AND2_2743( .ZN(g25351), .A1(g24683), .A2(g18120) );
  AND2_X1 AND2_2744( .ZN(g25356), .A1(g5898), .A2(g24607) );
  AND2_X1 AND2_2745( .ZN(g25360), .A1(g24664), .A2(g18200) );
  AND2_X1 AND2_2746( .ZN(g25362), .A1(g24683), .A2(g18217) );
  AND2_X1 AND2_2747( .ZN(g25365), .A1(g24700), .A2(g18236) );
  AND2_X1 AND2_2748( .ZN(g25371), .A1(g5937), .A2(g24619) );
  AND2_X1 AND2_2749( .ZN(g25375), .A1(g24683), .A2(g18307) );
  AND2_X1 AND2_2750( .ZN(g25377), .A1(g24700), .A2(g18324) );
  AND2_X1 AND2_2751( .ZN(g25388), .A1(g5971), .A2(g24630) );
  AND2_X1 AND2_2752( .ZN(g25392), .A1(g24700), .A2(g18400) );
  AND2_X1 AND2_2753( .ZN(g25453), .A1(g6142), .A2(g24763) );
  AND2_X1 AND2_2754( .ZN(g25457), .A1(g6163), .A2(g24784) );
  AND2_X1 AND2_2755( .ZN(g25461), .A1(g6190), .A2(g24805) );
  AND2_X1 AND2_2756( .ZN(g25466), .A1(g6222), .A2(g24827) );
  AND2_X1 AND2_2757( .ZN(g25470), .A1(g24479), .A2(g20400) );
  AND2_X1 AND2_2758( .ZN(g25475), .A1(g14148), .A2(g25087) );
  AND2_X1 AND2_2759( .ZN(g25482), .A1(g24480), .A2(g17567) );
  AND2_X1 AND2_2760( .ZN(g25483), .A1(g24481), .A2(g20421) );
  AND2_X1 AND2_2761( .ZN(g25487), .A1(g24485), .A2(g20425) );
  AND2_X1 AND2_2762( .ZN(g25505), .A1(g6707), .A2(g25094) );
  AND2_X1 AND2_2763( .ZN(g25506), .A1(g14263), .A2(g25095) );
  AND2_X1 AND2_2764( .ZN(g25513), .A1(g24487), .A2(g17664) );
  AND2_X1 AND2_2765( .ZN(g25514), .A1(g24488), .A2(g20443) );
  AND2_X1 AND2_2766( .ZN(g25518), .A1(g24489), .A2(g20447) );
  AND2_X1 AND2_2767( .ZN(g25552), .A1(g7009), .A2(g25104) );
  AND2_X1 AND2_2768( .ZN(g25553), .A1(g14385), .A2(g25105) );
  AND2_X1 AND2_2769( .ZN(g25560), .A1(g24494), .A2(g17764) );
  AND2_X1 AND2_2770( .ZN(g25561), .A1(g24495), .A2(g20462) );
  AND2_X1 AND2_2771( .ZN(g25565), .A1(g24496), .A2(g20466) );
  AND2_X1 AND2_2772( .ZN(g25618), .A1(g7259), .A2(g25110) );
  AND2_X1 AND2_2773( .ZN(g25619), .A1(g14497), .A2(g25111) );
  AND2_X1 AND2_2774( .ZN(g25626), .A1(g24504), .A2(g17865) );
  AND2_X1 AND2_2775( .ZN(g25627), .A1(g24505), .A2(g20477) );
  AND2_X1 AND2_2776( .ZN(g25628), .A1(g21008), .A2(g25115) );
  AND2_X1 AND2_2777( .ZN(g25629), .A1(g3024), .A2(g25116) );
  AND2_X1 AND2_2778( .ZN(g25697), .A1(g7455), .A2(g25120) );
  AND2_X1 AND2_2779( .ZN(g25881), .A1(g2908), .A2(g25126) );
  AND2_X1 AND2_2780( .ZN(g25951), .A1(g24800), .A2(g13670) );
  AND2_X1 AND2_2781( .ZN(g25953), .A1(g24783), .A2(g13699) );
  AND2_X1 AND2_2782( .ZN(g25957), .A1(g24782), .A2(g11869) );
  AND2_X1 AND2_2783( .ZN(g25961), .A1(g24770), .A2(g11901) );
  AND2_X1 AND2_2784( .ZN(g25963), .A1(g24756), .A2(g11944) );
  AND2_X1 AND2_2785( .ZN(g25968), .A1(g24871), .A2(g11986) );
  AND2_X1 AND2_2786( .ZN(g25972), .A1(g24859), .A2(g12042) );
  AND2_X1 AND2_2787( .ZN(g25973), .A1(g24847), .A2(g13838) );
  AND2_X1 AND2_2788( .ZN(g25975), .A1(g24606), .A2(g21917) );
  AND2_X1 AND2_2789( .ZN(g25977), .A1(g24845), .A2(g12089) );
  AND2_X1 AND2_2790( .ZN(g25978), .A1(g24836), .A2(g13850) );
  AND2_X1 AND2_2791( .ZN(g25980), .A1(g24663), .A2(g21928) );
  AND2_X1 AND2_2792( .ZN(g25981), .A1(g24819), .A2(g13858) );
  AND2_X1 AND2_2793( .ZN(g26023), .A1(g25422), .A2(g24912) );
  AND2_X1 AND2_2794( .ZN(g26024), .A1(g25301), .A2(g21102) );
  AND2_X1 AND2_2795( .ZN(g26026), .A1(g25431), .A2(g24929) );
  AND2_X1 AND2_2796( .ZN(g26027), .A1(g25418), .A2(g22271) );
  AND2_X1 AND2_2797( .ZN(g26028), .A1(g25438), .A2(g24941) );
  AND2_X1 AND2_2798( .ZN(g26029), .A1(g25445), .A2(g24952) );
  AND2_X1 AND2_2799( .ZN(g26030), .A1(g25429), .A2(g22304) );
  AND2_X1 AND2_2800( .ZN(g26032), .A1(g25379), .A2(g19415) );
  AND2_X1 AND2_2801( .ZN(g26033), .A1(g25395), .A2(g19452) );
  AND2_X1 AND2_2802( .ZN(g26034), .A1(g25405), .A2(g19479) );
  AND2_X1 AND2_2803( .ZN(g26035), .A1(g25523), .A2(g19483) );
  AND2_X1 AND2_2804( .ZN(g26036), .A1(g25413), .A2(g19502) );
  AND2_X1 AND2_2805( .ZN(g26038), .A1(g25589), .A2(g19504) );
  AND2_X1 AND2_2806( .ZN(g26039), .A1(g25668), .A2(g19523) );
  AND2_X1 AND2_2807( .ZN(g26040), .A1(g25745), .A2(g19533) );
  AND2_X1 AND2_2808( .ZN(g26051), .A1(g70), .A2(g25296) );
  AND2_X1 AND2_2809( .ZN(g26052), .A1(g25941), .A2(g21087) );
  AND2_X1 AND2_2810( .ZN(g26053), .A1(g758), .A2(g25306) );
  AND2_X1 AND2_2811( .ZN(g26054), .A1(g25944), .A2(g21099) );
  AND2_X1 AND2_2812( .ZN(g26060), .A1(g25943), .A2(g21108) );
  AND2_X1 AND2_2813( .ZN(g26061), .A1(g1444), .A2(g25315) );
  AND2_X1 AND2_2814( .ZN(g26062), .A1(g25947), .A2(g21113) );
  AND2_X1 AND2_2815( .ZN(g26067), .A1(g25946), .A2(g21125) );
  AND2_X1 AND2_2816( .ZN(g26068), .A1(g2138), .A2(g25324) );
  AND2_X1 AND2_2817( .ZN(g26069), .A1(g25949), .A2(g21130) );
  AND2_X1 AND2_2818( .ZN(g26074), .A1(g25948), .A2(g21144) );
  AND2_X1 AND2_2819( .ZN(g26075), .A1(g74), .A2(g25698) );
  AND2_X1 AND2_2820( .ZN(g26080), .A1(g25950), .A2(g21164) );
  AND2_X1 AND2_2821( .ZN(g26082), .A1(g762), .A2(g25771) );
  AND2_X1 AND2_2822( .ZN(g26085), .A1(g1448), .A2(g25825) );
  AND2_X1 AND2_2823( .ZN(g26091), .A1(g2142), .A2(g25860) );
  AND2_X1 AND2_2824( .ZN(g26157), .A1(g21825), .A2(g25630) );
  AND2_X1 AND2_2825( .ZN(g26158), .A1(g679), .A2(g25937) );
  AND2_X1 AND2_2826( .ZN(g26163), .A1(g1365), .A2(g25939) );
  AND2_X1 AND2_2827( .ZN(g26166), .A1(g686), .A2(g25454) );
  AND2_X1 AND2_2828( .ZN(g26171), .A1(g2059), .A2(g25942) );
  AND2_X1 AND2_2829( .ZN(g26186), .A1(g1372), .A2(g25458) );
  AND2_X1 AND2_2830( .ZN(g26188), .A1(g2753), .A2(g25945) );
  AND2_X1 AND2_2831( .ZN(g26207), .A1(g2066), .A2(g25463) );
  AND2_X1 AND2_2832( .ZN(g26212), .A1(g4217), .A2(g25467) );
  AND2_X1 AND2_2833( .ZN(g26213), .A1(g25895), .A2(g9306) );
  AND2_X1 AND2_2834( .ZN(g26231), .A1(g2760), .A2(g25472) );
  AND2_X1 AND2_2835( .ZN(g26233), .A1(g4340), .A2(g25476) );
  AND2_X1 AND2_2836( .ZN(g26234), .A1(g4343), .A2(g25479) );
  AND2_X1 AND2_2837( .ZN(g26235), .A1(g25895), .A2(g9368) );
  AND2_X1 AND2_2838( .ZN(g26236), .A1(g25899), .A2(g9371) );
  AND2_X1 AND2_2839( .ZN(g26243), .A1(g4372), .A2(g25484) );
  AND2_X1 AND2_2840( .ZN(g26244), .A1(g25903), .A2(g9387) );
  AND2_X1 AND2_2841( .ZN(g26257), .A1(g4465), .A2(g25493) );
  AND2_X1 AND2_2842( .ZN(g26258), .A1(g4468), .A2(g25496) );
  AND2_X1 AND2_2843( .ZN(g26259), .A1(g4471), .A2(g25499) );
  AND2_X1 AND2_2844( .ZN(g26260), .A1(g25254), .A2(g17649) );
  AND2_X1 AND2_2845( .ZN(g26261), .A1(g25895), .A2(g9443) );
  AND2_X1 AND2_2846( .ZN(g26262), .A1(g25899), .A2(g9446) );
  AND2_X1 AND2_2847( .ZN(g26263), .A1(g4476), .A2(g25502) );
  AND2_X1 AND2_2848( .ZN(g26268), .A1(g4509), .A2(g25507) );
  AND2_X1 AND2_2849( .ZN(g26269), .A1(g4512), .A2(g25510) );
  AND2_X1 AND2_2850( .ZN(g26270), .A1(g25903), .A2(g9465) );
  AND2_X1 AND2_2851( .ZN(g26271), .A1(g25907), .A2(g9468) );
  AND2_X1 AND2_2852( .ZN(g26278), .A1(g4541), .A2(g25515) );
  AND2_X1 AND2_2853( .ZN(g26279), .A1(g25911), .A2(g9484) );
  AND2_X1 AND2_2854( .ZN(g26288), .A1(g4592), .A2(g25524) );
  AND2_X1 AND2_2855( .ZN(g26289), .A1(g4595), .A2(g25527) );
  AND2_X1 AND2_2856( .ZN(g26290), .A1(g4598), .A2(g25530) );
  AND2_X2 AND2_2857( .ZN(g26291), .A1(g25899), .A2(g9524) );
  AND2_X2 AND2_2858( .ZN(g26292), .A1(g4603), .A2(g25533) );
  AND2_X1 AND2_2859( .ZN(g26293), .A1(g4606), .A2(g25536) );
  AND2_X1 AND2_2860( .ZN(g26298), .A1(g4641), .A2(g25540) );
  AND2_X1 AND2_2861( .ZN(g26299), .A1(g4644), .A2(g25543) );
  AND2_X1 AND2_2862( .ZN(g26300), .A1(g4647), .A2(g25546) );
  AND2_X1 AND2_2863( .ZN(g26301), .A1(g25258), .A2(g17749) );
  AND2_X1 AND2_2864( .ZN(g26302), .A1(g25903), .A2(g9585) );
  AND2_X1 AND2_2865( .ZN(g26303), .A1(g25907), .A2(g9588) );
  AND2_X1 AND2_2866( .ZN(g26307), .A1(g4652), .A2(g25549) );
  AND2_X1 AND2_2867( .ZN(g26309), .A1(g4685), .A2(g25554) );
  AND2_X1 AND2_2868( .ZN(g26310), .A1(g4688), .A2(g25557) );
  AND2_X1 AND2_2869( .ZN(g26311), .A1(g25911), .A2(g9607) );
  AND2_X1 AND2_2870( .ZN(g26312), .A1(g25915), .A2(g9610) );
  AND2_X1 AND2_2871( .ZN(g26316), .A1(g4717), .A2(g25562) );
  AND2_X1 AND2_2872( .ZN(g26317), .A1(g25919), .A2(g9626) );
  AND2_X1 AND2_2873( .ZN(g26318), .A1(g4737), .A2(g25573) );
  AND2_X1 AND2_2874( .ZN(g26319), .A1(g4740), .A2(g25576) );
  AND2_X1 AND2_2875( .ZN(g26324), .A1(g4743), .A2(g25579) );
  AND2_X1 AND2_2876( .ZN(g26325), .A1(g4746), .A2(g25582) );
  AND2_X1 AND2_2877( .ZN(g26326), .A1(g4749), .A2(g25585) );
  AND2_X1 AND2_2878( .ZN(g26332), .A1(g4769), .A2(g25590) );
  AND2_X1 AND2_2879( .ZN(g26333), .A1(g4772), .A2(g25593) );
  AND2_X1 AND2_2880( .ZN(g26334), .A1(g4775), .A2(g25596) );
  AND2_X1 AND2_2881( .ZN(g26335), .A1(g25907), .A2(g9666) );
  AND2_X1 AND2_2882( .ZN(g26339), .A1(g4780), .A2(g25599) );
  AND2_X1 AND2_2883( .ZN(g26340), .A1(g4783), .A2(g25602) );
  AND2_X1 AND2_2884( .ZN(g26342), .A1(g4818), .A2(g25606) );
  AND2_X1 AND2_2885( .ZN(g26343), .A1(g4821), .A2(g25609) );
  AND2_X1 AND2_2886( .ZN(g26344), .A1(g4824), .A2(g25612) );
  AND2_X1 AND2_2887( .ZN(g26345), .A1(g25261), .A2(g17850) );
  AND2_X1 AND2_2888( .ZN(g26346), .A1(g25911), .A2(g9727) );
  AND2_X1 AND2_2889( .ZN(g26347), .A1(g25915), .A2(g9730) );
  AND2_X1 AND2_2890( .ZN(g26348), .A1(g4829), .A2(g25615) );
  AND2_X1 AND2_2891( .ZN(g26350), .A1(g4862), .A2(g25620) );
  AND2_X1 AND2_2892( .ZN(g26351), .A1(g4865), .A2(g25623) );
  AND2_X1 AND2_2893( .ZN(g26352), .A1(g25919), .A2(g9749) );
  AND2_X1 AND2_2894( .ZN(g26353), .A1(g25923), .A2(g9752) );
  AND2_X1 AND2_2895( .ZN(g26357), .A1(g4882), .A2(g25634) );
  AND2_X1 AND2_2896( .ZN(g26361), .A1(g4888), .A2(g25637) );
  AND2_X1 AND2_2897( .ZN(g26362), .A1(g4891), .A2(g25640) );
  AND2_X1 AND2_2898( .ZN(g26363), .A1(g4894), .A2(g25643) );
  AND2_X1 AND2_2899( .ZN(g26365), .A1(g4913), .A2(g25652) );
  AND2_X1 AND2_2900( .ZN(g26366), .A1(g4916), .A2(g25655) );
  AND2_X1 AND2_2901( .ZN(g26371), .A1(g4919), .A2(g25658) );
  AND2_X1 AND2_2902( .ZN(g26372), .A1(g4922), .A2(g25661) );
  AND2_X1 AND2_2903( .ZN(g26373), .A1(g4925), .A2(g25664) );
  AND2_X1 AND2_2904( .ZN(g26379), .A1(g4945), .A2(g25669) );
  AND2_X1 AND2_2905( .ZN(g26380), .A1(g4948), .A2(g25672) );
  AND2_X1 AND2_2906( .ZN(g26381), .A1(g4951), .A2(g25675) );
  AND2_X1 AND2_2907( .ZN(g26382), .A1(g25915), .A2(g9812) );
  AND2_X1 AND2_2908( .ZN(g26383), .A1(g4956), .A2(g25678) );
  AND2_X1 AND2_2909( .ZN(g26384), .A1(g4959), .A2(g25681) );
  AND2_X1 AND2_2910( .ZN(g26386), .A1(g4994), .A2(g25685) );
  AND2_X1 AND2_2911( .ZN(g26387), .A1(g4997), .A2(g25688) );
  AND2_X1 AND2_2912( .ZN(g26388), .A1(g5000), .A2(g25691) );
  AND2_X1 AND2_2913( .ZN(g26389), .A1(g25264), .A2(g17962) );
  AND2_X1 AND2_2914( .ZN(g26390), .A1(g25919), .A2(g9873) );
  AND2_X1 AND2_2915( .ZN(g26391), .A1(g25923), .A2(g9876) );
  AND2_X1 AND2_2916( .ZN(g26392), .A1(g5005), .A2(g25694) );
  AND2_X1 AND2_2917( .ZN(g26396), .A1(g5027), .A2(g25700) );
  AND2_X1 AND2_2918( .ZN(g26397), .A1(g5030), .A2(g25703) );
  AND2_X1 AND2_2919( .ZN(g26400), .A1(g5041), .A2(g25711) );
  AND2_X1 AND2_2920( .ZN(g26404), .A1(g5047), .A2(g25714) );
  AND2_X1 AND2_2921( .ZN(g26405), .A1(g5050), .A2(g25717) );
  AND2_X1 AND2_2922( .ZN(g26406), .A1(g5053), .A2(g25720) );
  AND2_X1 AND2_2923( .ZN(g26408), .A1(g5072), .A2(g25729) );
  AND2_X1 AND2_2924( .ZN(g26409), .A1(g5075), .A2(g25732) );
  AND2_X1 AND2_2925( .ZN(g26414), .A1(g5078), .A2(g25735) );
  AND2_X1 AND2_2926( .ZN(g26415), .A1(g5081), .A2(g25738) );
  AND2_X1 AND2_2927( .ZN(g26416), .A1(g5084), .A2(g25741) );
  AND2_X1 AND2_2928( .ZN(g26422), .A1(g5104), .A2(g25746) );
  AND2_X1 AND2_2929( .ZN(g26423), .A1(g5107), .A2(g25749) );
  AND2_X1 AND2_2930( .ZN(g26424), .A1(g5110), .A2(g25752) );
  AND2_X1 AND2_2931( .ZN(g26425), .A1(g25923), .A2(g9958) );
  AND2_X1 AND2_2932( .ZN(g26426), .A1(g5115), .A2(g25755) );
  AND2_X1 AND2_2933( .ZN(g26427), .A1(g5118), .A2(g25758) );
  AND2_X1 AND2_2934( .ZN(g26432), .A1(g5145), .A2(g25767) );
  AND2_X1 AND2_2935( .ZN(g26437), .A1(g5156), .A2(g25773) );
  AND2_X1 AND2_2936( .ZN(g26438), .A1(g5159), .A2(g25776) );
  AND2_X1 AND2_2937( .ZN(g26441), .A1(g5170), .A2(g25784) );
  AND2_X1 AND2_2938( .ZN(g26445), .A1(g5176), .A2(g25787) );
  AND2_X1 AND2_2939( .ZN(g26446), .A1(g5179), .A2(g25790) );
  AND2_X1 AND2_2940( .ZN(g26447), .A1(g5182), .A2(g25793) );
  AND2_X1 AND2_2941( .ZN(g26449), .A1(g5201), .A2(g25802) );
  AND2_X1 AND2_2942( .ZN(g26450), .A1(g5204), .A2(g25805) );
  AND2_X1 AND2_2943( .ZN(g26455), .A1(g5207), .A2(g25808) );
  AND2_X1 AND2_2944( .ZN(g26456), .A1(g5210), .A2(g25811) );
  AND2_X1 AND2_2945( .ZN(g26457), .A1(g5213), .A2(g25814) );
  AND2_X1 AND2_2946( .ZN(g26464), .A1(g5238), .A2(g25821) );
  AND2_X1 AND2_2947( .ZN(g26469), .A1(g5249), .A2(g25827) );
  AND2_X1 AND2_2948( .ZN(g26470), .A1(g5252), .A2(g25830) );
  AND2_X1 AND2_2949( .ZN(g26473), .A1(g5263), .A2(g25838) );
  AND2_X1 AND2_2950( .ZN(g26477), .A1(g5269), .A2(g25841) );
  AND2_X1 AND2_2951( .ZN(g26478), .A1(g5272), .A2(g25844) );
  AND2_X1 AND2_2952( .ZN(g26479), .A1(g5275), .A2(g25847) );
  AND2_X1 AND2_2953( .ZN(g26488), .A1(g5301), .A2(g25856) );
  AND2_X1 AND2_2954( .ZN(g26493), .A1(g5312), .A2(g25862) );
  AND2_X1 AND2_2955( .ZN(g26494), .A1(g5315), .A2(g25865) );
  AND2_X1 AND2_2956( .ZN(g26504), .A1(g5338), .A2(g25877) );
  AND2_X1 AND2_2957( .ZN(g26663), .A1(g25274), .A2(g21066) );
  AND2_X1 AND2_2958( .ZN(g26668), .A1(g25283), .A2(g21076) );
  AND2_X1 AND2_2959( .ZN(g26673), .A1(g12431), .A2(g25318) );
  AND2_X1 AND2_2960( .ZN(g26674), .A1(g25291), .A2(g21090) );
  AND2_X1 AND2_2961( .ZN(g26754), .A1(g14657), .A2(g26508) );
  AND2_X1 AND2_2962( .ZN(g26755), .A1(g26083), .A2(g22239) );
  AND2_X1 AND2_2963( .ZN(g26756), .A1(g26113), .A2(g22240) );
  AND3_X1 AND3_247( .ZN(g26758), .A1(g16614), .A2(g26521), .A3(g13637) );
  AND2_X1 AND2_2964( .ZN(g26759), .A1(g26356), .A2(g19251) );
  AND2_X1 AND2_2965( .ZN(g26760), .A1(g26137), .A2(g22256) );
  AND2_X1 AND2_2966( .ZN(g26761), .A1(g26154), .A2(g22257) );
  AND2_X1 AND2_2967( .ZN(g26763), .A1(g14691), .A2(g26516) );
  AND3_X1 AND3_248( .ZN(g26764), .A1(g16632), .A2(g26525), .A3(g13649) );
  AND2_X1 AND2_2968( .ZN(g26765), .A1(g26399), .A2(g19265) );
  AND2_X1 AND2_2969( .ZN(g26766), .A1(g14725), .A2(g26521) );
  AND2_X2 AND2_2970( .ZN(g26767), .A1(g26087), .A2(g22287) );
  AND2_X2 AND2_2971( .ZN(g26768), .A1(g26440), .A2(g19280) );
  AND2_X1 AND2_2972( .ZN(g26769), .A1(g14753), .A2(g26525) );
  AND2_X1 AND2_2973( .ZN(g26770), .A1(g26059), .A2(g19287) );
  AND3_X1 AND3_249( .ZN(g26771), .A1(g24912), .A2(g26508), .A3(g13614) );
  AND2_X1 AND2_2974( .ZN(g26773), .A1(g26145), .A2(g22303) );
  AND2_X1 AND2_2975( .ZN(g26774), .A1(g26472), .A2(g19299) );
  AND2_X1 AND2_2976( .ZN(g26775), .A1(g26099), .A2(g22318) );
  AND2_X1 AND2_2977( .ZN(g26777), .A1(g26066), .A2(g19305) );
  AND3_X1 AND3_250( .ZN(g26778), .A1(g24929), .A2(g26516), .A3(g13626) );
  AND2_X1 AND2_2978( .ZN(g26780), .A1(g26119), .A2(g16622) );
  AND2_X1 AND2_2979( .ZN(g26783), .A1(g26073), .A2(g19326) );
  AND3_X1 AND3_251( .ZN(g26784), .A1(g24941), .A2(g26521), .A3(g13637) );
  AND2_X1 AND2_2980( .ZN(g26787), .A1(g26129), .A2(g16636) );
  AND2_X1 AND2_2981( .ZN(g26790), .A1(g26079), .A2(g19353) );
  AND3_X1 AND3_252( .ZN(g26791), .A1(g24952), .A2(g26525), .A3(g13649) );
  AND2_X1 AND2_2982( .ZN(g26794), .A1(g26143), .A2(g16647) );
  AND2_X1 AND2_2983( .ZN(g26797), .A1(g26148), .A2(g16659) );
  AND2_X1 AND2_2984( .ZN(g26829), .A1(g5623), .A2(g26209) );
  AND2_X1 AND2_2985( .ZN(g26833), .A1(g5651), .A2(g26237) );
  AND2_X1 AND2_2986( .ZN(g26842), .A1(g5689), .A2(g26275) );
  AND2_X1 AND2_2987( .ZN(g26845), .A1(g5664), .A2(g26056) );
  AND2_X1 AND2_2988( .ZN(g26851), .A1(g5741), .A2(g26313) );
  AND2_X1 AND2_2989( .ZN(g26853), .A1(g5716), .A2(g26063) );
  AND2_X1 AND2_2990( .ZN(g26860), .A1(g5774), .A2(g26070) );
  AND2_X1 AND2_2991( .ZN(g26866), .A1(g5833), .A2(g26076) );
  AND2_X1 AND2_2992( .ZN(g26955), .A1(g6157), .A2(g26533) );
  AND2_X1 AND2_2993( .ZN(g26958), .A1(g6184), .A2(g26538) );
  AND2_X1 AND2_2994( .ZN(g26961), .A1(g13907), .A2(g26175) );
  AND2_X1 AND2_2995( .ZN(g26962), .A1(g6180), .A2(g26178) );
  AND2_X1 AND2_2996( .ZN(g26963), .A1(g6216), .A2(g26539) );
  AND2_X1 AND2_2997( .ZN(g26965), .A1(g23320), .A2(g26540) );
  AND2_X1 AND2_2998( .ZN(g26966), .A1(g13963), .A2(g26196) );
  AND2_X1 AND2_2999( .ZN(g26967), .A1(g6212), .A2(g26202) );
  AND2_X1 AND2_3000( .ZN(g26968), .A1(g6305), .A2(g26542) );
  AND2_X1 AND2_3001( .ZN(g26969), .A1(g23320), .A2(g26543) );
  AND2_X1 AND2_3002( .ZN(g26970), .A1(g21976), .A2(g26544) );
  AND2_X1 AND2_3003( .ZN(g26971), .A1(g23325), .A2(g26546) );
  AND2_X1 AND2_3004( .ZN(g26972), .A1(g14033), .A2(g26223) );
  AND2_X1 AND2_3005( .ZN(g26973), .A1(g6301), .A2(g26226) );
  AND2_X1 AND2_3006( .ZN(g26977), .A1(g23320), .A2(g26550) );
  AND2_X1 AND2_3007( .ZN(g26978), .A1(g21976), .A2(g26551) );
  AND2_X1 AND2_3008( .ZN(g26979), .A1(g23331), .A2(g26552) );
  AND2_X1 AND2_3009( .ZN(g26980), .A1(g23360), .A2(g26554) );
  AND2_X1 AND2_3010( .ZN(g26981), .A1(g23325), .A2(g26555) );
  AND2_X1 AND2_3011( .ZN(g26982), .A1(g21983), .A2(g26556) );
  AND2_X1 AND2_3012( .ZN(g26984), .A1(g23335), .A2(g26558) );
  AND2_X1 AND2_3013( .ZN(g26985), .A1(g14124), .A2(g26251) );
  AND2_X1 AND2_3014( .ZN(g26986), .A1(g6438), .A2(g26254) );
  AND2_X1 AND2_3015( .ZN(g26993), .A1(g21976), .A2(g26561) );
  AND2_X1 AND2_3016( .ZN(g26994), .A1(g23331), .A2(g26562) );
  AND2_X1 AND2_3017( .ZN(g26995), .A1(g21991), .A2(g26563) );
  AND2_X1 AND2_3018( .ZN(g26996), .A1(g23360), .A2(g26564) );
  AND2_X1 AND2_3019( .ZN(g26997), .A1(g22050), .A2(g26565) );
  AND2_X1 AND2_3020( .ZN(g26998), .A1(g23325), .A2(g26566) );
  AND2_X1 AND2_3021( .ZN(g26999), .A1(g21983), .A2(g26567) );
  AND2_X1 AND2_3022( .ZN(g27000), .A1(g23340), .A2(g26568) );
  AND2_X1 AND2_3023( .ZN(g27001), .A1(g23364), .A2(g26570) );
  AND2_X1 AND2_3024( .ZN(g27002), .A1(g23335), .A2(g26571) );
  AND2_X1 AND2_3025( .ZN(g27003), .A1(g21996), .A2(g26572) );
  AND2_X1 AND2_3026( .ZN(g27004), .A1(g23344), .A2(g26574) );
  AND2_X1 AND2_3027( .ZN(g27005), .A1(g23331), .A2(g26578) );
  AND2_X1 AND2_3028( .ZN(g27006), .A1(g21991), .A2(g26579) );
  AND2_X1 AND2_3029( .ZN(g27007), .A1(g23360), .A2(g26580) );
  AND2_X1 AND2_3030( .ZN(g27008), .A1(g22050), .A2(g26581) );
  AND2_X1 AND2_3031( .ZN(g27009), .A1(g23368), .A2(g26582) );
  AND2_X1 AND2_3032( .ZN(g27016), .A1(g21983), .A2(g26584) );
  AND2_X1 AND2_3033( .ZN(g27017), .A1(g23340), .A2(g26585) );
  AND2_X1 AND2_3034( .ZN(g27018), .A1(g22005), .A2(g26586) );
  AND2_X1 AND2_3035( .ZN(g27019), .A1(g23364), .A2(g26587) );
  AND2_X1 AND2_3036( .ZN(g27020), .A1(g22069), .A2(g26588) );
  AND2_X1 AND2_3037( .ZN(g27021), .A1(g23335), .A2(g26589) );
  AND2_X1 AND2_3038( .ZN(g27022), .A1(g21996), .A2(g26590) );
  AND2_X1 AND2_3039( .ZN(g27023), .A1(g23349), .A2(g26591) );
  AND2_X1 AND2_3040( .ZN(g27024), .A1(g23372), .A2(g26593) );
  AND2_X1 AND2_3041( .ZN(g27025), .A1(g23344), .A2(g26594) );
  AND2_X1 AND2_3042( .ZN(g27026), .A1(g22009), .A2(g26595) );
  AND2_X1 AND2_3043( .ZN(g27027), .A1(g21991), .A2(g26598) );
  AND2_X1 AND2_3044( .ZN(g27028), .A1(g22050), .A2(g26599) );
  AND2_X1 AND2_3045( .ZN(g27029), .A1(g23368), .A2(g26600) );
  AND2_X1 AND2_3046( .ZN(g27030), .A1(g22083), .A2(g26601) );
  AND2_X1 AND2_3047( .ZN(g27031), .A1(g23340), .A2(g26602) );
  AND2_X1 AND2_3048( .ZN(g27032), .A1(g22005), .A2(g26603) );
  AND2_X1 AND2_3049( .ZN(g27033), .A1(g23364), .A2(g26604) );
  AND2_X1 AND2_3050( .ZN(g27034), .A1(g22069), .A2(g26605) );
  AND2_X1 AND2_3051( .ZN(g27035), .A1(g23377), .A2(g26606) );
  AND2_X1 AND2_3052( .ZN(g27042), .A1(g21996), .A2(g26608) );
  AND2_X1 AND2_3053( .ZN(g27043), .A1(g23349), .A2(g26609) );
  AND2_X1 AND2_3054( .ZN(g27044), .A1(g22016), .A2(g26610) );
  AND2_X1 AND2_3055( .ZN(g27045), .A1(g23372), .A2(g26611) );
  AND2_X1 AND2_3056( .ZN(g27046), .A1(g22093), .A2(g26612) );
  AND2_X1 AND2_3057( .ZN(g27047), .A1(g23344), .A2(g26613) );
  AND2_X1 AND2_3058( .ZN(g27048), .A1(g22009), .A2(g26614) );
  AND2_X1 AND2_3059( .ZN(g27049), .A1(g23353), .A2(g26615) );
  AND2_X1 AND2_3060( .ZN(g27050), .A1(g23381), .A2(g26617) );
  AND2_X1 AND2_3061( .ZN(g27052), .A1(g4885), .A2(g26358) );
  AND2_X1 AND2_3062( .ZN(g27053), .A1(g23368), .A2(g26619) );
  AND2_X1 AND2_3063( .ZN(g27054), .A1(g22083), .A2(g26620) );
  AND2_X1 AND2_3064( .ZN(g27055), .A1(g22005), .A2(g26621) );
  AND2_X1 AND2_3065( .ZN(g27056), .A1(g22069), .A2(g26622) );
  AND2_X1 AND2_3066( .ZN(g27057), .A1(g23377), .A2(g26623) );
  AND2_X1 AND2_3067( .ZN(g27058), .A1(g22108), .A2(g26624) );
  AND2_X1 AND2_3068( .ZN(g27059), .A1(g23349), .A2(g26625) );
  AND2_X1 AND2_3069( .ZN(g27060), .A1(g22016), .A2(g26626) );
  AND2_X1 AND2_3070( .ZN(g27061), .A1(g23372), .A2(g26627) );
  AND2_X1 AND2_3071( .ZN(g27062), .A1(g22093), .A2(g26628) );
  AND2_X1 AND2_3072( .ZN(g27063), .A1(g23388), .A2(g26629) );
  AND2_X1 AND2_3073( .ZN(g27070), .A1(g22009), .A2(g26631) );
  AND2_X1 AND2_3074( .ZN(g27071), .A1(g23353), .A2(g26632) );
  AND2_X1 AND2_3075( .ZN(g27072), .A1(g22021), .A2(g26633) );
  AND2_X1 AND2_3076( .ZN(g27073), .A1(g23381), .A2(g26634) );
  AND2_X1 AND2_3077( .ZN(g27074), .A1(g22118), .A2(g26635) );
  AND2_X1 AND2_3078( .ZN(g27076), .A1(g5024), .A2(g26393) );
  AND2_X1 AND2_3079( .ZN(g27077), .A1(g22083), .A2(g26636) );
  AND2_X1 AND2_3080( .ZN(g27079), .A1(g5044), .A2(g26401) );
  AND2_X1 AND2_3081( .ZN(g27080), .A1(g23377), .A2(g26637) );
  AND2_X1 AND2_3082( .ZN(g27081), .A1(g22108), .A2(g26638) );
  AND2_X1 AND2_3083( .ZN(g27082), .A1(g22016), .A2(g26639) );
  AND2_X2 AND2_3084( .ZN(g27083), .A1(g22093), .A2(g26640) );
  AND2_X2 AND2_3085( .ZN(g27084), .A1(g23388), .A2(g26641) );
  AND2_X1 AND2_3086( .ZN(g27085), .A1(g22134), .A2(g26642) );
  AND2_X1 AND2_3087( .ZN(g27086), .A1(g23353), .A2(g26643) );
  AND2_X1 AND2_3088( .ZN(g27087), .A1(g22021), .A2(g26644) );
  AND2_X1 AND2_3089( .ZN(g27088), .A1(g23381), .A2(g26645) );
  AND2_X1 AND2_3090( .ZN(g27089), .A1(g22118), .A2(g26646) );
  AND2_X1 AND2_3091( .ZN(g27090), .A1(g23395), .A2(g26647) );
  AND2_X1 AND2_3092( .ZN(g27091), .A1(g5142), .A2(g26429) );
  AND2_X1 AND2_3093( .ZN(g27092), .A1(g5153), .A2(g26434) );
  AND2_X1 AND2_3094( .ZN(g27093), .A1(g22108), .A2(g26648) );
  AND2_X1 AND2_3095( .ZN(g27095), .A1(g5173), .A2(g26442) );
  AND2_X1 AND2_3096( .ZN(g27096), .A1(g23388), .A2(g26649) );
  AND2_X1 AND2_3097( .ZN(g27097), .A1(g22134), .A2(g26650) );
  AND2_X1 AND2_3098( .ZN(g27098), .A1(g22021), .A2(g26651) );
  AND2_X1 AND2_3099( .ZN(g27099), .A1(g22118), .A2(g26652) );
  AND2_X1 AND2_3100( .ZN(g27100), .A1(g23395), .A2(g26653) );
  AND2_X1 AND2_3101( .ZN(g27101), .A1(g22157), .A2(g26654) );
  AND2_X1 AND2_3102( .ZN(g27103), .A1(g5235), .A2(g26461) );
  AND2_X1 AND2_3103( .ZN(g27104), .A1(g5246), .A2(g26466) );
  AND2_X1 AND2_3104( .ZN(g27105), .A1(g22134), .A2(g26656) );
  AND2_X1 AND2_3105( .ZN(g27107), .A1(g5266), .A2(g26474) );
  AND2_X1 AND2_3106( .ZN(g27108), .A1(g23395), .A2(g26657) );
  AND2_X1 AND2_3107( .ZN(g27109), .A1(g22157), .A2(g26658) );
  AND2_X1 AND2_3108( .ZN(g27110), .A1(g5298), .A2(g26485) );
  AND2_X1 AND2_3109( .ZN(g27111), .A1(g5309), .A2(g26490) );
  AND2_X1 AND2_3110( .ZN(g27112), .A1(g22157), .A2(g26662) );
  AND2_X1 AND2_3111( .ZN(g27115), .A1(g5335), .A2(g26501) );
  AND2_X1 AND2_3112( .ZN(g27178), .A1(g26110), .A2(g22213) );
  AND3_X1 AND3_253( .ZN(g27181), .A1(g16570), .A2(g26508), .A3(g13614) );
  AND2_X1 AND2_3113( .ZN(g27182), .A1(g26151), .A2(g22217) );
  AND2_X1 AND2_3114( .ZN(g27185), .A1(g26126), .A2(g22230) );
  AND3_X1 AND3_254( .ZN(g27187), .A1(g16594), .A2(g26516), .A3(g13626) );
  AND2_X1 AND2_3115( .ZN(g27240), .A1(g26905), .A2(g22241) );
  AND2_X1 AND2_3116( .ZN(g27241), .A1(g10730), .A2(g26934) );
  AND2_X1 AND2_3117( .ZN(g27242), .A1(g26793), .A2(g8357) );
  AND2_X1 AND2_3118( .ZN(g27244), .A1(g26914), .A2(g22258) );
  AND2_X1 AND2_3119( .ZN(g27245), .A1(g26877), .A2(g22286) );
  AND2_X1 AND2_3120( .ZN(g27246), .A1(g26988), .A2(g16676) );
  AND2_X1 AND2_3121( .ZN(g27247), .A1(g27011), .A2(g16702) );
  AND2_X1 AND2_3122( .ZN(g27248), .A1(g27037), .A2(g16733) );
  AND2_X1 AND2_3123( .ZN(g27249), .A1(g27065), .A2(g16775) );
  AND2_X1 AND2_3124( .ZN(g27355), .A1(g61), .A2(g26837) );
  AND2_X1 AND2_3125( .ZN(g27356), .A1(g65), .A2(g26987) );
  AND2_X1 AND2_3126( .ZN(g27358), .A1(g749), .A2(g26846) );
  AND2_X1 AND2_3127( .ZN(g27359), .A1(g753), .A2(g27010) );
  AND2_X1 AND2_3128( .ZN(g27364), .A1(g1435), .A2(g26855) );
  AND2_X1 AND2_3129( .ZN(g27365), .A1(g1439), .A2(g27036) );
  AND2_X1 AND2_3130( .ZN(g27370), .A1(g27126), .A2(g8874) );
  AND2_X1 AND2_3131( .ZN(g27371), .A1(g2129), .A2(g26861) );
  AND2_X1 AND2_3132( .ZN(g27372), .A1(g2133), .A2(g27064) );
  AND2_X1 AND2_3133( .ZN(g27394), .A1(g17802), .A2(g27134) );
  AND2_X1 AND2_3134( .ZN(g27396), .A1(g692), .A2(g27135) );
  AND2_X1 AND2_3135( .ZN(g27407), .A1(g17914), .A2(g27136) );
  AND2_X1 AND2_3136( .ZN(g27409), .A1(g1378), .A2(g27137) );
  AND2_X1 AND2_3137( .ZN(g27425), .A1(g18025), .A2(g27138) );
  AND2_X1 AND2_3138( .ZN(g27427), .A1(g2072), .A2(g27139) );
  AND2_X1 AND2_3139( .ZN(g27446), .A1(g18142), .A2(g27141) );
  AND2_X1 AND2_3140( .ZN(g27448), .A1(g2766), .A2(g27142) );
  AND2_X1 AND2_3141( .ZN(g27495), .A1(g23945), .A2(g27146) );
  AND2_X1 AND2_3142( .ZN(g27509), .A1(g23945), .A2(g27148) );
  AND2_X2 AND2_3143( .ZN(g27516), .A1(g23974), .A2(g27151) );
  AND2_X2 AND2_3144( .ZN(g27530), .A1(g23945), .A2(g27153) );
  AND2_X1 AND2_3145( .ZN(g27534), .A1(g23974), .A2(g27155) );
  AND2_X1 AND2_3146( .ZN(g27541), .A1(g24004), .A2(g27159) );
  AND2_X1 AND2_3147( .ZN(g27552), .A1(g23974), .A2(g27162) );
  AND2_X1 AND2_3148( .ZN(g27554), .A1(g24004), .A2(g27164) );
  AND2_X1 AND2_3149( .ZN(g27561), .A1(g24038), .A2(g27167) );
  AND2_X1 AND2_3150( .ZN(g27568), .A1(g24004), .A2(g27172) );
  AND2_X1 AND2_3151( .ZN(g27570), .A1(g24038), .A2(g27173) );
  AND2_X1 AND2_3152( .ZN(g27578), .A1(g24038), .A2(g27177) );
  AND2_X1 AND2_3153( .ZN(g27656), .A1(g26796), .A2(g11004) );
  AND2_X1 AND2_3154( .ZN(g27657), .A1(g27114), .A2(g11051) );
  AND2_X1 AND2_3155( .ZN(g27659), .A1(g27132), .A2(g11114) );
  AND2_X1 AND2_3156( .ZN(g27660), .A1(g26835), .A2(g11117) );
  AND2_X1 AND2_3157( .ZN(g27661), .A1(g26841), .A2(g11173) );
  AND2_X1 AND2_3158( .ZN(g27666), .A1(g26849), .A2(g11243) );
  AND2_X1 AND2_3159( .ZN(g27671), .A1(g26885), .A2(g22212) );
  AND2_X1 AND2_3160( .ZN(g27673), .A1(g26854), .A2(g11312) );
  AND2_X1 AND2_3161( .ZN(g27679), .A1(g26782), .A2(g11386) );
  AND2_X1 AND2_3162( .ZN(g27680), .A1(g26983), .A2(g11392) );
  AND2_X1 AND2_3163( .ZN(g27681), .A1(g26788), .A2(g11456) );
  AND2_X1 AND2_3164( .ZN(g27719), .A1(g27496), .A2(g20649) );
  AND2_X1 AND2_3165( .ZN(g27720), .A1(g27481), .A2(g20652) );
  AND2_X1 AND2_3166( .ZN(g27721), .A1(g27579), .A2(g20655) );
  AND2_X1 AND2_3167( .ZN(g27723), .A1(g27464), .A2(g20679) );
  AND2_X1 AND2_3168( .ZN(g27725), .A1(g27532), .A2(g20704) );
  AND2_X1 AND2_3169( .ZN(g27726), .A1(g27531), .A2(g20732) );
  AND2_X1 AND2_3170( .ZN(g27727), .A1(g27414), .A2(g19301) );
  AND2_X1 AND2_3171( .ZN(g27728), .A1(g27564), .A2(g20766) );
  AND2_X1 AND2_3172( .ZN(g27729), .A1(g27435), .A2(g19322) );
  AND2_X1 AND2_3173( .ZN(g27730), .A1(g27454), .A2(g19349) );
  AND2_X1 AND2_3174( .ZN(g27731), .A1(g27470), .A2(g19383) );
  AND2_X1 AND2_3175( .ZN(g27732), .A1(g27492), .A2(g16758) );
  AND2_X1 AND2_3176( .ZN(g27733), .A1(g27513), .A2(g16785) );
  AND2_X1 AND2_3177( .ZN(g27734), .A1(g27538), .A2(g16814) );
  AND2_X1 AND2_3178( .ZN(g27737), .A1(g27558), .A2(g16832) );
  AND2_X1 AND2_3179( .ZN(g27770), .A1(g5642), .A2(g27449) );
  AND2_X1 AND2_3180( .ZN(g27772), .A1(g5680), .A2(g27465) );
  AND2_X1 AND2_3181( .ZN(g27773), .A1(g5732), .A2(g27484) );
  AND2_X1 AND2_3182( .ZN(g27774), .A1(g5702), .A2(g27361) );
  AND2_X1 AND2_3183( .ZN(g27775), .A1(g5790), .A2(g27506) );
  AND2_X1 AND2_3184( .ZN(g27779), .A1(g5760), .A2(g27367) );
  AND2_X1 AND2_3185( .ZN(g27783), .A1(g5819), .A2(g27373) );
  AND2_X1 AND2_3186( .ZN(g27790), .A1(g5875), .A2(g27376) );
  AND2_X1 AND2_3187( .ZN(g27904), .A1(g13873), .A2(g27387) );
  AND2_X1 AND2_3188( .ZN(g27908), .A1(g13886), .A2(g27391) );
  AND2_X1 AND2_3189( .ZN(g27909), .A1(g13895), .A2(g27397) );
  AND2_X1 AND2_3190( .ZN(g27913), .A1(g4017), .A2(g27401) );
  AND2_X1 AND2_3191( .ZN(g27914), .A1(g13927), .A2(g27404) );
  AND2_X1 AND2_3192( .ZN(g27915), .A1(g13936), .A2(g27410) );
  AND2_X1 AND2_3193( .ZN(g27922), .A1(g4112), .A2(g27416) );
  AND2_X1 AND2_3194( .ZN(g27923), .A1(g4144), .A2(g27419) );
  AND2_X1 AND2_3195( .ZN(g27924), .A1(g13983), .A2(g27422) );
  AND2_X2 AND2_3196( .ZN(g27926), .A1(g13992), .A2(g27428) );
  AND2_X2 AND2_3197( .ZN(g27931), .A1(g4221), .A2(g27432) );
  AND2_X2 AND2_3198( .ZN(g27935), .A1(g4251), .A2(g27437) );
  AND2_X1 AND2_3199( .ZN(g27936), .A1(g4283), .A2(g27440) );
  AND2_X1 AND2_3200( .ZN(g27938), .A1(g14053), .A2(g27443) );
  AND2_X1 AND2_3201( .ZN(g27945), .A1(g4376), .A2(g27451) );
  AND2_X1 AND2_3202( .ZN(g27949), .A1(g4406), .A2(g27456) );
  AND2_X1 AND2_3203( .ZN(g27951), .A1(g4438), .A2(g27459) );
  AND2_X1 AND2_3204( .ZN(g27963), .A1(g4545), .A2(g27467) );
  AND2_X1 AND2_3205( .ZN(g27968), .A1(g4575), .A2(g27472) );
  AND2_X1 AND2_3206( .ZN(g27970), .A1(g14238), .A2(g27475) );
  AND2_X1 AND2_3207( .ZN(g27984), .A1(g4721), .A2(g27486) );
  AND2_X1 AND2_3208( .ZN(g27985), .A1(g14342), .A2(g27489) );
  AND2_X1 AND2_3209( .ZN(g27991), .A1(g14360), .A2(g27498) );
  AND2_X1 AND2_3210( .ZN(g28008), .A1(g27590), .A2(g9770) );
  AND2_X1 AND2_3211( .ZN(g28009), .A1(g14454), .A2(g27510) );
  AND2_X1 AND2_3212( .ZN(g28015), .A1(g14472), .A2(g27518) );
  AND2_X1 AND2_3213( .ZN(g28027), .A1(g27590), .A2(g9895) );
  AND2_X1 AND2_3214( .ZN(g28028), .A1(g27595), .A2(g9898) );
  AND2_X1 AND2_3215( .ZN(g28035), .A1(g27599), .A2(g9916) );
  AND2_X1 AND2_3216( .ZN(g28036), .A1(g14541), .A2(g27535) );
  AND2_X1 AND2_3217( .ZN(g28042), .A1(g14559), .A2(g27543) );
  AND2_X1 AND2_3218( .ZN(g28050), .A1(g27590), .A2(g10018) );
  AND2_X1 AND2_3219( .ZN(g28051), .A1(g27595), .A2(g10021) );
  AND2_X1 AND2_3220( .ZN(g28057), .A1(g27599), .A2(g10049) );
  AND2_X1 AND2_3221( .ZN(g28058), .A1(g27604), .A2(g10052) );
  AND2_X1 AND2_3222( .ZN(g28065), .A1(g27608), .A2(g10070) );
  AND2_X1 AND2_3223( .ZN(g28066), .A1(g14596), .A2(g27555) );
  AND2_X1 AND2_3224( .ZN(g28073), .A1(g27595), .A2(g10109) );
  AND2_X1 AND2_3225( .ZN(g28079), .A1(g27599), .A2(g10127) );
  AND2_X1 AND2_3226( .ZN(g28080), .A1(g27604), .A2(g10130) );
  AND2_X1 AND2_3227( .ZN(g28086), .A1(g27608), .A2(g10158) );
  AND2_X1 AND2_3228( .ZN(g28087), .A1(g27613), .A2(g10161) );
  AND2_X1 AND2_3229( .ZN(g28094), .A1(g27617), .A2(g10179) );
  AND2_X1 AND2_3230( .ZN(g28098), .A1(g27604), .A2(g10214) );
  AND2_X1 AND2_3231( .ZN(g28104), .A1(g27608), .A2(g10232) );
  AND2_X1 AND2_3232( .ZN(g28105), .A1(g27613), .A2(g10235) );
  AND2_X1 AND2_3233( .ZN(g28111), .A1(g27617), .A2(g10263) );
  AND2_X1 AND2_3234( .ZN(g28112), .A1(g27622), .A2(g10266) );
  AND2_X1 AND2_3235( .ZN(g28116), .A1(g27613), .A2(g10316) );
  AND2_X1 AND2_3236( .ZN(g28122), .A1(g27617), .A2(g10334) );
  AND2_X1 AND2_3237( .ZN(g28123), .A1(g27622), .A2(g10337) );
  AND2_X1 AND2_3238( .ZN(g28127), .A1(g27622), .A2(g10409) );
  AND2_X1 AND2_3239( .ZN(g28171), .A1(g27349), .A2(g10898) );
  AND2_X1 AND2_3240( .ZN(g28176), .A1(g27349), .A2(g10940) );
  AND2_X1 AND2_3241( .ZN(g28188), .A1(g27349), .A2(g11008) );
  AND2_X1 AND2_3242( .ZN(g28193), .A1(g27573), .A2(g21914) );
  AND2_X1 AND2_3243( .ZN(g28319), .A1(g27855), .A2(g22246) );
  AND2_X1 AND2_3244( .ZN(g28320), .A1(g27854), .A2(g20637) );
  AND2_X1 AND2_3245( .ZN(g28322), .A1(g27937), .A2(g13868) );
  AND2_X1 AND2_3246( .ZN(g28323), .A1(g8580), .A2(g27838) );
  AND2_X1 AND2_3247( .ZN(g28324), .A1(g27810), .A2(g20659) );
  AND2_X1 AND2_3248( .ZN(g28326), .A1(g27865), .A2(g22274) );
  AND2_X1 AND2_3249( .ZN(g28327), .A1(g27900), .A2(g22275) );
  AND2_X1 AND2_3250( .ZN(g28329), .A1(g27823), .A2(g20708) );
  AND2_X1 AND2_3251( .ZN(g28330), .A1(g27864), .A2(g20711) );
  AND2_X1 AND2_3252( .ZN(g28331), .A1(g27802), .A2(g22307) );
  AND2_X1 AND2_3253( .ZN(g28332), .A1(g27883), .A2(g22331) );
  AND2_X1 AND2_3254( .ZN(g28333), .A1(g27882), .A2(g20772) );
  AND2_X1 AND2_3255( .ZN(g28334), .A1(g27842), .A2(g20793) );
  AND2_X2 AND2_3256( .ZN(g28335), .A1(g27814), .A2(g22343) );
  AND2_X2 AND2_3257( .ZN(g28336), .A1(g27896), .A2(g20810) );
  AND2_X1 AND2_3258( .ZN(g28337), .A1(g28002), .A2(g19448) );
  AND2_X1 AND2_3259( .ZN(g28338), .A1(g28029), .A2(g19475) );
  AND2_X1 AND2_3260( .ZN(g28339), .A1(g28059), .A2(g19498) );
  AND2_X1 AND2_3261( .ZN(g28340), .A1(g28088), .A2(g19519) );
  AND2_X1 AND2_3262( .ZN(g28373), .A1(g56), .A2(g27969) );
  AND2_X1 AND2_3263( .ZN(g28376), .A1(g744), .A2(g27990) );
  AND2_X1 AND2_3264( .ZN(g28378), .A1(g52), .A2(g27776) );
  AND3_X1 AND3_255( .ZN(g28379), .A1(g27868), .A2(g19390), .A3(g19369) );
  AND2_X1 AND2_3265( .ZN(g28380), .A1(g1430), .A2(g28014) );
  AND2_X1 AND2_3266( .ZN(g28381), .A1(g28157), .A2(g9815) );
  AND2_X1 AND2_3267( .ZN(g28383), .A1(g740), .A2(g27780) );
  AND2_X1 AND2_3268( .ZN(g28385), .A1(g2124), .A2(g28041) );
  AND2_X1 AND2_3269( .ZN(g28387), .A1(g1426), .A2(g27787) );
  AND2_X1 AND2_3270( .ZN(g28389), .A1(g2120), .A2(g27794) );
  AND2_X1 AND2_3271( .ZN(g28396), .A1(g7754), .A2(g27806) );
  AND2_X1 AND2_3272( .ZN(g28398), .A1(g7769), .A2(g27817) );
  AND2_X1 AND2_3273( .ZN(g28399), .A1(g7776), .A2(g27820) );
  AND2_X1 AND2_3274( .ZN(g28401), .A1(g7782), .A2(g27831) );
  AND2_X1 AND2_3275( .ZN(g28402), .A1(g7785), .A2(g27839) );
  AND2_X1 AND2_3276( .ZN(g28404), .A1(g7792), .A2(g27843) );
  AND2_X1 AND2_3277( .ZN(g28405), .A1(g7796), .A2(g27847) );
  AND2_X1 AND2_3278( .ZN(g28407), .A1(g7799), .A2(g27858) );
  AND2_X1 AND2_3279( .ZN(g28408), .A1(g7806), .A2(g27861) );
  AND2_X1 AND2_3280( .ZN(g28411), .A1(g7809), .A2(g27872) );
  AND2_X1 AND2_3281( .ZN(g28412), .A1(g7812), .A2(g27879) );
  AND2_X1 AND2_3282( .ZN(g28416), .A1(g7823), .A2(g27889) );
  AND2_X1 AND2_3283( .ZN(g28422), .A1(g17640), .A2(g28150) );
  AND2_X1 AND2_3284( .ZN(g28423), .A1(g17724), .A2(g28152) );
  AND2_X1 AND2_3285( .ZN(g28424), .A1(g17741), .A2(g28153) );
  AND2_X1 AND2_3286( .ZN(g28426), .A1(g28128), .A2(g9170) );
  AND2_X1 AND2_3287( .ZN(g28427), .A1(g26092), .A2(g28154) );
  AND2_X1 AND2_3288( .ZN(g28428), .A1(g17825), .A2(g28155) );
  AND2_X1 AND2_3289( .ZN(g28429), .A1(g17842), .A2(g28156) );
  AND2_X1 AND2_3290( .ZN(g28430), .A1(g28128), .A2(g9196) );
  AND2_X1 AND2_3291( .ZN(g28431), .A1(g26092), .A2(g28158) );
  AND2_X1 AND2_3292( .ZN(g28433), .A1(g28133), .A2(g9212) );
  AND2_X1 AND2_3293( .ZN(g28434), .A1(g26114), .A2(g28159) );
  AND2_X1 AND2_3294( .ZN(g28435), .A1(g17937), .A2(g28160) );
  AND2_X1 AND2_3295( .ZN(g28436), .A1(g17954), .A2(g28161) );
  AND2_X1 AND2_3296( .ZN(g28438), .A1(g17882), .A2(g27919) );
  AND2_X1 AND2_3297( .ZN(g28439), .A1(g28128), .A2(g9242) );
  AND2_X2 AND2_3298( .ZN(g28440), .A1(g26092), .A2(g28162) );
  AND2_X2 AND2_3299( .ZN(g28441), .A1(g28133), .A2(g9257) );
  AND2_X1 AND2_3300( .ZN(g28442), .A1(g26114), .A2(g28163) );
  AND2_X1 AND2_3301( .ZN(g28444), .A1(g28137), .A2(g9273) );
  AND2_X1 AND2_3302( .ZN(g28445), .A1(g26121), .A2(g28164) );
  AND2_X1 AND2_3303( .ZN(g28446), .A1(g18048), .A2(g28165) );
  AND2_X1 AND2_3304( .ZN(g28448), .A1(g17974), .A2(g27928) );
  AND2_X1 AND2_3305( .ZN(g28450), .A1(g17993), .A2(g27932) );
  AND2_X1 AND2_3306( .ZN(g28451), .A1(g28133), .A2(g9320) );
  AND2_X1 AND2_3307( .ZN(g28452), .A1(g26114), .A2(g28166) );
  AND2_X1 AND2_3308( .ZN(g28453), .A1(g28137), .A2(g9335) );
  AND2_X1 AND2_3309( .ZN(g28454), .A1(g26121), .A2(g28167) );
  AND2_X1 AND2_3310( .ZN(g28456), .A1(g28141), .A2(g9351) );
  AND2_X1 AND2_3311( .ZN(g28457), .A1(g26131), .A2(g28168) );
  AND2_X1 AND2_3312( .ZN(g28459), .A1(g18074), .A2(g27939) );
  AND2_X1 AND2_3313( .ZN(g28460), .A1(g18091), .A2(g27942) );
  AND2_X1 AND2_3314( .ZN(g28462), .A1(g18110), .A2(g27946) );
  AND2_X1 AND2_3315( .ZN(g28463), .A1(g28137), .A2(g9401) );
  AND2_X1 AND2_3316( .ZN(g28464), .A1(g26121), .A2(g28169) );
  AND2_X1 AND2_3317( .ZN(g28465), .A1(g28141), .A2(g9416) );
  AND2_X1 AND2_3318( .ZN(g28466), .A1(g26131), .A2(g28170) );
  AND2_X1 AND2_3319( .ZN(g28468), .A1(g18265), .A2(g28172) );
  AND2_X1 AND2_3320( .ZN(g28469), .A1(g18179), .A2(g27952) );
  AND2_X1 AND2_3321( .ZN(g28471), .A1(g18190), .A2(g27956) );
  AND2_X1 AND2_3322( .ZN(g28472), .A1(g18207), .A2(g27959) );
  AND2_X1 AND2_3323( .ZN(g28474), .A1(g18226), .A2(g27965) );
  AND2_X1 AND2_3324( .ZN(g28475), .A1(g28141), .A2(g9498) );
  AND2_X1 AND2_3325( .ZN(g28476), .A1(g26131), .A2(g28173) );
  AND2_X1 AND2_3326( .ZN(g28477), .A1(g18341), .A2(g28174) );
  AND2_X1 AND2_3327( .ZN(g28478), .A1(g18358), .A2(g28175) );
  AND2_X1 AND2_3328( .ZN(g28479), .A1(g18286), .A2(g27973) );
  AND2_X1 AND2_3329( .ZN(g28480), .A1(g18297), .A2(g27977) );
  AND2_X1 AND2_3330( .ZN(g28481), .A1(g18314), .A2(g27981) );
  AND2_X1 AND2_3331( .ZN(g28484), .A1(g18436), .A2(g28177) );
  AND2_X1 AND2_3332( .ZN(g28485), .A1(g18453), .A2(g28178) );
  AND2_X1 AND2_3333( .ZN(g28486), .A1(g18379), .A2(g27994) );
  AND2_X1 AND2_3334( .ZN(g28487), .A1(g18390), .A2(g27999) );
  AND2_X1 AND2_3335( .ZN(g28492), .A1(g18509), .A2(g28186) );
  AND2_X1 AND2_3336( .ZN(g28493), .A1(g18526), .A2(g28187) );
  AND2_X1 AND2_3337( .ZN(g28494), .A1(g18474), .A2(g28018) );
  AND2_X1 AND2_3338( .ZN(g28497), .A1(g18573), .A2(g28190) );
  AND2_X1 AND2_3339( .ZN(g28657), .A1(g27925), .A2(g13700) );
  AND2_X1 AND2_3340( .ZN(g28659), .A1(g27917), .A2(g13736) );
  AND2_X1 AND2_3341( .ZN(g28660), .A1(g27916), .A2(g11911) );
  AND2_X1 AND2_3342( .ZN(g28662), .A1(g27911), .A2(g11951) );
  AND2_X1 AND2_3343( .ZN(g28663), .A1(g27906), .A2(g11997) );
  AND2_X1 AND2_3344( .ZN(g28664), .A1(g27997), .A2(g12055) );
  AND2_X1 AND2_3345( .ZN(g28665), .A1(g27827), .A2(g22222) );
  AND2_X1 AND2_3346( .ZN(g28666), .A1(g27980), .A2(g12106) );
  AND2_X1 AND2_3347( .ZN(g28667), .A1(g27964), .A2(g13852) );
  AND2_X1 AND2_3348( .ZN(g28669), .A1(g27897), .A2(g22233) );
  AND2_X1 AND2_3349( .ZN(g28670), .A1(g27798), .A2(g21935) );
  AND2_X1 AND2_3350( .ZN(g28671), .A1(g27962), .A2(g12161) );
  AND2_X1 AND2_3351( .ZN(g28672), .A1(g27950), .A2(g13859) );
  AND2_X1 AND2_3352( .ZN(g28707), .A1(g12436), .A2(g28379) );
  AND2_X1 AND2_3353( .ZN(g28708), .A1(g28392), .A2(g22260) );
  AND2_X1 AND2_3354( .ZN(g28709), .A1(g28400), .A2(g22261) );
  AND2_X1 AND2_3355( .ZN(g28710), .A1(g28403), .A2(g22262) );
  AND2_X1 AND2_3356( .ZN(g28711), .A1(g10749), .A2(g28415) );
  AND2_X1 AND2_3357( .ZN(g28712), .A1(g28406), .A2(g22276) );
  AND2_X1 AND2_3358( .ZN(g28713), .A1(g28410), .A2(g22290) );
  AND2_X1 AND2_3359( .ZN(g28714), .A1(g28394), .A2(g22306) );
  AND2_X1 AND2_3360( .ZN(g28715), .A1(g28414), .A2(g22332) );
  AND2_X1 AND2_3361( .ZN(g28716), .A1(g28449), .A2(g19319) );
  AND2_X1 AND2_3362( .ZN(g28717), .A1(g28461), .A2(g19346) );
  AND2_X1 AND2_3363( .ZN(g28718), .A1(g28473), .A2(g19380) );
  AND2_X1 AND2_3364( .ZN(g28719), .A1(g28482), .A2(g19412) );
  AND2_X2 AND2_3365( .ZN(g28722), .A1(g28523), .A2(g16694) );
  AND2_X1 AND2_3366( .ZN(g28724), .A1(g28551), .A2(g16725) );
  AND2_X1 AND2_3367( .ZN(g28726), .A1(g28578), .A2(g16767) );
  AND2_X1 AND2_3368( .ZN(g28729), .A1(g28606), .A2(g16794) );
  AND2_X1 AND2_3369( .ZN(g28834), .A1(g5751), .A2(g28483) );
  AND2_X1 AND2_3370( .ZN(g28836), .A1(g5810), .A2(g28491) );
  AND2_X1 AND2_3371( .ZN(g28838), .A1(g5866), .A2(g28496) );
  AND2_X1 AND2_3372( .ZN(g28840), .A1(g5913), .A2(g28500) );
  AND2_X1 AND2_3373( .ZN(g28841), .A1(g27834), .A2(g28554) );
  AND2_X1 AND2_3374( .ZN(g28843), .A1(g27834), .A2(g28581) );
  AND2_X1 AND2_3375( .ZN(g28844), .A1(g27850), .A2(g28582) );
  AND2_X1 AND2_3376( .ZN(g28846), .A1(g27834), .A2(g28608) );
  AND2_X1 AND2_3377( .ZN(g28847), .A1(g27850), .A2(g28609) );
  AND2_X1 AND2_3378( .ZN(g28848), .A1(g27875), .A2(g28610) );
  AND2_X2 AND2_3379( .ZN(g28849), .A1(g27850), .A2(g28616) );
  AND2_X1 AND2_3380( .ZN(g28850), .A1(g27875), .A2(g28617) );
  AND2_X1 AND2_3381( .ZN(g28851), .A1(g27892), .A2(g28618) );
  AND2_X1 AND2_3382( .ZN(g28852), .A1(g27875), .A2(g28623) );
  AND2_X1 AND2_3383( .ZN(g28853), .A1(g27892), .A2(g28624) );
  AND2_X1 AND2_3384( .ZN(g28854), .A1(g27892), .A2(g28629) );
  AND2_X1 AND2_3385( .ZN(g28880), .A1(g13946), .A2(g28639) );
  AND2_X1 AND2_3386( .ZN(g28881), .A1(g28612), .A2(g9199) );
  AND2_X1 AND2_3387( .ZN(g28892), .A1(g14001), .A2(g28640) );
  AND2_X1 AND2_3388( .ZN(g28893), .A1(g28612), .A2(g9245) );
  AND2_X1 AND2_3389( .ZN(g28897), .A1(g14016), .A2(g28641) );
  AND2_X1 AND2_3390( .ZN(g28898), .A1(g28619), .A2(g9260) );
  AND2_X1 AND2_3391( .ZN(g28909), .A1(g14062), .A2(g28642) );
  AND2_X1 AND2_3392( .ZN(g28910), .A1(g28612), .A2(g9303) );
  AND2_X1 AND2_3393( .ZN(g28914), .A1(g14092), .A2(g28643) );
  AND2_X1 AND2_3394( .ZN(g28915), .A1(g28619), .A2(g9323) );
  AND2_X1 AND2_3395( .ZN(g28919), .A1(g14107), .A2(g28644) );
  AND2_X1 AND2_3396( .ZN(g28923), .A1(g28625), .A2(g9338) );
  AND2_X1 AND2_3397( .ZN(g28931), .A1(g14153), .A2(g28645) );
  AND2_X1 AND2_3398( .ZN(g28935), .A1(g14177), .A2(g28646) );
  AND2_X1 AND2_3399( .ZN(g28936), .A1(g28619), .A2(g9384) );
  AND2_X1 AND2_3400( .ZN(g28940), .A1(g14207), .A2(g28647) );
  AND2_X1 AND2_3401( .ZN(g28944), .A1(g28625), .A2(g9404) );
  AND2_X1 AND2_3402( .ZN(g28948), .A1(g14222), .A2(g28648) );
  AND2_X1 AND2_3403( .ZN(g28949), .A1(g28630), .A2(g9419) );
  AND2_X1 AND2_3404( .ZN(g28958), .A1(g14268), .A2(g28649) );
  AND2_X1 AND2_3405( .ZN(g28962), .A1(g14292), .A2(g28650) );
  AND2_X1 AND2_3406( .ZN(g28966), .A1(g28625), .A2(g9481) );
  AND2_X1 AND2_3407( .ZN(g28970), .A1(g14322), .A2(g28651) );
  AND2_X1 AND2_3408( .ZN(g28971), .A1(g28630), .A2(g9501) );
  AND2_X1 AND2_3409( .ZN(g28986), .A1(g14390), .A2(g28652) );
  AND2_X2 AND2_3410( .ZN(g28996), .A1(g14414), .A2(g28653) );
  AND2_X2 AND2_3411( .ZN(g28997), .A1(g28630), .A2(g9623) );
  AND2_X2 AND2_3412( .ZN(g29022), .A1(g14502), .A2(g28655) );
  AND2_X2 AND2_3413( .ZN(g29130), .A1(g28397), .A2(g22221) );
  AND2_X2 AND2_3414( .ZN(g29174), .A1(g29031), .A2(g20684) );
  AND2_X2 AND2_3415( .ZN(g29175), .A1(g29009), .A2(g20687) );
  AND2_X2 AND2_3416( .ZN(g29176), .A1(g29097), .A2(g20690) );
  AND2_X2 AND2_3417( .ZN(g29180), .A1(g28982), .A2(g20714) );
  AND2_X2 AND2_3418( .ZN(g29183), .A1(g29064), .A2(g20739) );
  AND2_X1 AND2_3419( .ZN(g29186), .A1(g29063), .A2(g20769) );
  AND2_X1 AND2_3420( .ZN(g29188), .A1(g29083), .A2(g20796) );
  AND2_X1 AND2_3421( .ZN(g29196), .A1(g15022), .A2(g28741) );
  AND2_X1 AND2_3422( .ZN(g29200), .A1(g15096), .A2(g28751) );
  AND2_X1 AND2_3423( .ZN(g29203), .A1(g15118), .A2(g28755) );
  AND2_X1 AND2_3424( .ZN(g29208), .A1(g15188), .A2(g28764) );
  AND2_X1 AND2_3425( .ZN(g29211), .A1(g15210), .A2(g28768) );
  AND2_X1 AND2_3426( .ZN(g29217), .A1(g15274), .A2(g28775) );
  AND2_X1 AND2_3427( .ZN(g29220), .A1(g15296), .A2(g28779) );
  AND2_X1 AND2_3428( .ZN(g29225), .A1(g15366), .A2(g28785) );
  AND2_X1 AND2_3429( .ZN(g29229), .A1(g9293), .A2(g28791) );
  AND2_X1 AND2_3430( .ZN(g29232), .A1(g9356), .A2(g28796) );
  AND2_X1 AND2_3431( .ZN(g29233), .A1(g9374), .A2(g28799) );
  AND2_X1 AND2_3432( .ZN(g29234), .A1(g9427), .A2(g28804) );
  AND2_X1 AND2_3433( .ZN(g29235), .A1(g9453), .A2(g28807) );
  AND2_X1 AND2_3434( .ZN(g29236), .A1(g9471), .A2(g28810) );
  AND2_X1 AND2_3435( .ZN(g29238), .A1(g9569), .A2(g28814) );
  AND2_X1 AND2_3436( .ZN(g29239), .A1(g9595), .A2(g28817) );
  AND2_X1 AND2_3437( .ZN(g29240), .A1(g9613), .A2(g28820) );
  AND2_X1 AND2_3438( .ZN(g29241), .A1(g9711), .A2(g28823) );
  AND2_X1 AND2_3439( .ZN(g29242), .A1(g9737), .A2(g28826) );
  AND2_X1 AND2_3440( .ZN(g29243), .A1(g9857), .A2(g28829) );
  AND2_X1 AND2_3441( .ZN(g29248), .A1(g28855), .A2(g8836) );
  AND2_X1 AND2_3442( .ZN(g29251), .A1(g28855), .A2(g8856) );
  AND2_X1 AND2_3443( .ZN(g29252), .A1(g28859), .A2(g8863) );
  AND2_X1 AND2_3444( .ZN(g29255), .A1(g28855), .A2(g8885) );
  AND2_X1 AND2_3445( .ZN(g29256), .A1(g28859), .A2(g8894) );
  AND2_X1 AND2_3446( .ZN(g29257), .A1(g28863), .A2(g8901) );
  AND2_X1 AND2_3447( .ZN(g29259), .A1(g28859), .A2(g8925) );
  AND2_X1 AND2_3448( .ZN(g29260), .A1(g28863), .A2(g8934) );
  AND2_X1 AND2_3449( .ZN(g29261), .A1(g28867), .A2(g8941) );
  AND2_X1 AND2_3450( .ZN(g29262), .A1(g28863), .A2(g8965) );
  AND2_X1 AND2_3451( .ZN(g29263), .A1(g28867), .A2(g8974) );
  AND2_X1 AND2_3452( .ZN(g29264), .A1(g28867), .A2(g8997) );
  AND2_X1 AND2_3453( .ZN(g29284), .A1(g29001), .A2(g28871) );
  AND2_X1 AND2_3454( .ZN(g29289), .A1(g29030), .A2(g28883) );
  AND2_X1 AND2_3455( .ZN(g29294), .A1(g29053), .A2(g28900) );
  AND2_X1 AND2_3456( .ZN(g29300), .A1(g29072), .A2(g28925) );
  AND2_X1 AND2_3457( .ZN(g29302), .A1(g29026), .A2(g28928) );
  AND2_X1 AND2_3458( .ZN(g29310), .A1(g28978), .A2(g28951) );
  AND2_X1 AND2_3459( .ZN(g29312), .A1(g29049), .A2(g28955) );
  AND2_X1 AND2_3460( .ZN(g29320), .A1(g29088), .A2(g28972) );
  AND2_X1 AND2_3461( .ZN(g29321), .A1(g29008), .A2(g28979) );
  AND2_X1 AND2_3462( .ZN(g29323), .A1(g29068), .A2(g28983) );
  AND2_X1 AND2_3463( .ZN(g29329), .A1(g29096), .A2(g29002) );
  AND2_X1 AND2_3464( .ZN(g29330), .A1(g29038), .A2(g29010) );
  AND2_X1 AND2_3465( .ZN(g29332), .A1(g29080), .A2(g29019) );
  AND2_X1 AND2_3466( .ZN(g29336), .A1(g29045), .A2(g29023) );
  AND2_X1 AND2_3467( .ZN(g29337), .A1(g29103), .A2(g29032) );
  AND2_X1 AND2_3468( .ZN(g29338), .A1(g29060), .A2(g29042) );
  AND2_X1 AND2_3469( .ZN(g29341), .A1(g29062), .A2(g29046) );
  AND2_X1 AND2_3470( .ZN(g29342), .A1(g29107), .A2(g29054) );
  AND2_X1 AND2_3471( .ZN(g29344), .A1(g29076), .A2(g29065) );
  AND2_X1 AND2_3472( .ZN(g29346), .A1(g29087), .A2(g29077) );
  AND2_X1 AND2_3473( .ZN(g29411), .A1(g29090), .A2(g21932) );
  AND2_X1 AND2_3474( .ZN(g29464), .A1(g29190), .A2(g8375) );
  AND2_X1 AND2_3475( .ZN(g29465), .A1(g29191), .A2(g8424) );
  AND2_X1 AND2_3476( .ZN(g29466), .A1(g8587), .A2(g29265) );
  AND2_X1 AND2_3477( .ZN(g29467), .A1(g29340), .A2(g19467) );
  AND2_X1 AND2_3478( .ZN(g29468), .A1(g29343), .A2(g19490) );
  AND2_X1 AND2_3479( .ZN(g29469), .A1(g29345), .A2(g19511) );
  AND2_X1 AND2_3480( .ZN(g29470), .A1(g29347), .A2(g19530) );
  AND2_X1 AND2_3481( .ZN(g29471), .A1(g21461), .A2(g29266) );
  AND2_X1 AND2_3482( .ZN(g29472), .A1(g21461), .A2(g29268) );
  AND2_X1 AND2_3483( .ZN(g29473), .A1(g21508), .A2(g29269) );
  AND2_X1 AND2_3484( .ZN(g29474), .A1(g21508), .A2(g29271) );
  AND2_X1 AND2_3485( .ZN(g29475), .A1(g21544), .A2(g29272) );
  AND2_X1 AND2_3486( .ZN(g29476), .A1(g21544), .A2(g29274) );
  AND2_X1 AND2_3487( .ZN(g29477), .A1(g21580), .A2(g29275) );
  AND2_X1 AND2_3488( .ZN(g29478), .A1(g21580), .A2(g29277) );
  AND2_X1 AND2_3489( .ZN(g29479), .A1(g21461), .A2(g29280) );
  AND2_X1 AND2_3490( .ZN(g29480), .A1(g21461), .A2(g29282) );
  AND2_X1 AND2_3491( .ZN(g29481), .A1(g21508), .A2(g29283) );
  AND2_X1 AND2_3492( .ZN(g29482), .A1(g21461), .A2(g29285) );
  AND2_X1 AND2_3493( .ZN(g29483), .A1(g21508), .A2(g29286) );
  AND2_X1 AND2_3494( .ZN(g29484), .A1(g21544), .A2(g29287) );
  AND2_X1 AND2_3495( .ZN(g29485), .A1(g21508), .A2(g29290) );
  AND2_X1 AND2_3496( .ZN(g29486), .A1(g21544), .A2(g29291) );
  AND2_X1 AND2_3497( .ZN(g29487), .A1(g21580), .A2(g29292) );
  AND2_X1 AND2_3498( .ZN(g29488), .A1(g21544), .A2(g29295) );
  AND2_X1 AND2_3499( .ZN(g29489), .A1(g21580), .A2(g29296) );
  AND2_X1 AND2_3500( .ZN(g29490), .A1(g21580), .A2(g29301) );
  AND2_X1 AND2_3501( .ZN(g29502), .A1(g29350), .A2(g8912) );
  AND2_X1 AND2_3502( .ZN(g29518), .A1(g28728), .A2(g29360) );
  AND2_X1 AND2_3503( .ZN(g29520), .A1(g28731), .A2(g29361) );
  AND2_X1 AND2_3504( .ZN(g29521), .A1(g28733), .A2(g29362) );
  AND2_X1 AND2_3505( .ZN(g29522), .A1(g27735), .A2(g29363) );
  AND2_X1 AND2_3506( .ZN(g29523), .A1(g28737), .A2(g29364) );
  AND2_X1 AND2_3507( .ZN(g29524), .A1(g28739), .A2(g29365) );
  AND2_X1 AND2_3508( .ZN(g29525), .A1(g29195), .A2(g29366) );
  AND2_X1 AND2_3509( .ZN(g29526), .A1(g27741), .A2(g29367) );
  AND2_X1 AND2_3510( .ZN(g29527), .A1(g28748), .A2(g29368) );
  AND2_X1 AND2_3511( .ZN(g29528), .A1(g28750), .A2(g29369) );
  AND2_X1 AND2_3512( .ZN(g29529), .A1(g29199), .A2(g29370) );
  AND2_X1 AND2_3513( .ZN(g29531), .A1(g29202), .A2(g29371) );
  AND2_X1 AND2_3514( .ZN(g29532), .A1(g27746), .A2(g29372) );
  AND2_X1 AND2_3515( .ZN(g29533), .A1(g28762), .A2(g29373) );
  AND2_X1 AND2_3516( .ZN(g29534), .A1(g29206), .A2(g29374) );
  AND2_X1 AND2_3517( .ZN(g29536), .A1(g29207), .A2(g29375) );
  AND2_X1 AND2_3518( .ZN(g29538), .A1(g29210), .A2(g29376) );
  AND2_X1 AND2_3519( .ZN(g29539), .A1(g27754), .A2(g29377) );
  AND2_X1 AND2_3520( .ZN(g29540), .A1(g26041), .A2(g29378) );
  AND2_X1 AND2_3521( .ZN(g29541), .A1(g29214), .A2(g29379) );
  AND2_X1 AND2_3522( .ZN(g29543), .A1(g29215), .A2(g29380) );
  AND2_X1 AND2_3523( .ZN(g29545), .A1(g29216), .A2(g29381) );
  AND2_X1 AND2_3524( .ZN(g29547), .A1(g29219), .A2(g29382) );
  AND2_X1 AND2_3525( .ZN(g29548), .A1(g28784), .A2(g29383) );
  AND2_X1 AND2_3526( .ZN(g29549), .A1(g26043), .A2(g29384) );
  AND2_X1 AND2_3527( .ZN(g29550), .A1(g29222), .A2(g29385) );
  AND2_X1 AND2_3528( .ZN(g29553), .A1(g29223), .A2(g29386) );
  AND2_X1 AND2_3529( .ZN(g29555), .A1(g29224), .A2(g29387) );
  AND2_X1 AND2_3530( .ZN(g29557), .A1(g28789), .A2(g29388) );
  AND2_X1 AND2_3531( .ZN(g29558), .A1(g28790), .A2(g29389) );
  AND2_X1 AND2_3532( .ZN(g29559), .A1(g26045), .A2(g29390) );
  AND2_X1 AND2_3533( .ZN(g29560), .A1(g29227), .A2(g29391) );
  AND2_X1 AND2_3534( .ZN(g29562), .A1(g29228), .A2(g29392) );
  AND2_X1 AND2_3535( .ZN(g29564), .A1(g28794), .A2(g29393) );
  AND2_X1 AND2_3536( .ZN(g29565), .A1(g28795), .A2(g29394) );
  AND2_X1 AND2_3537( .ZN(g29566), .A1(g26047), .A2(g29395) );
  AND2_X1 AND2_3538( .ZN(g29567), .A1(g29231), .A2(g29396) );
  AND2_X1 AND2_3539( .ZN(g29572), .A1(g28802), .A2(g29397) );
  AND2_X1 AND2_3540( .ZN(g29573), .A1(g28803), .A2(g29398) );
  AND2_X1 AND2_3541( .ZN(g29575), .A1(g28813), .A2(g29402) );
  AND2_X1 AND2_3542( .ZN(g29607), .A1(g29193), .A2(g11056) );
  AND2_X1 AND2_3543( .ZN(g29610), .A1(g29349), .A2(g11123) );
  AND2_X2 AND2_3544( .ZN(g29614), .A1(g29359), .A2(g11182) );
  AND2_X2 AND2_3545( .ZN(g29615), .A1(g29245), .A2(g11185) );
  AND2_X2 AND2_3546( .ZN(g29619), .A1(g29247), .A2(g11259) );
  AND2_X2 AND2_3547( .ZN(g29622), .A1(g29250), .A2(g11327) );
  AND2_X2 AND2_3548( .ZN(g29624), .A1(g29254), .A2(g11407) );
  AND2_X1 AND2_3549( .ZN(g29625), .A1(g29189), .A2(g11472) );
  AND2_X1 AND2_3550( .ZN(g29626), .A1(g29318), .A2(g11478) );
  AND2_X1 AND2_3551( .ZN(g29790), .A1(g29491), .A2(g10918) );
  AND2_X1 AND2_3552( .ZN(g29792), .A1(g29491), .A2(g10977) );
  AND2_X1 AND2_3553( .ZN(g29793), .A1(g29491), .A2(g11063) );
  AND2_X1 AND2_3554( .ZN(g29810), .A1(g29748), .A2(g22248) );
  AND2_X1 AND2_3555( .ZN(g29811), .A1(g29703), .A2(g20644) );
  AND2_X1 AND2_3556( .ZN(g29812), .A1(g29762), .A2(g12223) );
  AND2_X1 AND2_3557( .ZN(g29813), .A1(g29760), .A2(g13869) );
  AND2_X1 AND2_3558( .ZN(g29814), .A1(g29728), .A2(g22266) );
  AND2_X1 AND2_3559( .ZN(g29815), .A1(g29727), .A2(g20662) );
  AND2_X1 AND2_3560( .ZN(g29816), .A1(g29759), .A2(g13883) );
  AND2_X1 AND2_3561( .ZN(g29817), .A1(g29709), .A2(g20694) );
  AND2_X1 AND2_3562( .ZN(g29818), .A1(g29732), .A2(g22293) );
  AND2_X1 AND2_3563( .ZN(g29819), .A1(g29751), .A2(g22294) );
  AND2_X1 AND2_3564( .ZN(g29820), .A1(g29717), .A2(g20743) );
  AND2_X1 AND2_3565( .ZN(g29821), .A1(g29731), .A2(g20746) );
  AND2_X1 AND2_3566( .ZN(g29822), .A1(g29705), .A2(g22335) );
  AND2_X1 AND2_3567( .ZN(g29827), .A1(g29741), .A2(g22356) );
  AND2_X1 AND2_3568( .ZN(g29828), .A1(g29740), .A2(g20802) );
  AND2_X1 AND2_3569( .ZN(g29833), .A1(g29725), .A2(g20813) );
  AND2_X1 AND2_3570( .ZN(g29834), .A1(g29713), .A2(g22366) );
  AND2_X1 AND2_3571( .ZN(g29839), .A1(g29747), .A2(g20827) );
  AND3_X1 AND3_256( .ZN(g29909), .A1(g29735), .A2(g19420), .A3(g19401) );
  AND2_X1 AND2_3572( .ZN(g29910), .A1(g29779), .A2(g9961) );
  AND2_X1 AND2_3573( .ZN(g29942), .A1(g29771), .A2(g28877) );
  AND2_X1 AND2_3574( .ZN(g29944), .A1(g29782), .A2(g28889) );
  AND2_X1 AND2_3575( .ZN(g29945), .A1(g29773), .A2(g28894) );
  AND2_X1 AND2_3576( .ZN(g29946), .A1(g29778), .A2(g28906) );
  AND2_X1 AND2_3577( .ZN(g29947), .A1(g29785), .A2(g28911) );
  AND2_X1 AND2_3578( .ZN(g29948), .A1(g29775), .A2(g28916) );
  AND2_X1 AND2_3579( .ZN(g29949), .A1(g29781), .A2(g28932) );
  AND2_X1 AND2_3580( .ZN(g29950), .A1(g29788), .A2(g28937) );
  AND2_X1 AND2_3581( .ZN(g29951), .A1(g29777), .A2(g28945) );
  AND2_X1 AND2_3582( .ZN(g29952), .A1(g29784), .A2(g28959) );
  AND2_X1 AND2_3583( .ZN(g29953), .A1(g29791), .A2(g28967) );
  AND2_X1 AND2_3584( .ZN(g29954), .A1(g29770), .A2(g28975) );
  AND2_X1 AND2_3585( .ZN(g29955), .A1(g29787), .A2(g28993) );
  AND2_X1 AND2_3586( .ZN(g29956), .A1(g29780), .A2(g28998) );
  AND2_X1 AND2_3587( .ZN(g29957), .A1(g29772), .A2(g29005) );
  AND2_X1 AND2_3588( .ZN(g29958), .A1(g29783), .A2(g29027) );
  AND2_X1 AND2_3589( .ZN(g29959), .A1(g29774), .A2(g29035) );
  AND2_X1 AND2_3590( .ZN(g29960), .A1(g29786), .A2(g29050) );
  AND2_X1 AND2_3591( .ZN(g29961), .A1(g29776), .A2(g29057) );
  AND2_X1 AND2_3592( .ZN(g29962), .A1(g29789), .A2(g29069) );
  AND2_X1 AND2_3593( .ZN(g29963), .A1(g29758), .A2(g13737) );
  AND2_X1 AND2_3594( .ZN(g29964), .A1(g29757), .A2(g13786) );
  AND2_X1 AND2_3595( .ZN(g29965), .A1(g29756), .A2(g11961) );
  AND2_X1 AND2_3596( .ZN(g29966), .A1(g29755), .A2(g12004) );
  AND2_X1 AND2_3597( .ZN(g29967), .A1(g29754), .A2(g12066) );
  AND2_X1 AND2_3598( .ZN(g29968), .A1(g29765), .A2(g12119) );
  AND2_X1 AND2_3599( .ZN(g29969), .A1(g29721), .A2(g22237) );
  AND2_X1 AND2_3600( .ZN(g29970), .A1(g29764), .A2(g12178) );
  AND2_X1 AND2_3601( .ZN(g29971), .A1(g29763), .A2(g13861) );
  AND2_X1 AND2_3602( .ZN(g29980), .A1(g29881), .A2(g8324) );
  AND2_X1 AND2_3603( .ZN(g29981), .A1(g29869), .A2(g8330) );
  AND2_X1 AND2_3604( .ZN(g29982), .A1(g29893), .A2(g8336) );
  AND2_X1 AND2_3605( .ZN(g29983), .A1(g29885), .A2(g8344) );
  AND2_X1 AND2_3606( .ZN(g29984), .A1(g29873), .A2(g8351) );
  AND2_X1 AND2_3607( .ZN(g29985), .A1(g29897), .A2(g8363) );
  AND2_X1 AND2_3608( .ZN(g29986), .A1(g29877), .A2(g8366) );
  AND2_X1 AND2_3609( .ZN(g29987), .A1(g29889), .A2(g8369) );
  AND2_X1 AND2_3610( .ZN(g29988), .A1(g29881), .A2(g8382) );
  AND2_X1 AND2_3611( .ZN(g29989), .A1(g29893), .A2(g8391) );
  AND2_X1 AND2_3612( .ZN(g29990), .A1(g29885), .A2(g8397) );
  AND2_X1 AND2_3613( .ZN(g29991), .A1(g29901), .A2(g8403) );
  AND2_X1 AND2_3614( .ZN(g29992), .A1(g12441), .A2(g29909) );
  AND2_X1 AND2_3615( .ZN(g29993), .A1(g29897), .A2(g8411) );
  AND2_X1 AND2_3616( .ZN(g29994), .A1(g29889), .A2(g8418) );
  AND2_X1 AND2_3617( .ZN(g29995), .A1(g29893), .A2(g8434) );
  AND2_X1 AND2_3618( .ZN(g29996), .A1(g29901), .A2(g8443) );
  AND2_X1 AND2_3619( .ZN(g29997), .A1(g29918), .A2(g22277) );
  AND2_X1 AND2_3620( .ZN(g29998), .A1(g29922), .A2(g22278) );
  AND2_X1 AND2_3621( .ZN(g29999), .A1(g29924), .A2(g22279) );
  AND2_X1 AND2_3622( .ZN(g30000), .A1(g10767), .A2(g29930) );
  AND2_X1 AND2_3623( .ZN(g30001), .A1(g29897), .A2(g8449) );
  AND2_X1 AND2_3624( .ZN(g30002), .A1(g29905), .A2(g8455) );
  AND2_X1 AND2_3625( .ZN(g30003), .A1(g29901), .A2(g8469) );
  AND2_X1 AND2_3626( .ZN(g30004), .A1(g29926), .A2(g22295) );
  AND2_X1 AND2_3627( .ZN(g30005), .A1(g29905), .A2(g8478) );
  AND2_X1 AND2_3628( .ZN(g30006), .A1(g29928), .A2(g22310) );
  AND2_X1 AND2_3629( .ZN(g30007), .A1(g29905), .A2(g8494) );
  AND2_X1 AND2_3630( .ZN(g30008), .A1(g29919), .A2(g22334) );
  AND2_X1 AND2_3631( .ZN(g30009), .A1(g29929), .A2(g22357) );
  AND2_X1 AND2_3632( .ZN(g30077), .A1(g29823), .A2(g10963) );
  AND2_X1 AND2_3633( .ZN(g30079), .A1(g29823), .A2(g10988) );
  AND2_X1 AND2_3634( .ZN(g30080), .A1(g29829), .A2(g10996) );
  AND2_X1 AND2_3635( .ZN(g30081), .A1(g29823), .A2(g11022) );
  AND2_X1 AND2_3636( .ZN(g30082), .A1(g29829), .A2(g11036) );
  AND2_X1 AND2_3637( .ZN(g30083), .A1(g29835), .A2(g11048) );
  AND2_X1 AND2_3638( .ZN(g30085), .A1(g29829), .A2(g11092) );
  AND2_X1 AND2_3639( .ZN(g30086), .A1(g29835), .A2(g11108) );
  AND2_X1 AND2_3640( .ZN(g30087), .A1(g29840), .A2(g11120) );
  AND2_X1 AND2_3641( .ZN(g30088), .A1(g29844), .A2(g11138) );
  AND2_X1 AND2_3642( .ZN(g30089), .A1(g29835), .A2(g11160) );
  AND2_X1 AND2_3643( .ZN(g30090), .A1(g29840), .A2(g11176) );
  AND2_X1 AND2_3644( .ZN(g30091), .A1(g29844), .A2(g11202) );
  AND2_X1 AND2_3645( .ZN(g30092), .A1(g29849), .A2(g11205) );
  AND2_X1 AND2_3646( .ZN(g30093), .A1(g29853), .A2(g11222) );
  AND2_X1 AND2_3647( .ZN(g30094), .A1(g29840), .A2(g11246) );
  AND2_X1 AND2_3648( .ZN(g30095), .A1(g29857), .A2(g11265) );
  AND2_X1 AND2_3649( .ZN(g30096), .A1(g29844), .A2(g11268) );
  AND2_X1 AND2_3650( .ZN(g30097), .A1(g29849), .A2(g11271) );
  AND2_X1 AND2_3651( .ZN(g30098), .A1(g29853), .A2(g11284) );
  AND2_X1 AND2_3652( .ZN(g30099), .A1(g29861), .A2(g11287) );
  AND2_X1 AND2_3653( .ZN(g30100), .A1(g29865), .A2(g11306) );
  AND2_X1 AND2_3654( .ZN(g30101), .A1(g29857), .A2(g11341) );
  AND2_X1 AND2_3655( .ZN(g30102), .A1(g29849), .A2(g11348) );
  AND2_X1 AND2_3656( .ZN(g30103), .A1(g29869), .A2(g11358) );
  AND2_X1 AND2_3657( .ZN(g30104), .A1(g29853), .A2(g11361) );
  AND2_X1 AND2_3658( .ZN(g30105), .A1(g29861), .A2(g11364) );
  AND2_X1 AND2_3659( .ZN(g30106), .A1(g29865), .A2(g11379) );
  AND2_X1 AND2_3660( .ZN(g30107), .A1(g29873), .A2(g11382) );
  AND2_X1 AND2_3661( .ZN(g30108), .A1(g29877), .A2(g11401) );
  AND2_X1 AND2_3662( .ZN(g30109), .A1(g29857), .A2(g11411) );
  AND2_X1 AND2_3663( .ZN(g30110), .A1(g29881), .A2(g11417) );
  AND2_X1 AND2_3664( .ZN(g30111), .A1(g29869), .A2(g11425) );
  AND2_X1 AND2_3665( .ZN(g30112), .A1(g29861), .A2(g11432) );
  AND2_X1 AND2_3666( .ZN(g30113), .A1(g29885), .A2(g11444) );
  AND2_X1 AND2_3667( .ZN(g30114), .A1(g29865), .A2(g11447) );
  AND2_X1 AND2_3668( .ZN(g30115), .A1(g29873), .A2(g11450) );
  AND2_X1 AND2_3669( .ZN(g30116), .A1(g29921), .A2(g22236) );
  AND2_X1 AND2_3670( .ZN(g30117), .A1(g29877), .A2(g11465) );
  AND2_X1 AND2_3671( .ZN(g30118), .A1(g29889), .A2(g11468) );
  AND2_X1 AND2_3672( .ZN(g30123), .A1(g30070), .A2(g20641) );
  AND2_X1 AND2_3673( .ZN(g30127), .A1(g30065), .A2(g20719) );
  AND2_X1 AND2_3674( .ZN(g30128), .A1(g30062), .A2(g20722) );
  AND2_X1 AND2_3675( .ZN(g30129), .A1(g30071), .A2(g20725) );
  AND2_X1 AND2_3676( .ZN(g30131), .A1(g30059), .A2(g20749) );
  AND2_X1 AND2_3677( .ZN(g30132), .A1(g30068), .A2(g20776) );
  AND2_X1 AND2_3678( .ZN(g30133), .A1(g30067), .A2(g20799) );
  AND2_X1 AND2_3679( .ZN(g30138), .A1(g30069), .A2(g20816) );
  AND2_X1 AND2_3680( .ZN(g30216), .A1(g30036), .A2(g8921) );
  AND2_X1 AND2_3681( .ZN(g30217), .A1(g30036), .A2(g8955) );
  AND2_X1 AND2_3682( .ZN(g30218), .A1(g30040), .A2(g8961) );
  AND2_X1 AND2_3683( .ZN(g30219), .A1(g30036), .A2(g8980) );
  AND2_X1 AND2_3684( .ZN(g30220), .A1(g30040), .A2(g8987) );
  AND2_X1 AND2_3685( .ZN(g30221), .A1(g30044), .A2(g8993) );
  AND2_X1 AND2_3686( .ZN(g30222), .A1(g30040), .A2(g9010) );
  AND2_X1 AND2_3687( .ZN(g30223), .A1(g30044), .A2(g9016) );
  AND2_X1 AND2_3688( .ZN(g30224), .A1(g30048), .A2(g9022) );
  AND2_X1 AND2_3689( .ZN(g30225), .A1(g30044), .A2(g9035) );
  AND2_X1 AND2_3690( .ZN(g30226), .A1(g30048), .A2(g9041) );
  AND2_X1 AND2_3691( .ZN(g30227), .A1(g30048), .A2(g9058) );
  AND2_X1 AND2_3692( .ZN(g30327), .A1(g30187), .A2(g8321) );
  AND2_X1 AND2_3693( .ZN(g30330), .A1(g30195), .A2(g8333) );
  AND2_X1 AND2_3694( .ZN(g30333), .A1(g30191), .A2(g8341) );
  AND2_X1 AND2_3695( .ZN(g30334), .A1(g30203), .A2(g8347) );
  AND2_X1 AND2_3696( .ZN(g30337), .A1(g30199), .A2(g8354) );
  AND2_X1 AND2_3697( .ZN(g30340), .A1(g30207), .A2(g8372) );
  AND2_X1 AND2_3698( .ZN(g30345), .A1(g30195), .A2(g8388) );
  AND2_X1 AND2_3699( .ZN(g30348), .A1(g30203), .A2(g8400) );
  AND2_X1 AND2_3700( .ZN(g30351), .A1(g30199), .A2(g8408) );
  AND2_X1 AND2_3701( .ZN(g30352), .A1(g30211), .A2(g8414) );
  AND2_X1 AND2_3702( .ZN(g30355), .A1(g30207), .A2(g8421) );
  AND2_X1 AND2_3703( .ZN(g30361), .A1(g30203), .A2(g8440) );
  AND2_X1 AND2_3704( .ZN(g30364), .A1(g30211), .A2(g8452) );
  AND2_X1 AND2_3705( .ZN(g30367), .A1(g30207), .A2(g8460) );
  AND2_X1 AND2_3706( .ZN(g30372), .A1(g8594), .A2(g30228) );
  AND2_X1 AND2_3707( .ZN(g30374), .A1(g30211), .A2(g8475) );
  AND2_X1 AND2_3708( .ZN(g30387), .A1(g30229), .A2(g8888) );
  AND2_X1 AND2_3709( .ZN(g30388), .A1(g30229), .A2(g8918) );
  AND2_X1 AND2_3710( .ZN(g30389), .A1(g30233), .A2(g8928) );
  AND2_X1 AND2_3711( .ZN(g30390), .A1(g30229), .A2(g8952) );
  AND2_X1 AND2_3712( .ZN(g30391), .A1(g30233), .A2(g8958) );
  AND2_X1 AND2_3713( .ZN(g30392), .A1(g30237), .A2(g8968) );
  AND2_X1 AND2_3714( .ZN(g30393), .A1(g30233), .A2(g8984) );
  AND2_X1 AND2_3715( .ZN(g30394), .A1(g30237), .A2(g8990) );
  AND2_X1 AND2_3716( .ZN(g30395), .A1(g30241), .A2(g9000) );
  AND2_X1 AND2_3717( .ZN(g30396), .A1(g30237), .A2(g9013) );
  AND2_X1 AND2_3718( .ZN(g30397), .A1(g30241), .A2(g9019) );
  AND2_X1 AND2_3719( .ZN(g30398), .A1(g30241), .A2(g9038) );
  AND2_X1 AND2_3720( .ZN(g30407), .A1(g30134), .A2(g10991) );
  AND2_X1 AND2_3721( .ZN(g30409), .A1(g30134), .A2(g11025) );
  AND2_X2 AND2_3722( .ZN(g30410), .A1(g30139), .A2(g11028) );
  AND2_X1 AND2_3723( .ZN(g30411), .A1(g30143), .A2(g11039) );
  AND2_X1 AND2_3724( .ZN(g30436), .A1(g30134), .A2(g11079) );
  AND2_X1 AND2_3725( .ZN(g30437), .A1(g30139), .A2(g11082) );
  AND2_X1 AND2_3726( .ZN(g30438), .A1(g30147), .A2(g11085) );
  AND2_X1 AND2_3727( .ZN(g30440), .A1(g30143), .A2(g11095) );
  AND2_X1 AND2_3728( .ZN(g30441), .A1(g30151), .A2(g11098) );
  AND2_X1 AND2_3729( .ZN(g30442), .A1(g30155), .A2(g11111) );
  AND2_X1 AND2_3730( .ZN(g30444), .A1(g30139), .A2(g11132) );
  AND2_X1 AND2_3731( .ZN(g30445), .A1(g30147), .A2(g11135) );
  AND2_X1 AND2_3732( .ZN(g30447), .A1(g30143), .A2(g11145) );
  AND2_X1 AND2_3733( .ZN(g30448), .A1(g30151), .A2(g11148) );
  AND2_X1 AND2_3734( .ZN(g30449), .A1(g30159), .A2(g11151) );
  AND2_X1 AND2_3735( .ZN(g30451), .A1(g30155), .A2(g11163) );
  AND2_X1 AND2_3736( .ZN(g30452), .A1(g30163), .A2(g11166) );
  AND2_X1 AND2_3737( .ZN(g30453), .A1(g30167), .A2(g11179) );
  AND2_X1 AND2_3738( .ZN(g30454), .A1(g30147), .A2(g11199) );
  AND2_X1 AND2_3739( .ZN(g30457), .A1(g30151), .A2(g11216) );
  AND2_X1 AND2_3740( .ZN(g30458), .A1(g30159), .A2(g11219) );
  AND2_X1 AND2_3741( .ZN(g30460), .A1(g30155), .A2(g11231) );
  AND2_X1 AND2_3742( .ZN(g30461), .A1(g30163), .A2(g11234) );
  AND2_X1 AND2_3743( .ZN(g30462), .A1(g30171), .A2(g11237) );
  AND2_X1 AND2_3744( .ZN(g30464), .A1(g30167), .A2(g11249) );
  AND2_X1 AND2_3745( .ZN(g30465), .A1(g30175), .A2(g11252) );
  AND2_X1 AND2_3746( .ZN(g30467), .A1(g30179), .A2(g11274) );
  AND2_X1 AND2_3747( .ZN(g30469), .A1(g30159), .A2(g11281) );
  AND2_X1 AND2_3748( .ZN(g30472), .A1(g30163), .A2(g11300) );
  AND2_X1 AND2_3749( .ZN(g30473), .A1(g30171), .A2(g11303) );
  AND2_X1 AND2_3750( .ZN(g30475), .A1(g30167), .A2(g11315) );
  AND2_X1 AND2_3751( .ZN(g30476), .A1(g30175), .A2(g11318) );
  AND2_X1 AND2_3752( .ZN(g30477), .A1(g30183), .A2(g11321) );
  AND2_X1 AND2_3753( .ZN(g30478), .A1(g30187), .A2(g11344) );
  AND2_X1 AND2_3754( .ZN(g30481), .A1(g30179), .A2(g11351) );
  AND2_X1 AND2_3755( .ZN(g30484), .A1(g30191), .A2(g11367) );
  AND2_X1 AND2_3756( .ZN(g30486), .A1(g30171), .A2(g11376) );
  AND2_X1 AND2_3757( .ZN(g30489), .A1(g30175), .A2(g11395) );
  AND2_X1 AND2_3758( .ZN(g30490), .A1(g30183), .A2(g11398) );
  AND2_X1 AND2_3759( .ZN(g30492), .A1(g30187), .A2(g11414) );
  AND2_X1 AND2_3760( .ZN(g30495), .A1(g30179), .A2(g11422) );
  AND2_X1 AND2_3761( .ZN(g30496), .A1(g30195), .A2(g11428) );
  AND2_X1 AND2_3762( .ZN(g30499), .A1(g30191), .A2(g11435) );
  AND2_X1 AND2_3763( .ZN(g30502), .A1(g30199), .A2(g11453) );
  AND2_X1 AND2_3764( .ZN(g30504), .A1(g30183), .A2(g11462) );
  AND2_X1 AND2_3765( .ZN(g30696), .A1(g30383), .A2(g10943) );
  AND2_X1 AND2_3766( .ZN(g30697), .A1(g30383), .A2(g11011) );
  AND2_X1 AND2_3767( .ZN(g30698), .A1(g30383), .A2(g11126) );
  AND2_X1 AND2_3768( .ZN(g30728), .A1(g30605), .A2(g22252) );
  AND2_X1 AND2_3769( .ZN(g30735), .A1(g30629), .A2(g22268) );
  AND2_X1 AND2_3770( .ZN(g30736), .A1(g30584), .A2(g20669) );
  AND2_X1 AND2_3771( .ZN(g30743), .A1(g30610), .A2(g22283) );
  AND2_X1 AND2_3772( .ZN(g30744), .A1(g30609), .A2(g20697) );
  AND2_X1 AND2_3773( .ZN(g30750), .A1(g30593), .A2(g20729) );
  AND2_X1 AND2_3774( .ZN(g30754), .A1(g30614), .A2(g22313) );
  AND2_X1 AND2_3775( .ZN(g30755), .A1(g30632), .A2(g22314) );
  AND2_X1 AND2_3776( .ZN(g30757), .A1(g30601), .A2(g20780) );
  AND2_X1 AND2_3777( .ZN(g30758), .A1(g30613), .A2(g20783) );
  AND2_X1 AND2_3778( .ZN(g30759), .A1(g30588), .A2(g22360) );
  AND2_X1 AND2_3779( .ZN(g30760), .A1(g30622), .A2(g22379) );
  AND2_X1 AND2_3780( .ZN(g30761), .A1(g30621), .A2(g20822) );
  AND2_X1 AND2_3781( .ZN(g30762), .A1(g30608), .A2(g20830) );
  AND2_X1 AND2_3782( .ZN(g30763), .A1(g30597), .A2(g22386) );
  AND2_X1 AND2_3783( .ZN(g30764), .A1(g30628), .A2(g20837) );
  AND3_X1 AND3_257( .ZN(g30766), .A1(g30617), .A2(g19457), .A3(g19431) );
  AND2_X1 AND2_3784( .ZN(g30916), .A1(g30785), .A2(g22251) );
  AND2_X1 AND2_3785( .ZN(g30917), .A1(g12446), .A2(g30766) );
  AND2_X1 AND2_3786( .ZN(g30918), .A1(g30780), .A2(g22296) );
  AND2_X1 AND2_3787( .ZN(g30919), .A1(g30786), .A2(g22297) );
  AND2_X1 AND2_3788( .ZN(g30920), .A1(g30787), .A2(g22298) );
  AND2_X1 AND2_3789( .ZN(g30921), .A1(g10773), .A2(g30791) );
  AND2_X1 AND2_3790( .ZN(g30922), .A1(g30788), .A2(g22315) );
  AND2_X1 AND2_3791( .ZN(g30923), .A1(g30789), .A2(g22338) );
  AND2_X1 AND2_3792( .ZN(g30924), .A1(g30783), .A2(g22359) );
  AND2_X1 AND2_3793( .ZN(g30925), .A1(g30790), .A2(g22380) );
  AND2_X1 AND2_3794( .ZN(g30944), .A1(g30935), .A2(g20666) );
  AND2_X1 AND2_3795( .ZN(g30945), .A1(g30931), .A2(g20754) );
  AND2_X1 AND2_3796( .ZN(g30946), .A1(g30930), .A2(g20757) );
  AND2_X1 AND2_3797( .ZN(g30947), .A1(g30936), .A2(g20760) );
  AND2_X1 AND2_3798( .ZN(g30948), .A1(g30929), .A2(g20786) );
  AND2_X1 AND2_3799( .ZN(g30949), .A1(g30933), .A2(g20806) );
  AND2_X1 AND2_3800( .ZN(g30950), .A1(g30932), .A2(g20819) );
  AND2_X2 AND2_3801( .ZN(g30951), .A1(g30934), .A2(g20833) );
  AND2_X1 AND2_3802( .ZN(g30953), .A1(g8605), .A2(g30952) );
  OR2_X1 OR2_0( .ZN(g9144), .A1(g2986), .A2(g5389) );
  OR2_X1 OR2_1( .ZN(g10778), .A1(g2929), .A2(g8022) );
  OR2_X1 OR2_2( .ZN(g12377), .A1(g7553), .A2(g11059) );
  OR2_X1 OR2_3( .ZN(g12407), .A1(g7573), .A2(g10779) );
  OR2_X1 OR2_4( .ZN(g12886), .A1(g9534), .A2(g3398) );
  OR2_X1 OR2_5( .ZN(g12926), .A1(g9676), .A2(g3554) );
  OR2_X1 OR2_6( .ZN(g12955), .A1(g9822), .A2(g3710) );
  OR2_X1 OR2_7( .ZN(g12984), .A1(g9968), .A2(g3866) );
  OR2_X1 OR2_8( .ZN(g16539), .A1(g15880), .A2(g14657) );
  OR2_X1 OR2_9( .ZN(g16571), .A1(g15913), .A2(g14691) );
  OR2_X1 OR2_10( .ZN(g16595), .A1(g15942), .A2(g14725) );
  OR2_X1 OR2_11( .ZN(g16615), .A1(g15971), .A2(g14753) );
  OR2_X1 OR2_12( .ZN(g17973), .A1(g11623), .A2(g15659) );
  OR2_X1 OR2_13( .ZN(g19181), .A1(g17729), .A2(g17979) );
  OR2_X1 OR2_14( .ZN(g19186), .A1(g18419), .A2(g17887) );
  OR2_X1 OR2_15( .ZN(g19187), .A1(g18419), .A2(g17729) );
  OR2_X1 OR2_16( .ZN(g19188), .A1(g17830), .A2(g18096) );
  OR2_X1 OR2_17( .ZN(g19191), .A1(g17807), .A2(g17887) );
  OR2_X1 OR2_18( .ZN(g19192), .A1(g18183), .A2(g18270) );
  OR2_X1 OR2_19( .ZN(g19193), .A1(g18492), .A2(g17998) );
  OR2_X1 OR2_20( .ZN(g19194), .A1(g18492), .A2(g17830) );
  OR2_X1 OR2_21( .ZN(g19195), .A1(g17942), .A2(g18212) );
  OR2_X1 OR2_22( .ZN(g19200), .A1(g18346), .A2(g18424) );
  OR2_X1 OR2_23( .ZN(g19201), .A1(g18183), .A2(g18424) );
  OR2_X1 OR2_24( .ZN(g19202), .A1(g17919), .A2(g17998) );
  OR2_X1 OR2_25( .ZN(g19203), .A1(g18290), .A2(g18363) );
  OR2_X1 OR2_26( .ZN(g19204), .A1(g18556), .A2(g18115) );
  OR2_X1 OR2_27( .ZN(g19205), .A1(g18556), .A2(g17942) );
  OR2_X1 OR2_28( .ZN(g19206), .A1(g18053), .A2(g18319) );
  OR2_X1 OR2_29( .ZN(g19209), .A1(g18079), .A2(g18346) );
  OR2_X1 OR2_30( .ZN(g19210), .A1(g18079), .A2(g18183) );
  OR2_X1 OR2_31( .ZN(g19211), .A1(g18441), .A2(g18497) );
  OR2_X1 OR2_32( .ZN(g19212), .A1(g18290), .A2(g18497) );
  OR2_X2 OR2_33( .ZN(g19213), .A1(g18030), .A2(g18115) );
  OR2_X2 OR2_34( .ZN(g19214), .A1(g18383), .A2(g18458) );
  OR2_X1 OR2_35( .ZN(g19215), .A1(g18606), .A2(g18231) );
  OR2_X1 OR2_36( .ZN(g19216), .A1(g18606), .A2(g18053) );
  OR2_X1 OR2_37( .ZN(g19221), .A1(g18270), .A2(g18346) );
  OR2_X1 OR2_38( .ZN(g19222), .A1(g18195), .A2(g18441) );
  OR2_X1 OR2_39( .ZN(g19223), .A1(g18195), .A2(g18290) );
  OR2_X1 OR2_40( .ZN(g19224), .A1(g18514), .A2(g18561) );
  OR2_X1 OR2_41( .ZN(g19225), .A1(g18383), .A2(g18561) );
  OR2_X1 OR2_42( .ZN(g19226), .A1(g18147), .A2(g18231) );
  OR2_X1 OR2_43( .ZN(g19227), .A1(g18478), .A2(g18531) );
  OR3_X1 OR3_0( .ZN(II25477), .A1(g17024), .A2(g17000), .A3(g16992) );
  OR3_X1 OR3_1( .ZN(g19230), .A1(g16985), .A2(g16965), .A3(II25477) );
  OR2_X1 OR2_44( .ZN(g19231), .A1(g18363), .A2(g18441) );
  OR2_X1 OR2_45( .ZN(g19232), .A1(g18302), .A2(g18514) );
  OR2_X1 OR2_46( .ZN(g19233), .A1(g18302), .A2(g18383) );
  OR2_X1 OR2_47( .ZN(g19234), .A1(g18578), .A2(g18611) );
  OR2_X1 OR2_48( .ZN(g19235), .A1(g18478), .A2(g18611) );
  OR3_X1 OR3_2( .ZN(II25495), .A1(g17158), .A2(g17137), .A3(g17115) );
  OR3_X1 OR3_3( .ZN(g19240), .A1(g17083), .A2(g17050), .A3(II25495) );
  OR2_X1 OR2_49( .ZN(g19242), .A1(g14244), .A2(g16501) );
  OR3_X1 OR3_4( .ZN(II25500), .A1(g17058), .A2(g17030), .A3(g17016) );
  OR3_X1 OR3_5( .ZN(g19243), .A1(g16995), .A2(g16986), .A3(II25500) );
  OR2_X1 OR2_50( .ZN(g19244), .A1(g18458), .A2(g18514) );
  OR2_X1 OR2_51( .ZN(g19245), .A1(g18395), .A2(g18578) );
  OR2_X1 OR2_52( .ZN(g19246), .A1(g18395), .A2(g18478) );
  OR2_X1 OR2_53( .ZN(g19250), .A1(g17729), .A2(g17807) );
  OR3_X1 OR3_6( .ZN(II25516), .A1(g17173), .A2(g17160), .A3(g17142) );
  OR3_X1 OR3_7( .ZN(g19253), .A1(g17121), .A2(g17085), .A3(II25516) );
  OR2_X1 OR2_54( .ZN(g19255), .A1(g14366), .A2(g16523) );
  OR3_X1 OR3_8( .ZN(II25521), .A1(g17093), .A2(g17064), .A3(g17046) );
  OR3_X1 OR3_9( .ZN(g19256), .A1(g17019), .A2(g16996), .A3(II25521) );
  OR2_X1 OR2_55( .ZN(g19257), .A1(g18531), .A2(g18578) );
  OR2_X1 OR2_56( .ZN(g19263), .A1(g17887), .A2(g17979) );
  OR2_X1 OR2_57( .ZN(g19264), .A1(g17830), .A2(g17919) );
  OR3_X1 OR3_10( .ZN(II25549), .A1(g17190), .A2(g17175), .A3(g17165) );
  OR3_X1 OR3_11( .ZN(g19266), .A1(g17148), .A2(g17123), .A3(II25549) );
  OR2_X1 OR2_58( .ZN(g19268), .A1(g14478), .A2(g16554) );
  OR3_X1 OR3_12( .ZN(II25554), .A1(g17131), .A2(g17099), .A3(g17080) );
  OR3_X1 OR3_13( .ZN(g19269), .A1(g17049), .A2(g17020), .A3(II25554) );
  OR3_X1 OR3_14( .ZN(g19275), .A1(g16867), .A2(g16515), .A3(g19001) );
  OR2_X1 OR2_59( .ZN(g19278), .A1(g17998), .A2(g18096) );
  OR2_X1 OR2_60( .ZN(g19279), .A1(g17942), .A2(g18030) );
  OR3_X1 OR3_15( .ZN(II25588), .A1(g17201), .A2(g17192), .A3(g17180) );
  OR3_X1 OR3_16( .ZN(g19281), .A1(g17171), .A2(g17150), .A3(II25588) );
  OR2_X1 OR2_61( .ZN(g19283), .A1(g14565), .A2(g16586) );
  OR3_X1 OR3_17( .ZN(g19294), .A1(g16895), .A2(g16546), .A3(g16507) );
  OR2_X1 OR2_62( .ZN(g19297), .A1(g18115), .A2(g18212) );
  OR2_X1 OR2_63( .ZN(g19298), .A1(g18053), .A2(g18147) );
  OR3_X1 OR3_18( .ZN(g19312), .A1(g16924), .A2(g16578), .A3(g16529) );
  OR2_X1 OR2_64( .ZN(g19315), .A1(g18231), .A2(g18319) );
  OR3_X1 OR3_19( .ZN(g19333), .A1(g16954), .A2(g16602), .A3(g16560) );
  OR2_X1 OR2_65( .ZN(g19450), .A1(g14837), .A2(g16682) );
  OR2_X1 OR2_66( .ZN(g19477), .A1(g14910), .A2(g16708) );
  OR2_X1 OR2_67( .ZN(g19500), .A1(g14991), .A2(g16739) );
  OR3_X1 OR3_20( .ZN(g19503), .A1(g16884), .A2(g16697), .A3(g16665) );
  OR2_X1 OR2_68( .ZN(g19521), .A1(g15080), .A2(g16781) );
  OR3_X1 OR3_21( .ZN(g19522), .A1(g16913), .A2(g16728), .A3(g16686) );
  OR3_X1 OR3_22( .ZN(g19532), .A1(g16943), .A2(g16770), .A3(g16712) );
  OR3_X1 OR3_23( .ZN(g19542), .A1(g16974), .A2(g16797), .A3(g16743) );
  OR3_X1 OR3_24( .ZN(II26429), .A1(g17979), .A2(g17887), .A3(g17807) );
  OR3_X1 OR3_25( .ZN(g19981), .A1(g17729), .A2(g18419), .A3(II26429) );
  OR3_X1 OR3_26( .ZN(II26455), .A1(g18424), .A2(g18346), .A3(g18270) );
  OR3_X1 OR3_27( .ZN(g20015), .A1(g18183), .A2(g18079), .A3(II26455) );
  OR3_X1 OR3_28( .ZN(II26461), .A1(g18096), .A2(g17998), .A3(g17919) );
  OR3_X1 OR3_29( .ZN(g20019), .A1(g17830), .A2(g18492), .A3(II26461) );
  OR3_X1 OR3_30( .ZN(II26491), .A1(g18497), .A2(g18441), .A3(g18363) );
  OR3_X1 OR3_31( .ZN(g20057), .A1(g18290), .A2(g18195), .A3(II26491) );
  OR3_X1 OR3_32( .ZN(II26497), .A1(g18212), .A2(g18115), .A3(g18030) );
  OR3_X1 OR3_33( .ZN(g20061), .A1(g17942), .A2(g18556), .A3(II26497) );
  OR3_X1 OR3_34( .ZN(II26532), .A1(g18561), .A2(g18514), .A3(g18458) );
  OR3_X1 OR3_35( .ZN(g20098), .A1(g18383), .A2(g18302), .A3(II26532) );
  OR3_X1 OR3_36( .ZN(II26538), .A1(g18319), .A2(g18231), .A3(g18147) );
  OR3_X1 OR3_37( .ZN(g20102), .A1(g18053), .A2(g18606), .A3(II26538) );
  OR3_X1 OR3_38( .ZN(II26571), .A1(g18611), .A2(g18578), .A3(g18531) );
  OR3_X1 OR3_39( .ZN(g20123), .A1(g18478), .A2(g18395), .A3(II26571) );
  OR3_X1 OR3_40( .ZN(g21120), .A1(g19484), .A2(g16515), .A3(g14071) );
  OR3_X1 OR3_41( .ZN(g21139), .A1(g19505), .A2(g16546), .A3(g14186) );
  OR3_X1 OR3_42( .ZN(g21159), .A1(g19524), .A2(g16578), .A3(g14301) );
  OR3_X1 OR3_43( .ZN(g21179), .A1(g19534), .A2(g16602), .A3(g14423) );
  OR3_X1 OR3_44( .ZN(g21244), .A1(g19578), .A2(g16697), .A3(g14776) );
  OR3_X1 OR3_45( .ZN(g21253), .A1(g19608), .A2(g16728), .A3(g14811) );
  OR3_X1 OR3_46( .ZN(g21261), .A1(g19641), .A2(g16770), .A3(g14863) );
  OR3_X1 OR3_47( .ZN(g21269), .A1(g19681), .A2(g16797), .A3(g14936) );
  OR3_X1 OR3_48( .ZN(g21501), .A1(g20522), .A2(g16867), .A3(g14071) );
  OR3_X1 OR3_49( .ZN(g21536), .A1(g20522), .A2(g19484), .A3(g19001) );
  OR3_X1 OR3_50( .ZN(g21540), .A1(g20542), .A2(g16895), .A3(g14186) );
  OR3_X1 OR3_51( .ZN(g21572), .A1(g20542), .A2(g19505), .A3(g16507) );
  OR3_X1 OR3_52( .ZN(g21576), .A1(g19067), .A2(g16924), .A3(g14301) );
  OR3_X1 OR3_53( .ZN(g21605), .A1(g19067), .A2(g19524), .A3(g16529) );
  OR3_X1 OR3_54( .ZN(g21609), .A1(g19084), .A2(g16954), .A3(g14423) );
  OR3_X1 OR3_55( .ZN(g21634), .A1(g19084), .A2(g19534), .A3(g16560) );
  OR3_X1 OR3_56( .ZN(g21774), .A1(g19121), .A2(g16884), .A3(g14776) );
  OR3_X1 OR3_57( .ZN(g21787), .A1(g19121), .A2(g19578), .A3(g16665) );
  OR3_X1 OR3_58( .ZN(II28305), .A1(g20197), .A2(g20177), .A3(g20145) );
  OR3_X1 OR3_59( .ZN(g21788), .A1(g20117), .A2(g20094), .A3(II28305) );
  OR3_X1 OR3_60( .ZN(g21789), .A1(g19128), .A2(g16913), .A3(g14811) );
  OR3_X1 OR3_61( .ZN(II28318), .A1(g19092), .A2(g19088), .A3(g19079) );
  OR4_X1 OR4_0( .ZN(g21799), .A1(g16505), .A2(g20538), .A3(g18994), .A4(II28318) );
  OR4_X1 OR4_1( .ZN(g21800), .A1(g18665), .A2(g20270), .A3(g20248), .A4(g18647) );
  OR3_X1 OR3_62( .ZN(g21801), .A1(g19128), .A2(g19608), .A3(g16686) );
  OR3_X1 OR3_63( .ZN(II28323), .A1(g20227), .A2(g20211), .A3(g20183) );
  OR3_X1 OR3_64( .ZN(g21802), .A1(g20147), .A2(g20119), .A3(II28323) );
  OR3_X1 OR3_65( .ZN(g21803), .A1(g19135), .A2(g16943), .A3(g14863) );
  OR4_X1 OR4_2( .ZN(g21806), .A1(g20116), .A2(g20093), .A3(g18547), .A4(g19097) );
  OR3_X1 OR3_66( .ZN(II28330), .A1(g19099), .A2(g19094), .A3(g19089) );
  OR4_X1 OR4_3( .ZN(g21807), .A1(g16527), .A2(g19063), .A3(g19007), .A4(II28330) );
  OR4_X1 OR4_4( .ZN(g21808), .A1(g18688), .A2(g20282), .A3(g20271), .A4(g18650) );
  OR3_X1 OR3_67( .ZN(g21809), .A1(g19135), .A2(g19641), .A3(g16712) );
  OR3_X1 OR3_68( .ZN(II28335), .A1(g20254), .A2(g20241), .A3(g20217) );
  OR3_X1 OR3_69( .ZN(g21810), .A1(g20185), .A2(g20149), .A3(II28335) );
  OR3_X1 OR3_70( .ZN(g21811), .A1(g19138), .A2(g16974), .A3(g14936) );
  OR4_X1 OR4_5( .ZN(g21813), .A1(g20146), .A2(g20118), .A3(g18597), .A4(g19104) );
  OR3_X1 OR3_71( .ZN(II28341), .A1(g19106), .A2(g19101), .A3(g19095) );
  OR4_X1 OR4_6( .ZN(g21814), .A1(g16558), .A2(g19080), .A3(g16513), .A4(II28341) );
  OR4_X1 OR4_7( .ZN(g21815), .A1(g18717), .A2(g20293), .A3(g20283), .A4(g18654) );
  OR3_X1 OR3_72( .ZN(g21816), .A1(g19138), .A2(g19681), .A3(g16743) );
  OR3_X1 OR3_73( .ZN(II28346), .A1(g20277), .A2(g20268), .A3(g20247) );
  OR3_X1 OR3_74( .ZN(g21817), .A1(g20219), .A2(g20187), .A3(II28346) );
  OR4_X1 OR4_8( .ZN(g21819), .A1(g20184), .A2(g20148), .A3(g18629), .A4(g19109) );
  OR3_X1 OR3_75( .ZN(II28351), .A1(g19111), .A2(g19108), .A3(g19102) );
  OR4_X1 OR4_9( .ZN(g21820), .A1(g16590), .A2(g19090), .A3(g16535), .A4(II28351) );
  OR4_X1 OR4_10( .ZN(g21821), .A1(g18753), .A2(g20309), .A3(g20294), .A4(g18668) );
  OR4_X1 OR4_11( .ZN(g21823), .A1(g20218), .A2(g20186), .A3(g18638), .A4(g19116) );
  OR3_X1 OR3_76( .ZN(II28365), .A1(g20280), .A2(g18652), .A3(g18649) );
  OR3_X1 OR3_77( .ZN(g21844), .A1(g20222), .A2(g18645), .A3(II28365) );
  OR3_X1 OR3_78( .ZN(II28369), .A1(g20291), .A2(g18666), .A3(g18653) );
  OR3_X1 OR3_79( .ZN(g21846), .A1(g20249), .A2(g18648), .A3(II28369) );
  OR3_X1 OR3_80( .ZN(II28374), .A1(g20307), .A2(g18689), .A3(g18667) );
  OR3_X1 OR3_81( .ZN(g21849), .A1(g20272), .A2(g18651), .A3(II28374) );
  OR3_X1 OR3_82( .ZN(II28380), .A1(g20326), .A2(g18718), .A3(g18690) );
  OR3_X1 OR3_83( .ZN(g21856), .A1(g20284), .A2(g18655), .A3(II28380) );
  OR2_X2 OR2_69( .ZN(g22175), .A1(g16075), .A2(g20842) );
  OR2_X2 OR2_70( .ZN(g22190), .A1(g16113), .A2(g20850) );
  OR2_X2 OR2_71( .ZN(g22199), .A1(g16164), .A2(g20858) );
  OR2_X1 OR2_72( .ZN(g22205), .A1(g16223), .A2(g20866) );
  OR4_X1 OR4_12( .ZN(g22811), .A1(g562), .A2(g559), .A3(g12451), .A4(g21851) );
  OR3_X1 OR3_84( .ZN(g23052), .A1(g21800), .A2(g21788), .A3(g21844) );
  OR3_X1 OR3_85( .ZN(g23071), .A1(g21808), .A2(g21802), .A3(g21846) );
  OR3_X1 OR3_86( .ZN(g23084), .A1(g21815), .A2(g21810), .A3(g21849) );
  OR2_X1 OR2_73( .ZN(g23089), .A1(g21806), .A2(g21799) );
  OR3_X1 OR3_87( .ZN(g23100), .A1(g21821), .A2(g21817), .A3(g21856) );
  OR2_X1 OR2_74( .ZN(g23107), .A1(g21813), .A2(g21807) );
  OR2_X1 OR2_75( .ZN(g23120), .A1(g21819), .A2(g21814) );
  OR2_X1 OR2_76( .ZN(g23129), .A1(g21823), .A2(g21820) );
  OR2_X1 OR2_77( .ZN(g23319), .A1(g14493), .A2(g22385) );
  OR2_X1 OR2_78( .ZN(g23688), .A1(g23106), .A2(g21906) );
  OR2_X1 OR2_79( .ZN(g23742), .A1(g23119), .A2(g21920) );
  OR2_X1 OR2_80( .ZN(g23797), .A1(g23128), .A2(g21938) );
  OR2_X1 OR2_81( .ZN(g23850), .A1(g23139), .A2(g20647) );
  OR2_X1 OR2_82( .ZN(g23919), .A1(g22666), .A2(g23140) );
  OR2_X1 OR2_83( .ZN(g24239), .A1(g19387), .A2(g22401) );
  OR2_X1 OR2_84( .ZN(g24244), .A1(g14144), .A2(g22317) );
  OR2_X1 OR2_85( .ZN(g24245), .A1(g19417), .A2(g22402) );
  OR2_X1 OR2_86( .ZN(g24252), .A1(g14259), .A2(g22342) );
  OR2_X1 OR2_87( .ZN(g24254), .A1(g19454), .A2(g22403) );
  OR2_X1 OR2_88( .ZN(g24257), .A1(g14381), .A2(g22365) );
  OR2_X1 OR2_89( .ZN(g24258), .A1(g19481), .A2(g22404) );
  OR2_X1 OR2_90( .ZN(g24633), .A1(g24094), .A2(g20842) );
  OR2_X1 OR2_91( .ZN(g24653), .A1(g24095), .A2(g20850) );
  OR2_X1 OR2_92( .ZN(g24672), .A1(g24097), .A2(g20858) );
  OR2_X1 OR2_93( .ZN(g24691), .A1(g24103), .A2(g20866) );
  OR2_X1 OR2_94( .ZN(g24890), .A1(g23639), .A2(g23144) );
  OR2_X1 OR2_95( .ZN(g24909), .A1(g23726), .A2(g23142) );
  OR2_X1 OR2_96( .ZN(g24925), .A1(g23772), .A2(g23141) );
  OR2_X1 OR2_97( .ZN(g24965), .A1(g23922), .A2(g23945) );
  OR2_X1 OR2_98( .ZN(g24978), .A1(g23954), .A2(g23974) );
  OR2_X1 OR2_99( .ZN(g24989), .A1(g23983), .A2(g24004) );
  OR2_X1 OR2_100( .ZN(g25000), .A1(g24013), .A2(g24038) );
  OR2_X1 OR2_101( .ZN(g25183), .A1(g24958), .A2(g24893) );
  OR2_X1 OR2_102( .ZN(g25186), .A1(g24969), .A2(g24916) );
  OR2_X1 OR2_103( .ZN(g25190), .A1(g24982), .A2(g24933) );
  OR2_X1 OR2_104( .ZN(g25195), .A1(g24993), .A2(g24945) );
  OR2_X1 OR2_105( .ZN(g25489), .A1(g24795), .A2(g16466) );
  OR2_X1 OR2_106( .ZN(g25490), .A1(g24759), .A2(g23146) );
  OR2_X1 OR2_107( .ZN(g25520), .A1(g24813), .A2(g23145) );
  OR2_X1 OR2_108( .ZN(g25566), .A1(g24843), .A2(g23143) );
  OR2_X1 OR2_109( .ZN(g26320), .A1(g25852), .A2(g25870) );
  OR2_X1 OR2_110( .ZN(g26367), .A1(g25873), .A2(g25882) );
  OR2_X1 OR2_111( .ZN(g26410), .A1(g25885), .A2(g25887) );
  OR2_X1 OR2_112( .ZN(g26451), .A1(g25890), .A2(g25892) );
  OR2_X1 OR2_113( .ZN(g26974), .A1(g26157), .A2(g23147) );
  OR3_X1 OR3_88( .ZN(g27113), .A1(g1248), .A2(g1245), .A3(g26534) );
  OR2_X1 OR2_114( .ZN(g28501), .A1(g27738), .A2(g25764) );
  OR2_X1 OR2_115( .ZN(g28512), .A1(g26481), .A2(g27738) );
  OR2_X1 OR2_116( .ZN(g28529), .A1(g27743), .A2(g25818) );
  OR2_X1 OR2_117( .ZN(g28540), .A1(g26497), .A2(g27743) );
  OR2_X1 OR2_118( .ZN(g28556), .A1(g27751), .A2(g25853) );
  OR2_X2 OR2_119( .ZN(g28567), .A1(g26512), .A2(g27751) );
  OR2_X2 OR2_120( .ZN(g28584), .A1(g27756), .A2(g25874) );
  OR2_X2 OR2_121( .ZN(g28595), .A1(g26520), .A2(g27756) );
  OR3_X2 OR3_89( .ZN(g29348), .A1(g1942), .A2(g1939), .A3(g29113) );
  OR3_X2 OR3_90( .ZN(g30305), .A1(g2636), .A2(g2633), .A3(g30072) );
  NAND2_X1 NAND2_0( .ZN(II15167), .A1(g2981), .A2(g2874) );
  NAND2_X1 NAND2_1( .ZN(II15168), .A1(g2981), .A2(II15167) );
  NAND2_X1 NAND2_2( .ZN(II15169), .A1(g2874), .A2(II15167) );
  NAND2_X1 NAND2_3( .ZN(g7855), .A1(II15168), .A2(II15169) );
  NAND2_X1 NAND2_4( .ZN(II15183), .A1(g2975), .A2(g2978) );
  NAND2_X1 NAND2_5( .ZN(II15184), .A1(g2975), .A2(II15183) );
  NAND2_X1 NAND2_6( .ZN(II15185), .A1(g2978), .A2(II15183) );
  NAND2_X1 NAND2_7( .ZN(g7875), .A1(II15184), .A2(II15185) );
  NAND2_X1 NAND2_8( .ZN(II15190), .A1(g2956), .A2(g2959) );
  NAND2_X1 NAND2_9( .ZN(II15191), .A1(g2956), .A2(II15190) );
  NAND2_X1 NAND2_10( .ZN(II15192), .A1(g2959), .A2(II15190) );
  NAND2_X1 NAND2_11( .ZN(g7876), .A1(II15191), .A2(II15192) );
  NAND2_X2 NAND2_12( .ZN(II15204), .A1(g2969), .A2(g2972) );
  NAND2_X2 NAND2_13( .ZN(II15205), .A1(g2969), .A2(II15204) );
  NAND2_X1 NAND2_14( .ZN(II15206), .A1(g2972), .A2(II15204) );
  NAND2_X1 NAND2_15( .ZN(g7895), .A1(II15205), .A2(II15206) );
  NAND2_X1 NAND2_16( .ZN(II15211), .A1(g2947), .A2(g2953) );
  NAND2_X1 NAND2_17( .ZN(II15212), .A1(g2947), .A2(II15211) );
  NAND2_X1 NAND2_18( .ZN(II15213), .A1(g2953), .A2(II15211) );
  NAND2_X1 NAND2_19( .ZN(g7896), .A1(II15212), .A2(II15213) );
  NAND2_X1 NAND2_20( .ZN(II15237), .A1(g2963), .A2(g2966) );
  NAND2_X1 NAND2_21( .ZN(II15238), .A1(g2963), .A2(II15237) );
  NAND2_X1 NAND2_22( .ZN(II15239), .A1(g2966), .A2(II15237) );
  NAND2_X1 NAND2_23( .ZN(g7922), .A1(II15238), .A2(II15239) );
  NAND2_X1 NAND2_24( .ZN(II15244), .A1(g2941), .A2(g2944) );
  NAND2_X1 NAND2_25( .ZN(II15245), .A1(g2941), .A2(II15244) );
  NAND2_X1 NAND2_26( .ZN(II15246), .A1(g2944), .A2(II15244) );
  NAND2_X1 NAND2_27( .ZN(g7923), .A1(II15245), .A2(II15246) );
  NAND2_X1 NAND2_28( .ZN(II15276), .A1(g2935), .A2(g2938) );
  NAND2_X1 NAND2_29( .ZN(II15277), .A1(g2935), .A2(II15276) );
  NAND2_X1 NAND2_30( .ZN(II15278), .A1(g2938), .A2(II15276) );
  NAND2_X1 NAND2_31( .ZN(g7970), .A1(II15277), .A2(II15278) );
  NAND4_X1 NAND4_0( .ZN(g8381), .A1(g8182), .A2(g8120), .A3(g8044), .A4(g7989) );
  NAND2_X1 NAND2_32( .ZN(g8533), .A1(g3398), .A2(g3366) );
  NAND2_X1 NAND2_33( .ZN(g8547), .A1(g3398), .A2(g3366) );
  NAND2_X1 NAND2_34( .ZN(g8550), .A1(g3554), .A2(g3522) );
  NAND2_X1 NAND2_35( .ZN(g8560), .A1(g3554), .A2(g3522) );
  NAND2_X1 NAND2_36( .ZN(g8563), .A1(g3710), .A2(g3678) );
  NAND2_X1 NAND2_37( .ZN(g8571), .A1(g3710), .A2(g3678) );
  NAND2_X1 NAND2_38( .ZN(g8574), .A1(g3866), .A2(g3834) );
  NAND2_X1 NAND2_39( .ZN(g8577), .A1(g3866), .A2(g3834) );
  NAND2_X1 NAND2_40( .ZN(II16879), .A1(g4203), .A2(g3998) );
  NAND2_X1 NAND2_41( .ZN(II16880), .A1(g4203), .A2(II16879) );
  NAND2_X1 NAND2_42( .ZN(II16881), .A1(g3998), .A2(II16879) );
  NAND2_X1 NAND2_43( .ZN(g9883), .A1(II16880), .A2(II16881) );
  NAND2_X1 NAND2_44( .ZN(II16965), .A1(g4734), .A2(g4452) );
  NAND2_X1 NAND2_45( .ZN(II16966), .A1(g4734), .A2(II16965) );
  NAND2_X1 NAND2_46( .ZN(II16967), .A1(g4452), .A2(II16965) );
  NAND2_X1 NAND2_47( .ZN(g10003), .A1(II16966), .A2(II16967) );
  NAND2_X1 NAND2_48( .ZN(g10038), .A1(g7772), .A2(g3366) );
  NAND2_X1 NAND2_49( .ZN(II17059), .A1(g6637), .A2(g6309) );
  NAND2_X1 NAND2_50( .ZN(II17060), .A1(g6637), .A2(II17059) );
  NAND2_X1 NAND2_51( .ZN(II17061), .A1(g6309), .A2(II17059) );
  NAND2_X1 NAND2_52( .ZN(g10095), .A1(II17060), .A2(II17061) );
  NAND2_X1 NAND2_53( .ZN(g10147), .A1(g7788), .A2(g3522) );
  NAND2_X1 NAND2_54( .ZN(II17149), .A1(g7465), .A2(g7142) );
  NAND2_X2 NAND2_55( .ZN(II17150), .A1(g7465), .A2(II17149) );
  NAND2_X2 NAND2_56( .ZN(II17151), .A1(g7142), .A2(II17149) );
  NAND2_X1 NAND2_57( .ZN(g10185), .A1(II17150), .A2(II17151) );
  NAND2_X1 NAND2_58( .ZN(g10252), .A1(g7802), .A2(g3678) );
  NAND2_X1 NAND2_59( .ZN(g10354), .A1(g7815), .A2(g3834) );
  NAND2_X1 NAND2_60( .ZN(g10649), .A1(g3398), .A2(g6912) );
  NAND2_X1 NAND2_61( .ZN(g10676), .A1(g3398), .A2(g6678) );
  NAND2_X1 NAND2_62( .ZN(g10677), .A1(g3398), .A2(g6912) );
  NAND2_X1 NAND2_63( .ZN(g10679), .A1(g3554), .A2(g7162) );
  NAND2_X1 NAND2_64( .ZN(g10703), .A1(g3398), .A2(g6678) );
  NAND2_X1 NAND2_65( .ZN(g10705), .A1(g3554), .A2(g6980) );
  NAND2_X1 NAND2_66( .ZN(g10706), .A1(g3554), .A2(g7162) );
  NAND2_X1 NAND2_67( .ZN(g10708), .A1(g3710), .A2(g7358) );
  NAND2_X1 NAND2_68( .ZN(g10723), .A1(g3554), .A2(g6980) );
  NAND2_X1 NAND2_69( .ZN(g10725), .A1(g3710), .A2(g7230) );
  NAND2_X1 NAND2_70( .ZN(g10726), .A1(g3710), .A2(g7358) );
  NAND2_X1 NAND2_71( .ZN(g10728), .A1(g3866), .A2(g7488) );
  NAND2_X1 NAND2_72( .ZN(g10744), .A1(g3710), .A2(g7230) );
  NAND2_X1 NAND2_73( .ZN(g10746), .A1(g3866), .A2(g7426) );
  NAND2_X1 NAND2_74( .ZN(g10747), .A1(g3866), .A2(g7488) );
  NAND2_X1 NAND2_75( .ZN(g10763), .A1(g3866), .A2(g7426) );
  NAND2_X1 NAND2_76( .ZN(II18106), .A1(g7875), .A2(g7855) );
  NAND2_X1 NAND2_77( .ZN(II18107), .A1(g7875), .A2(II18106) );
  NAND2_X1 NAND2_78( .ZN(II18108), .A1(g7855), .A2(II18106) );
  NAND2_X1 NAND2_79( .ZN(g11188), .A1(II18107), .A2(II18108) );
  NAND2_X1 NAND2_80( .ZN(II18113), .A1(g3997), .A2(g8181) );
  NAND2_X1 NAND2_81( .ZN(II18114), .A1(g3997), .A2(II18113) );
  NAND2_X1 NAND2_82( .ZN(II18115), .A1(g8181), .A2(II18113) );
  NAND2_X1 NAND2_83( .ZN(g11189), .A1(II18114), .A2(II18115) );
  NAND2_X1 NAND2_84( .ZN(II18190), .A1(g7922), .A2(g7895) );
  NAND2_X1 NAND2_85( .ZN(II18191), .A1(g7922), .A2(II18190) );
  NAND2_X1 NAND2_86( .ZN(II18192), .A1(g7895), .A2(II18190) );
  NAND2_X1 NAND2_87( .ZN(g11262), .A1(II18191), .A2(II18192) );
  NAND2_X1 NAND2_88( .ZN(II18197), .A1(g7896), .A2(g7876) );
  NAND2_X1 NAND2_89( .ZN(II18198), .A1(g7896), .A2(II18197) );
  NAND2_X1 NAND2_90( .ZN(II18199), .A1(g7876), .A2(II18197) );
  NAND2_X1 NAND2_91( .ZN(g11263), .A1(II18198), .A2(II18199) );
  NAND2_X1 NAND2_92( .ZN(II18204), .A1(g7975), .A2(g4202) );
  NAND2_X1 NAND2_93( .ZN(II18205), .A1(g7975), .A2(II18204) );
  NAND2_X1 NAND2_94( .ZN(II18206), .A1(g4202), .A2(II18204) );
  NAND2_X1 NAND2_95( .ZN(g11264), .A1(II18205), .A2(II18206) );
  NAND2_X1 NAND2_96( .ZN(II18280), .A1(g7970), .A2(g7923) );
  NAND2_X1 NAND2_97( .ZN(II18281), .A1(g7970), .A2(II18280) );
  NAND2_X1 NAND2_98( .ZN(II18282), .A1(g7923), .A2(II18280) );
  NAND2_X1 NAND2_99( .ZN(g11330), .A1(II18281), .A2(II18282) );
  NAND2_X1 NAND2_100( .ZN(II18287), .A1(g8256), .A2(g8102) );
  NAND2_X1 NAND2_101( .ZN(II18288), .A1(g8256), .A2(II18287) );
  NAND2_X1 NAND2_102( .ZN(II18289), .A1(g8102), .A2(II18287) );
  NAND2_X1 NAND2_103( .ZN(g11331), .A1(II18288), .A2(II18289) );
  NAND2_X1 NAND2_104( .ZN(II18368), .A1(g4325), .A2(g4093) );
  NAND2_X1 NAND2_105( .ZN(II18369), .A1(g4325), .A2(II18368) );
  NAND2_X1 NAND2_106( .ZN(II18370), .A1(g4093), .A2(II18368) );
  NAND2_X1 NAND2_107( .ZN(g11410), .A1(II18369), .A2(II18370) );
  NAND2_X1 NAND2_108( .ZN(g11617), .A1(g8313), .A2(g2883) );
  NAND2_X1 NAND2_109( .ZN(II18799), .A1(g11410), .A2(g11331) );
  NAND2_X1 NAND2_110( .ZN(II18800), .A1(g11410), .A2(II18799) );
  NAND2_X1 NAND2_111( .ZN(II18801), .A1(g11331), .A2(II18799) );
  NAND2_X1 NAND2_112( .ZN(g11621), .A1(II18800), .A2(II18801) );
  NAND2_X1 NAND2_113( .ZN(g11661), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_114( .ZN(g11662), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_115( .ZN(g11672), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_116( .ZN(g11673), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_117( .ZN(g11674), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_118( .ZN(g11683), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_119( .ZN(g11684), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_120( .ZN(g11685), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_121( .ZN(g11686), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_122( .ZN(g11691), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_123( .ZN(g11692), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_124( .ZN(g11693), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_125( .ZN(g11694), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_126( .ZN(g11695), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_127( .ZN(g11696), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_128( .ZN(g11698), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_129( .ZN(g11699), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_130( .ZN(g11700), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_131( .ZN(g11701), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_132( .ZN(g11702), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_133( .ZN(g11704), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_134( .ZN(g11705), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_135( .ZN(g11707), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_136( .ZN(g11708), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_137( .ZN(g11709), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_138( .ZN(g11710), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_139( .ZN(g11712), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_140( .ZN(g11713), .A1(g10481), .A2(g9144) );
  NAND2_X1 NAND2_141( .ZN(g11716), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_142( .ZN(g11717), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_143( .ZN(g11718), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_144( .ZN(g11719), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_145( .ZN(g11720), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_146( .ZN(g11721), .A1(g9534), .A2(g3366) );
  NAND2_X1 NAND2_147( .ZN(g11722), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_148( .ZN(g11723), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_149( .ZN(g11724), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_150( .ZN(g11725), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_151( .ZN(g11726), .A1(g9676), .A2(g3522) );
  NAND2_X1 NAND2_152( .ZN(g11727), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_153( .ZN(g11728), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_154( .ZN(g11729), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_155( .ZN(g11730), .A1(g9822), .A2(g3678) );
  NAND2_X1 NAND2_156( .ZN(g11731), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_157( .ZN(g11733), .A1(g9968), .A2(g3834) );
  NAND2_X1 NAND2_158( .ZN(g12433), .A1(g2879), .A2(g10778) );
  NAND2_X1 NAND2_159( .ZN(g12486), .A1(g8278), .A2(g6448) );
  NAND2_X1 NAND2_160( .ZN(g12503), .A1(g8278), .A2(g5438) );
  NAND2_X1 NAND2_161( .ZN(g12506), .A1(g8287), .A2(g6713) );
  NAND2_X1 NAND2_162( .ZN(g12520), .A1(g8287), .A2(g5473) );
  NAND2_X1 NAND2_163( .ZN(g12523), .A1(g8296), .A2(g7015) );
  NAND2_X1 NAND2_164( .ZN(g12535), .A1(g8296), .A2(g5512) );
  NAND2_X2 NAND2_165( .ZN(g12538), .A1(g8305), .A2(g7265) );
  NAND2_X2 NAND2_166( .ZN(g12544), .A1(g8305), .A2(g5556) );
  NAND2_X2 NAND2_167( .ZN(II20031), .A1(g10003), .A2(g9883) );
  NAND2_X1 NAND2_168( .ZN(II20032), .A1(g10003), .A2(II20031) );
  NAND2_X1 NAND2_169( .ZN(II20033), .A1(g9883), .A2(II20031) );
  NAND2_X1 NAND2_170( .ZN(g12988), .A1(II20032), .A2(II20033) );
  NAND2_X1 NAND2_171( .ZN(II20048), .A1(g10185), .A2(g10095) );
  NAND2_X1 NAND2_172( .ZN(II20049), .A1(g10185), .A2(II20048) );
  NAND2_X1 NAND2_173( .ZN(II20050), .A1(g10095), .A2(II20048) );
  NAND2_X1 NAND2_174( .ZN(g12999), .A1(II20049), .A2(II20050) );
  NAND2_X1 NAND2_175( .ZN(g13020), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_176( .ZN(g13021), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_177( .ZN(g13026), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_178( .ZN(g13027), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_179( .ZN(g13028), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_180( .ZN(g13029), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_181( .ZN(g13030), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_182( .ZN(g13034), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_183( .ZN(g13035), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_184( .ZN(g13037), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_185( .ZN(g13038), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_186( .ZN(g13039), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_187( .ZN(g13040), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_188( .ZN(g13041), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_189( .ZN(g13044), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_190( .ZN(g13045), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_191( .ZN(g13047), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_192( .ZN(g13048), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_193( .ZN(g13050), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_194( .ZN(g13051), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_195( .ZN(g13052), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_196( .ZN(g13053), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_197( .ZN(g13054), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_198( .ZN(g13058), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_199( .ZN(g13059), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_200( .ZN(g13061), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_201( .ZN(g13062), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_202( .ZN(g13064), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_203( .ZN(g13065), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_204( .ZN(g13067), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_205( .ZN(g13068), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_206( .ZN(g13069), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_207( .ZN(g13071), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_208( .ZN(g13072), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_209( .ZN(g13074), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_210( .ZN(g13075), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_211( .ZN(g13077), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_212( .ZN(g13078), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_213( .ZN(g13080), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_214( .ZN(g13081), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_215( .ZN(g13087), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_216( .ZN(g13088), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_217( .ZN(g13089), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_218( .ZN(g13090), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_219( .ZN(g13091), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_220( .ZN(g13093), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_221( .ZN(g13094), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_222( .ZN(g13096), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_223( .ZN(g13097), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_224( .ZN(g13098), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_225( .ZN(g13099), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_226( .ZN(g13100), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_227( .ZN(g13102), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_228( .ZN(g13103), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_229( .ZN(g13104), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_230( .ZN(g13105), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_231( .ZN(g13106), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_232( .ZN(g13108), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_233( .ZN(g13109), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_234( .ZN(g13112), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_235( .ZN(g13113), .A1(g9534), .A2(g6912) );
  NAND2_X1 NAND2_236( .ZN(g13114), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_237( .ZN(g13115), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_238( .ZN(g13116), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_239( .ZN(g13118), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_240( .ZN(g13119), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_241( .ZN(g13120), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_242( .ZN(g13121), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_243( .ZN(g13122), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_244( .ZN(g13123), .A1(g9534), .A2(g6678) );
  NAND2_X1 NAND2_245( .ZN(g13125), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_246( .ZN(g13126), .A1(g9676), .A2(g7162) );
  NAND2_X1 NAND2_247( .ZN(g13127), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_248( .ZN(g13128), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_249( .ZN(g13129), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_250( .ZN(g13131), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_251( .ZN(g13132), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_252( .ZN(g13133), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_253( .ZN(g13134), .A1(g9676), .A2(g6980) );
  NAND2_X1 NAND2_254( .ZN(g13136), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_255( .ZN(g13137), .A1(g9822), .A2(g7358) );
  NAND2_X1 NAND2_256( .ZN(g13138), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_257( .ZN(g13139), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_258( .ZN(g13140), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_259( .ZN(g13142), .A1(g9822), .A2(g7230) );
  NAND2_X1 NAND2_260( .ZN(g13144), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_261( .ZN(g13145), .A1(g9968), .A2(g7488) );
  NAND2_X1 NAND2_262( .ZN(g13146), .A1(g9968), .A2(g7426) );
  NAND2_X1 NAND2_263( .ZN(g13147), .A1(g8278), .A2(g3306) );
  NAND2_X1 NAND2_264( .ZN(g13150), .A1(g8287), .A2(g3462) );
  NAND2_X1 NAND2_265( .ZN(g13156), .A1(g8296), .A2(g3618) );
  NAND2_X1 NAND2_266( .ZN(g13165), .A1(g8305), .A2(g3774) );
  NAND2_X1 NAND2_267( .ZN(g13245), .A1(g10779), .A2(g7901) );
  NAND2_X1 NAND2_268( .ZN(g13305), .A1(g8317), .A2(g2993) );
  NAND2_X1 NAND2_269( .ZN(II20429), .A1(g11262), .A2(g11188) );
  NAND2_X1 NAND2_270( .ZN(II20430), .A1(g11262), .A2(II20429) );
  NAND2_X1 NAND2_271( .ZN(II20431), .A1(g11188), .A2(II20429) );
  NAND2_X1 NAND2_272( .ZN(g13348), .A1(II20430), .A2(II20431) );
  NAND2_X1 NAND2_273( .ZN(II20465), .A1(g11330), .A2(g11263) );
  NAND2_X1 NAND2_274( .ZN(II20466), .A1(g11330), .A2(II20465) );
  NAND2_X1 NAND2_275( .ZN(II20467), .A1(g11263), .A2(II20465) );
  NAND2_X1 NAND2_276( .ZN(g13370), .A1(II20466), .A2(II20467) );
  NAND2_X1 NAND2_277( .ZN(II20504), .A1(g11264), .A2(g11189) );
  NAND2_X1 NAND2_278( .ZN(II20505), .A1(g11264), .A2(II20504) );
  NAND2_X1 NAND2_279( .ZN(II20506), .A1(g11189), .A2(II20504) );
  NAND2_X1 NAND2_280( .ZN(g13399), .A1(II20505), .A2(II20506) );
  NAND2_X1 NAND2_281( .ZN(g13476), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_282( .ZN(g13478), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_283( .ZN(g13482), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_284( .ZN(g13494), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_285( .ZN(g13495), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_286( .ZN(g13497), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_287( .ZN(g13501), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_288( .ZN(II20743), .A1(g11621), .A2(g13399) );
  NAND2_X1 NAND2_289( .ZN(II20744), .A1(g11621), .A2(II20743) );
  NAND2_X1 NAND2_290( .ZN(II20745), .A1(g13399), .A2(II20743) );
  NAND2_X1 NAND2_291( .ZN(g13507), .A1(II20744), .A2(II20745) );
  NAND2_X1 NAND2_292( .ZN(g13510), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_293( .ZN(g13511), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_294( .ZN(g13512), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_295( .ZN(g13514), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_296( .ZN(g13518), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_297( .ZN(g13524), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_298( .ZN(g13525), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_299( .ZN(g13526), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_300( .ZN(g13528), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_301( .ZN(g13529), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_302( .ZN(g13535), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_303( .ZN(g13536), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_304( .ZN(g13537), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_305( .ZN(g13538), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_306( .ZN(g13539), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_307( .ZN(g13540), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_308( .ZN(g13546), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_309( .ZN(g13547), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_310( .ZN(g13548), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_311( .ZN(g13549), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_312( .ZN(g13550), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_313( .ZN(g13551), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_314( .ZN(g13557), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_315( .ZN(g13558), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_316( .ZN(g13559), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_317( .ZN(g13560), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_318( .ZN(g13561), .A1(g12657), .A2(g3566) );
  NAND2_X1 NAND2_319( .ZN(g13562), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_320( .ZN(g13563), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_321( .ZN(g13564), .A1(g12711), .A2(g3722) );
  NAND2_X1 NAND2_322( .ZN(g13599), .A1(g12886), .A2(g3366) );
  NAND2_X1 NAND2_323( .ZN(g13611), .A1(g12926), .A2(g3522) );
  NAND2_X1 NAND2_324( .ZN(g13621), .A1(g12955), .A2(g3678) );
  NAND2_X1 NAND2_325( .ZN(g13633), .A1(g12984), .A2(g3834) );
  NAND2_X1 NAND2_326( .ZN(g13893), .A1(g8580), .A2(g12463) );
  NAND3_X1 NAND3_0( .ZN(g13915), .A1(g8822), .A2(g12473), .A3(g12463) );
  NAND2_X1 NAND2_327( .ZN(g13934), .A1(g8587), .A2(g12478) );
  NAND2_X1 NAND2_328( .ZN(g13957), .A1(g10730), .A2(g12473) );
  NAND3_X1 NAND3_1( .ZN(g13971), .A1(g8846), .A2(g12490), .A3(g12478) );
  NAND2_X1 NAND2_329( .ZN(g13990), .A1(g8594), .A2(g12495) );
  NAND2_X1 NAND2_330( .ZN(g14027), .A1(g10749), .A2(g12490) );
  NAND3_X1 NAND3_2( .ZN(g14041), .A1(g8873), .A2(g12510), .A3(g12495) );
  NAND2_X1 NAND2_331( .ZN(g14060), .A1(g8605), .A2(g12515) );
  NAND2_X1 NAND2_332( .ZN(g14118), .A1(g10767), .A2(g12510) );
  NAND3_X1 NAND3_3( .ZN(g14132), .A1(g8911), .A2(g12527), .A3(g12515) );
  NAND2_X1 NAND2_333( .ZN(g14233), .A1(g10773), .A2(g12527) );
  NAND3_X1 NAND3_4( .ZN(g15454), .A1(g9232), .A2(g9150), .A3(g12780) );
  NAND3_X1 NAND3_5( .ZN(g15540), .A1(g9310), .A2(g9174), .A3(g12819) );
  NAND3_X1 NAND3_6( .ZN(g15618), .A1(g9391), .A2(g9216), .A3(g12857) );
  NAND2_X1 NAND2_334( .ZN(g15660), .A1(g13401), .A2(g12354) );
  NAND2_X1 NAND2_335( .ZN(g15664), .A1(g12565), .A2(g6314) );
  NAND3_X1 NAND3_7( .ZN(g15694), .A1(g9488), .A2(g9277), .A3(g12898) );
  NAND2_X1 NAND2_336( .ZN(g15718), .A1(g13286), .A2(g12354) );
  NAND2_X1 NAND2_337( .ZN(g15719), .A1(g13401), .A2(g12392) );
  NAND2_X1 NAND2_338( .ZN(g15720), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_339( .ZN(g15721), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_340( .ZN(g15723), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_341( .ZN(g15756), .A1(g13313), .A2(g12354) );
  NAND2_X1 NAND2_342( .ZN(g15757), .A1(g11622), .A2(g12392) );
  NAND2_X1 NAND2_343( .ZN(g15758), .A1(g12565), .A2(g6232) );
  NAND2_X2 NAND2_344( .ZN(g15759), .A1(g12565), .A2(g6314) );
  NAND2_X2 NAND2_345( .ZN(g15760), .A1(g12611), .A2(g6369) );
  NAND2_X2 NAND2_346( .ZN(g15761), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_347( .ZN(g15763), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_348( .ZN(g15782), .A1(g13332), .A2(g12354) );
  NAND2_X1 NAND2_349( .ZN(g15783), .A1(g11643), .A2(g12392) );
  NAND2_X1 NAND2_350( .ZN(g15784), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_351( .ZN(g15785), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_352( .ZN(g15786), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_353( .ZN(g15787), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_354( .ZN(g15788), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_355( .ZN(g15789), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_356( .ZN(g15791), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_357( .ZN(g15803), .A1(g13375), .A2(g12354) );
  NAND2_X1 NAND2_358( .ZN(g15804), .A1(g11660), .A2(g12392) );
  NAND2_X1 NAND2_359( .ZN(g15805), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_360( .ZN(g15806), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_361( .ZN(g15807), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_362( .ZN(g15808), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_363( .ZN(g15809), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_364( .ZN(g15810), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_365( .ZN(g15811), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_366( .ZN(g15812), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_367( .ZN(II22062), .A1(g12999), .A2(g12988) );
  NAND2_X1 NAND2_368( .ZN(II22063), .A1(g12999), .A2(II22062) );
  NAND2_X1 NAND2_369( .ZN(II22064), .A1(g12988), .A2(II22062) );
  NAND2_X1 NAND2_370( .ZN(g15814), .A1(II22063), .A2(II22064) );
  NAND2_X1 NAND2_371( .ZN(g15818), .A1(g13024), .A2(g12354) );
  NAND2_X1 NAND2_372( .ZN(g15819), .A1(g13286), .A2(g12392) );
  NAND2_X1 NAND2_373( .ZN(g15820), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_374( .ZN(g15821), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_375( .ZN(g15822), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_376( .ZN(g15823), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_377( .ZN(g15824), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_378( .ZN(g15825), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_379( .ZN(g15826), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_380( .ZN(g15827), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_381( .ZN(g15830), .A1(g13310), .A2(g12392) );
  NAND2_X1 NAND2_382( .ZN(g15831), .A1(g13313), .A2(g12392) );
  NAND2_X1 NAND2_383( .ZN(g15832), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_384( .ZN(g15833), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_385( .ZN(g15834), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_386( .ZN(g15835), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_387( .ZN(g15836), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_388( .ZN(g15837), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_389( .ZN(g15838), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_390( .ZN(g15839), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_391( .ZN(g15841), .A1(g13331), .A2(g12392) );
  NAND2_X1 NAND2_392( .ZN(g15842), .A1(g13332), .A2(g12392) );
  NAND2_X1 NAND2_393( .ZN(g15843), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_394( .ZN(g15844), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_395( .ZN(g15845), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_396( .ZN(g15846), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_397( .ZN(g15847), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_398( .ZN(g15848), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_399( .ZN(g15849), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_400( .ZN(g15850), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_401( .ZN(g15851), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_402( .ZN(g15853), .A1(g13310), .A2(g12354) );
  NAND2_X1 NAND2_403( .ZN(g15854), .A1(g13353), .A2(g12392) );
  NAND2_X1 NAND2_404( .ZN(g15855), .A1(g13354), .A2(g12392) );
  NAND2_X1 NAND2_405( .ZN(g15856), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_406( .ZN(g15857), .A1(g12565), .A2(g6314) );
  NAND2_X1 NAND2_407( .ZN(g15858), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_408( .ZN(g15866), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_409( .ZN(g15867), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_410( .ZN(g15868), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_411( .ZN(g15869), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_412( .ZN(g15870), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_413( .ZN(g15871), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_414( .ZN(g15872), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_415( .ZN(g15877), .A1(g13374), .A2(g12392) );
  NAND2_X1 NAND2_416( .ZN(g15878), .A1(g13375), .A2(g12392) );
  NAND2_X1 NAND2_417( .ZN(g15879), .A1(g12565), .A2(g6232) );
  NAND2_X1 NAND2_418( .ZN(g15887), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_419( .ZN(g15888), .A1(g12611), .A2(g6519) );
  NAND2_X1 NAND2_420( .ZN(g15889), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_421( .ZN(g15897), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_422( .ZN(g15898), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_423( .ZN(g15899), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_424( .ZN(g15900), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_425( .ZN(g15901), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_426( .ZN(g15903), .A1(g13404), .A2(g12392) );
  NAND2_X1 NAND2_427( .ZN(g15912), .A1(g12611), .A2(g6369) );
  NAND2_X1 NAND2_428( .ZN(g15920), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_429( .ZN(g15921), .A1(g12657), .A2(g6783) );
  NAND2_X1 NAND2_430( .ZN(g15922), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_431( .ZN(g15930), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_432( .ZN(g15931), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_433( .ZN(g15932), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_434( .ZN(g15941), .A1(g12657), .A2(g6574) );
  NAND2_X1 NAND2_435( .ZN(g15949), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_436( .ZN(g15950), .A1(g12711), .A2(g7085) );
  NAND2_X1 NAND2_437( .ZN(g15951), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_438( .ZN(g15970), .A1(g12711), .A2(g6838) );
  NAND2_X1 NAND2_439( .ZN(g15990), .A1(g12886), .A2(g6912) );
  NAND2_X1 NAND2_440( .ZN(g15992), .A1(g12886), .A2(g6678) );
  NAND2_X1 NAND2_441( .ZN(g15993), .A1(g12926), .A2(g7162) );
  NAND2_X1 NAND2_442( .ZN(g15995), .A1(g12926), .A2(g6980) );
  NAND2_X1 NAND2_443( .ZN(g15996), .A1(g12955), .A2(g7358) );
  NAND2_X1 NAND2_444( .ZN(g15999), .A1(g12955), .A2(g7230) );
  NAND2_X1 NAND2_445( .ZN(g16000), .A1(g12984), .A2(g7488) );
  NAND2_X1 NAND2_446( .ZN(g16006), .A1(g12984), .A2(g7426) );
  NAND2_X1 NAND2_447( .ZN(g16085), .A1(g12883), .A2(g633) );
  NAND2_X1 NAND2_448( .ZN(g16123), .A1(g12923), .A2(g1319) );
  NAND2_X1 NAND2_449( .ZN(II22282), .A1(g2962), .A2(g13348) );
  NAND2_X1 NAND2_450( .ZN(II22283), .A1(g2962), .A2(II22282) );
  NAND2_X1 NAND2_451( .ZN(II22284), .A1(g13348), .A2(II22282) );
  NAND2_X1 NAND2_452( .ZN(g16132), .A1(II22283), .A2(II22284) );
  NAND2_X1 NAND2_453( .ZN(g16174), .A1(g12952), .A2(g2013) );
  NAND2_X1 NAND2_454( .ZN(II22316), .A1(g2934), .A2(g13370) );
  NAND2_X1 NAND2_455( .ZN(II22317), .A1(g2934), .A2(II22316) );
  NAND2_X1 NAND2_456( .ZN(II22318), .A1(g13370), .A2(II22316) );
  NAND2_X1 NAND2_457( .ZN(g16181), .A1(II22317), .A2(II22318) );
  NAND2_X1 NAND2_458( .ZN(g16233), .A1(g12981), .A2(g2707) );
  NAND2_X1 NAND2_459( .ZN(g16341), .A1(g12377), .A2(g12407) );
  NAND2_X1 NAND2_460( .ZN(g16412), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_461( .ZN(g16439), .A1(g13082), .A2(g2912) );
  NAND2_X1 NAND2_462( .ZN(g16442), .A1(g12565), .A2(g3254) );
  NAND2_X1 NAND2_463( .ZN(g16446), .A1(g12611), .A2(g3410) );
  NAND2_X1 NAND2_464( .ZN(g16463), .A1(g13004), .A2(g3018) );
  NAND2_X1 NAND2_465( .ZN(g16536), .A1(g15873), .A2(g2896) );
  NAND2_X1 NAND2_466( .ZN(II22630), .A1(g13507), .A2(g15978) );
  NAND2_X1 NAND2_467( .ZN(II22631), .A1(g13507), .A2(II22630) );
  NAND2_X1 NAND2_468( .ZN(II22632), .A1(g15978), .A2(II22630) );
  NAND2_X1 NAND2_469( .ZN(g16566), .A1(II22631), .A2(II22632) );
  NAND2_X1 NAND2_470( .ZN(II22705), .A1(g13348), .A2(g15661) );
  NAND2_X1 NAND2_471( .ZN(II22706), .A1(g13348), .A2(II22705) );
  NAND2_X1 NAND2_472( .ZN(II22707), .A1(g15661), .A2(II22705) );
  NAND2_X1 NAND2_473( .ZN(g16662), .A1(II22706), .A2(II22707) );
  NAND2_X1 NAND2_474( .ZN(II22884), .A1(g13370), .A2(g15661) );
  NAND2_X1 NAND2_475( .ZN(II22885), .A1(g13370), .A2(II22884) );
  NAND2_X1 NAND2_476( .ZN(II22886), .A1(g15661), .A2(II22884) );
  NAND2_X1 NAND2_477( .ZN(g16935), .A1(II22885), .A2(II22886) );
  NAND2_X1 NAND2_478( .ZN(II22900), .A1(g15022), .A2(g14000) );
  NAND2_X1 NAND2_479( .ZN(II22901), .A1(g15022), .A2(II22900) );
  NAND2_X1 NAND2_480( .ZN(II22902), .A1(g14000), .A2(II22900) );
  NAND2_X1 NAND2_481( .ZN(g16965), .A1(II22901), .A2(II22902) );
  NAND2_X1 NAND2_482( .ZN(II22917), .A1(g15096), .A2(g13945) );
  NAND2_X1 NAND2_483( .ZN(II22918), .A1(g15096), .A2(II22917) );
  NAND2_X1 NAND2_484( .ZN(II22919), .A1(g13945), .A2(II22917) );
  NAND2_X1 NAND2_485( .ZN(g16985), .A1(II22918), .A2(II22919) );
  NAND2_X1 NAND2_486( .ZN(II22924), .A1(g15118), .A2(g14091) );
  NAND2_X1 NAND2_487( .ZN(II22925), .A1(g15118), .A2(II22924) );
  NAND2_X1 NAND2_488( .ZN(II22926), .A1(g14091), .A2(II22924) );
  NAND2_X1 NAND2_489( .ZN(g16986), .A1(II22925), .A2(II22926) );
  NAND2_X1 NAND2_490( .ZN(II22936), .A1(g9150), .A2(g13906) );
  NAND2_X1 NAND2_491( .ZN(II22937), .A1(g9150), .A2(II22936) );
  NAND2_X1 NAND2_492( .ZN(II22938), .A1(g13906), .A2(II22936) );
  NAND2_X1 NAND2_493( .ZN(g16992), .A1(II22937), .A2(II22938) );
  NAND2_X1 NAND2_494( .ZN(II22945), .A1(g15188), .A2(g14015) );
  NAND2_X1 NAND2_495( .ZN(II22946), .A1(g15188), .A2(II22945) );
  NAND2_X1 NAND2_496( .ZN(II22947), .A1(g14015), .A2(II22945) );
  NAND2_X1 NAND2_497( .ZN(g16995), .A1(II22946), .A2(II22947) );
  NAND2_X1 NAND2_498( .ZN(II22952), .A1(g15210), .A2(g14206) );
  NAND2_X1 NAND2_499( .ZN(II22953), .A1(g15210), .A2(II22952) );
  NAND2_X1 NAND2_500( .ZN(II22954), .A1(g14206), .A2(II22952) );
  NAND2_X1 NAND2_501( .ZN(g16996), .A1(II22953), .A2(II22954) );
  NAND2_X1 NAND2_502( .ZN(II22962), .A1(g9161), .A2(g13885) );
  NAND2_X1 NAND2_503( .ZN(II22963), .A1(g9161), .A2(II22962) );
  NAND2_X1 NAND2_504( .ZN(II22964), .A1(g13885), .A2(II22962) );
  NAND2_X1 NAND2_505( .ZN(g17000), .A1(II22963), .A2(II22964) );
  NAND2_X1 NAND2_506( .ZN(II22972), .A1(g9174), .A2(g13962) );
  NAND2_X1 NAND2_507( .ZN(II22973), .A1(g9174), .A2(II22972) );
  NAND2_X1 NAND2_508( .ZN(II22974), .A1(g13962), .A2(II22972) );
  NAND2_X2 NAND2_509( .ZN(g17016), .A1(II22973), .A2(II22974) );
  NAND2_X2 NAND2_510( .ZN(II22981), .A1(g15274), .A2(g14106) );
  NAND2_X2 NAND2_511( .ZN(II22982), .A1(g15274), .A2(II22981) );
  NAND2_X1 NAND2_512( .ZN(II22983), .A1(g14106), .A2(II22981) );
  NAND2_X1 NAND2_513( .ZN(g17019), .A1(II22982), .A2(II22983) );
  NAND2_X1 NAND2_514( .ZN(II22988), .A1(g15296), .A2(g14321) );
  NAND2_X1 NAND2_515( .ZN(II22989), .A1(g15296), .A2(II22988) );
  NAND2_X1 NAND2_516( .ZN(II22990), .A1(g14321), .A2(II22988) );
  NAND2_X1 NAND2_517( .ZN(g17020), .A1(II22989), .A2(II22990) );
  NAND2_X1 NAND2_518( .ZN(II22998), .A1(g9187), .A2(g13872) );
  NAND2_X1 NAND2_519( .ZN(II22999), .A1(g9187), .A2(II22998) );
  NAND2_X1 NAND2_520( .ZN(II23000), .A1(g13872), .A2(II22998) );
  NAND2_X1 NAND2_521( .ZN(g17024), .A1(II22999), .A2(II23000) );
  NAND2_X1 NAND2_522( .ZN(II23008), .A1(g9203), .A2(g13926) );
  NAND2_X1 NAND2_523( .ZN(II23009), .A1(g9203), .A2(II23008) );
  NAND2_X1 NAND2_524( .ZN(II23010), .A1(g13926), .A2(II23008) );
  NAND2_X1 NAND2_525( .ZN(g17030), .A1(II23009), .A2(II23010) );
  NAND2_X1 NAND2_526( .ZN(II23018), .A1(g9216), .A2(g14032) );
  NAND2_X1 NAND2_527( .ZN(II23019), .A1(g9216), .A2(II23018) );
  NAND2_X1 NAND2_528( .ZN(II23020), .A1(g14032), .A2(II23018) );
  NAND2_X1 NAND2_529( .ZN(g17046), .A1(II23019), .A2(II23020) );
  NAND2_X1 NAND2_530( .ZN(II23027), .A1(g15366), .A2(g14221) );
  NAND2_X1 NAND2_531( .ZN(II23028), .A1(g15366), .A2(II23027) );
  NAND2_X1 NAND2_532( .ZN(II23029), .A1(g14221), .A2(II23027) );
  NAND2_X1 NAND2_533( .ZN(g17049), .A1(II23028), .A2(II23029) );
  NAND2_X1 NAND2_534( .ZN(II23034), .A1(g9232), .A2(g13864) );
  NAND2_X1 NAND2_535( .ZN(II23035), .A1(g9232), .A2(II23034) );
  NAND2_X1 NAND2_536( .ZN(II23036), .A1(g13864), .A2(II23034) );
  NAND2_X1 NAND2_537( .ZN(g17050), .A1(II23035), .A2(II23036) );
  NAND2_X1 NAND2_538( .ZN(II23045), .A1(g9248), .A2(g13894) );
  NAND2_X1 NAND2_539( .ZN(II23046), .A1(g9248), .A2(II23045) );
  NAND2_X1 NAND2_540( .ZN(II23047), .A1(g13894), .A2(II23045) );
  NAND2_X1 NAND2_541( .ZN(g17058), .A1(II23046), .A2(II23047) );
  NAND2_X1 NAND2_542( .ZN(II23055), .A1(g9264), .A2(g13982) );
  NAND2_X1 NAND2_543( .ZN(II23056), .A1(g9264), .A2(II23055) );
  NAND2_X1 NAND2_544( .ZN(II23057), .A1(g13982), .A2(II23055) );
  NAND2_X1 NAND2_545( .ZN(g17064), .A1(II23056), .A2(II23057) );
  NAND2_X1 NAND2_546( .ZN(II23065), .A1(g9277), .A2(g14123) );
  NAND2_X1 NAND2_547( .ZN(II23066), .A1(g9277), .A2(II23065) );
  NAND2_X1 NAND2_548( .ZN(II23067), .A1(g14123), .A2(II23065) );
  NAND2_X1 NAND2_549( .ZN(g17080), .A1(II23066), .A2(II23067) );
  NAND2_X1 NAND2_550( .ZN(II23074), .A1(g9293), .A2(g13856) );
  NAND2_X1 NAND2_551( .ZN(II23075), .A1(g9293), .A2(II23074) );
  NAND2_X1 NAND2_552( .ZN(II23076), .A1(g13856), .A2(II23074) );
  NAND2_X1 NAND2_553( .ZN(g17083), .A1(II23075), .A2(II23076) );
  NAND2_X1 NAND2_554( .ZN(II23082), .A1(g9310), .A2(g13879) );
  NAND2_X1 NAND2_555( .ZN(II23083), .A1(g9310), .A2(II23082) );
  NAND2_X1 NAND2_556( .ZN(II23084), .A1(g13879), .A2(II23082) );
  NAND2_X1 NAND2_557( .ZN(g17085), .A1(II23083), .A2(II23084) );
  NAND2_X1 NAND2_558( .ZN(II23093), .A1(g9326), .A2(g13935) );
  NAND2_X1 NAND2_559( .ZN(II23094), .A1(g9326), .A2(II23093) );
  NAND2_X1 NAND2_560( .ZN(II23095), .A1(g13935), .A2(II23093) );
  NAND2_X1 NAND2_561( .ZN(g17093), .A1(II23094), .A2(II23095) );
  NAND2_X1 NAND2_562( .ZN(II23103), .A1(g9342), .A2(g14052) );
  NAND2_X1 NAND2_563( .ZN(II23104), .A1(g9342), .A2(II23103) );
  NAND2_X1 NAND2_564( .ZN(II23105), .A1(g14052), .A2(II23103) );
  NAND2_X1 NAND2_565( .ZN(g17099), .A1(II23104), .A2(II23105) );
  NAND2_X1 NAND2_566( .ZN(II23113), .A1(g9356), .A2(g13848) );
  NAND2_X1 NAND2_567( .ZN(II23114), .A1(g9356), .A2(II23113) );
  NAND2_X1 NAND2_568( .ZN(II23115), .A1(g13848), .A2(II23113) );
  NAND2_X1 NAND2_569( .ZN(g17115), .A1(II23114), .A2(II23115) );
  NAND2_X1 NAND2_570( .ZN(g17118), .A1(g13915), .A2(g13893) );
  NAND2_X1 NAND2_571( .ZN(II23123), .A1(g9374), .A2(g13866) );
  NAND2_X1 NAND2_572( .ZN(II23124), .A1(g9374), .A2(II23123) );
  NAND2_X1 NAND2_573( .ZN(II23125), .A1(g13866), .A2(II23123) );
  NAND2_X1 NAND2_574( .ZN(g17121), .A1(II23124), .A2(II23125) );
  NAND2_X1 NAND2_575( .ZN(II23131), .A1(g9391), .A2(g13901) );
  NAND2_X1 NAND2_576( .ZN(II23132), .A1(g9391), .A2(II23131) );
  NAND2_X1 NAND2_577( .ZN(II23133), .A1(g13901), .A2(II23131) );
  NAND2_X1 NAND2_578( .ZN(g17123), .A1(II23132), .A2(II23133) );
  NAND2_X1 NAND2_579( .ZN(II23142), .A1(g9407), .A2(g13991) );
  NAND2_X1 NAND2_580( .ZN(II23143), .A1(g9407), .A2(II23142) );
  NAND2_X1 NAND2_581( .ZN(II23144), .A1(g13991), .A2(II23142) );
  NAND2_X1 NAND2_582( .ZN(g17131), .A1(II23143), .A2(II23144) );
  NAND2_X1 NAND2_583( .ZN(II23152), .A1(g9427), .A2(g14061) );
  NAND2_X1 NAND2_584( .ZN(II23153), .A1(g9427), .A2(II23152) );
  NAND2_X1 NAND2_585( .ZN(II23154), .A1(g14061), .A2(II23152) );
  NAND2_X1 NAND2_586( .ZN(g17137), .A1(II23153), .A2(II23154) );
  NAND2_X1 NAND2_587( .ZN(g17139), .A1(g13957), .A2(g13915) );
  NAND2_X1 NAND2_588( .ZN(II23161), .A1(g9453), .A2(g13857) );
  NAND2_X1 NAND2_589( .ZN(II23162), .A1(g9453), .A2(II23161) );
  NAND2_X1 NAND2_590( .ZN(II23163), .A1(g13857), .A2(II23161) );
  NAND2_X1 NAND2_591( .ZN(g17142), .A1(II23162), .A2(II23163) );
  NAND2_X1 NAND2_592( .ZN(g17145), .A1(g13971), .A2(g13934) );
  NAND2_X1 NAND2_593( .ZN(II23171), .A1(g9471), .A2(g13881) );
  NAND2_X1 NAND2_594( .ZN(II23172), .A1(g9471), .A2(II23171) );
  NAND2_X1 NAND2_595( .ZN(II23173), .A1(g13881), .A2(II23171) );
  NAND2_X1 NAND2_596( .ZN(g17148), .A1(II23172), .A2(II23173) );
  NAND2_X1 NAND2_597( .ZN(II23179), .A1(g9488), .A2(g13942) );
  NAND2_X1 NAND2_598( .ZN(II23180), .A1(g9488), .A2(II23179) );
  NAND2_X1 NAND2_599( .ZN(II23181), .A1(g13942), .A2(II23179) );
  NAND2_X1 NAND2_600( .ZN(g17150), .A1(II23180), .A2(II23181) );
  NAND2_X1 NAND2_601( .ZN(II23190), .A1(g9507), .A2(g13999) );
  NAND2_X1 NAND2_602( .ZN(II23191), .A1(g9507), .A2(II23190) );
  NAND2_X1 NAND2_603( .ZN(II23192), .A1(g13999), .A2(II23190) );
  NAND2_X1 NAND2_604( .ZN(g17158), .A1(II23191), .A2(II23192) );
  NAND2_X1 NAND2_605( .ZN(g17159), .A1(g14642), .A2(g14657) );
  NAND2_X1 NAND2_606( .ZN(II23198), .A1(g9569), .A2(g14176) );
  NAND2_X1 NAND2_607( .ZN(II23199), .A1(g9569), .A2(II23198) );
  NAND2_X1 NAND2_608( .ZN(II23200), .A1(g14176), .A2(II23198) );
  NAND2_X1 NAND2_609( .ZN(g17160), .A1(II23199), .A2(II23200) );
  NAND2_X1 NAND2_610( .ZN(g17162), .A1(g14027), .A2(g13971) );
  NAND2_X1 NAND2_611( .ZN(II23207), .A1(g9595), .A2(g13867) );
  NAND2_X1 NAND2_612( .ZN(II23208), .A1(g9595), .A2(II23207) );
  NAND2_X1 NAND2_613( .ZN(II23209), .A1(g13867), .A2(II23207) );
  NAND2_X1 NAND2_614( .ZN(g17165), .A1(II23208), .A2(II23209) );
  NAND2_X1 NAND2_615( .ZN(g17168), .A1(g14041), .A2(g13990) );
  NAND2_X1 NAND2_616( .ZN(II23217), .A1(g9613), .A2(g13903) );
  NAND2_X1 NAND2_617( .ZN(II23218), .A1(g9613), .A2(II23217) );
  NAND2_X1 NAND2_618( .ZN(II23219), .A1(g13903), .A2(II23217) );
  NAND2_X1 NAND2_619( .ZN(g17171), .A1(II23218), .A2(II23219) );
  NAND2_X1 NAND2_620( .ZN(II23225), .A1(g9649), .A2(g14090) );
  NAND2_X1 NAND2_621( .ZN(II23226), .A1(g9649), .A2(II23225) );
  NAND2_X1 NAND2_622( .ZN(II23227), .A1(g14090), .A2(II23225) );
  NAND2_X1 NAND2_623( .ZN(g17173), .A1(II23226), .A2(II23227) );
  NAND2_X1 NAND2_624( .ZN(g17174), .A1(g14669), .A2(g14691) );
  NAND2_X1 NAND2_625( .ZN(II23233), .A1(g9711), .A2(g14291) );
  NAND2_X1 NAND2_626( .ZN(II23234), .A1(g9711), .A2(II23233) );
  NAND2_X1 NAND2_627( .ZN(II23235), .A1(g14291), .A2(II23233) );
  NAND2_X1 NAND2_628( .ZN(g17175), .A1(II23234), .A2(II23235) );
  NAND2_X1 NAND2_629( .ZN(g17177), .A1(g14118), .A2(g14041) );
  NAND2_X1 NAND2_630( .ZN(II23242), .A1(g9737), .A2(g13882) );
  NAND2_X1 NAND2_631( .ZN(II23243), .A1(g9737), .A2(II23242) );
  NAND2_X1 NAND2_632( .ZN(II23244), .A1(g13882), .A2(II23242) );
  NAND2_X1 NAND2_633( .ZN(g17180), .A1(II23243), .A2(II23244) );
  NAND2_X1 NAND2_634( .ZN(g17183), .A1(g14132), .A2(g14060) );
  NAND2_X1 NAND2_635( .ZN(II23256), .A1(g9795), .A2(g14205) );
  NAND2_X1 NAND2_636( .ZN(II23257), .A1(g9795), .A2(II23256) );
  NAND2_X1 NAND2_637( .ZN(II23258), .A1(g14205), .A2(II23256) );
  NAND2_X1 NAND2_638( .ZN(g17190), .A1(II23257), .A2(II23258) );
  NAND2_X1 NAND2_639( .ZN(g17191), .A1(g14703), .A2(g14725) );
  NAND2_X1 NAND2_640( .ZN(II23264), .A1(g9857), .A2(g14413) );
  NAND2_X1 NAND2_641( .ZN(II23265), .A1(g9857), .A2(II23264) );
  NAND2_X1 NAND2_642( .ZN(II23266), .A1(g14413), .A2(II23264) );
  NAND2_X1 NAND2_643( .ZN(g17192), .A1(II23265), .A2(II23266) );
  NAND2_X1 NAND2_644( .ZN(g17194), .A1(g14233), .A2(g14132) );
  NAND2_X1 NAND2_645( .ZN(II23277), .A1(g9941), .A2(g14320) );
  NAND2_X1 NAND2_646( .ZN(II23278), .A1(g9941), .A2(II23277) );
  NAND2_X1 NAND2_647( .ZN(II23279), .A1(g14320), .A2(II23277) );
  NAND2_X1 NAND2_648( .ZN(g17201), .A1(II23278), .A2(II23279) );
  NAND2_X1 NAND2_649( .ZN(g17202), .A1(g14737), .A2(g14753) );
  NAND2_X1 NAND2_650( .ZN(II23806), .A1(g14062), .A2(g9150) );
  NAND2_X1 NAND2_651( .ZN(II23807), .A1(g14062), .A2(II23806) );
  NAND2_X1 NAND2_652( .ZN(II23808), .A1(g9150), .A2(II23806) );
  NAND2_X1 NAND2_653( .ZN(g17729), .A1(II23807), .A2(II23808) );
  NAND2_X1 NAND2_654( .ZN(II23878), .A1(g14001), .A2(g9187) );
  NAND2_X1 NAND2_655( .ZN(II23879), .A1(g14001), .A2(II23878) );
  NAND2_X1 NAND2_656( .ZN(II23880), .A1(g9187), .A2(II23878) );
  NAND2_X1 NAND2_657( .ZN(g17807), .A1(II23879), .A2(II23880) );
  NAND2_X1 NAND2_658( .ZN(II23893), .A1(g14177), .A2(g9174) );
  NAND2_X1 NAND2_659( .ZN(II23894), .A1(g14177), .A2(II23893) );
  NAND2_X1 NAND2_660( .ZN(II23895), .A1(g9174), .A2(II23893) );
  NAND2_X1 NAND2_661( .ZN(g17830), .A1(II23894), .A2(II23895) );
  NAND2_X1 NAND2_662( .ZN(II23941), .A1(g13946), .A2(g9293) );
  NAND2_X1 NAND2_663( .ZN(II23942), .A1(g13946), .A2(II23941) );
  NAND2_X1 NAND2_664( .ZN(II23943), .A1(g9293), .A2(II23941) );
  NAND2_X1 NAND2_665( .ZN(g17887), .A1(II23942), .A2(II23943) );
  NAND2_X1 NAND2_666( .ZN(II23958), .A1(g6513), .A2(g14171) );
  NAND2_X1 NAND2_667( .ZN(II23959), .A1(g6513), .A2(II23958) );
  NAND2_X1 NAND2_668( .ZN(II23960), .A1(g14171), .A2(II23958) );
  NAND2_X1 NAND2_669( .ZN(g17913), .A1(II23959), .A2(II23960) );
  NAND2_X1 NAND2_670( .ZN(II23966), .A1(g14092), .A2(g9248) );
  NAND2_X1 NAND2_671( .ZN(II23967), .A1(g14092), .A2(II23966) );
  NAND2_X1 NAND2_672( .ZN(II23968), .A1(g9248), .A2(II23966) );
  NAND2_X1 NAND2_673( .ZN(g17919), .A1(II23967), .A2(II23968) );
  NAND2_X1 NAND2_674( .ZN(II23981), .A1(g14292), .A2(g9216) );
  NAND2_X1 NAND2_675( .ZN(II23982), .A1(g14292), .A2(II23981) );
  NAND2_X1 NAND2_676( .ZN(II23983), .A1(g9216), .A2(II23981) );
  NAND2_X1 NAND2_677( .ZN(g17942), .A1(II23982), .A2(II23983) );
  NAND2_X1 NAND2_678( .ZN(II24005), .A1(g7548), .A2(g15814) );
  NAND2_X1 NAND2_679( .ZN(II24006), .A1(g7548), .A2(II24005) );
  NAND2_X1 NAND2_680( .ZN(II24007), .A1(g15814), .A2(II24005) );
  NAND2_X1 NAND2_681( .ZN(g17968), .A1(II24006), .A2(II24007) );
  NAND2_X2 NAND2_682( .ZN(II24015), .A1(g13907), .A2(g9427) );
  NAND2_X2 NAND2_683( .ZN(II24016), .A1(g13907), .A2(II24015) );
  NAND2_X1 NAND2_684( .ZN(II24017), .A1(g9427), .A2(II24015) );
  NAND2_X1 NAND2_685( .ZN(g17979), .A1(II24016), .A2(II24017) );
  NAND2_X1 NAND2_686( .ZN(g17985), .A1(g14641), .A2(g9636) );
  NAND2_X1 NAND2_687( .ZN(II24028), .A1(g6201), .A2(g14086) );
  NAND2_X1 NAND2_688( .ZN(II24029), .A1(g6201), .A2(II24028) );
  NAND2_X1 NAND2_689( .ZN(II24030), .A1(g14086), .A2(II24028) );
  NAND2_X1 NAND2_690( .ZN(g17992), .A1(II24029), .A2(II24030) );
  NAND2_X1 NAND2_691( .ZN(II24036), .A1(g14016), .A2(g9374) );
  NAND2_X1 NAND2_692( .ZN(II24037), .A1(g14016), .A2(II24036) );
  NAND2_X1 NAND2_693( .ZN(II24038), .A1(g9374), .A2(II24036) );
  NAND2_X1 NAND2_694( .ZN(g17998), .A1(II24037), .A2(II24038) );
  NAND2_X1 NAND2_695( .ZN(II24053), .A1(g6777), .A2(g14286) );
  NAND2_X1 NAND2_696( .ZN(II24054), .A1(g6777), .A2(II24053) );
  NAND2_X1 NAND2_697( .ZN(II24055), .A1(g14286), .A2(II24053) );
  NAND2_X1 NAND2_698( .ZN(g18024), .A1(II24054), .A2(II24055) );
  NAND2_X1 NAND2_699( .ZN(II24061), .A1(g14207), .A2(g9326) );
  NAND2_X1 NAND2_700( .ZN(II24062), .A1(g14207), .A2(II24061) );
  NAND2_X1 NAND2_701( .ZN(II24063), .A1(g9326), .A2(II24061) );
  NAND2_X1 NAND2_702( .ZN(g18030), .A1(II24062), .A2(II24063) );
  NAND2_X1 NAND2_703( .ZN(II24076), .A1(g14414), .A2(g9277) );
  NAND2_X1 NAND2_704( .ZN(II24077), .A1(g14414), .A2(II24076) );
  NAND2_X1 NAND2_705( .ZN(II24078), .A1(g9277), .A2(II24076) );
  NAND2_X1 NAND2_706( .ZN(g18053), .A1(II24077), .A2(II24078) );
  NAND2_X1 NAND2_707( .ZN(II24091), .A1(g13886), .A2(g15096) );
  NAND2_X1 NAND2_708( .ZN(II24092), .A1(g13886), .A2(II24091) );
  NAND2_X1 NAND2_709( .ZN(II24093), .A1(g15096), .A2(II24091) );
  NAND2_X1 NAND2_710( .ZN(g18079), .A1(II24092), .A2(II24093) );
  NAND2_X1 NAND2_711( .ZN(II24102), .A1(g6363), .A2(g14011) );
  NAND2_X1 NAND2_712( .ZN(II24103), .A1(g6363), .A2(II24102) );
  NAND2_X1 NAND2_713( .ZN(II24104), .A1(g14011), .A2(II24102) );
  NAND2_X1 NAND2_714( .ZN(g18090), .A1(II24103), .A2(II24104) );
  NAND2_X1 NAND2_715( .ZN(II24110), .A1(g13963), .A2(g9569) );
  NAND2_X1 NAND2_716( .ZN(II24111), .A1(g13963), .A2(II24110) );
  NAND2_X1 NAND2_717( .ZN(II24112), .A1(g9569), .A2(II24110) );
  NAND2_X1 NAND2_718( .ZN(g18096), .A1(II24111), .A2(II24112) );
  NAND2_X1 NAND2_719( .ZN(g18102), .A1(g14668), .A2(g9782) );
  NAND2_X1 NAND2_720( .ZN(II24123), .A1(g6290), .A2(g14201) );
  NAND2_X1 NAND2_721( .ZN(II24124), .A1(g6290), .A2(II24123) );
  NAND2_X1 NAND2_722( .ZN(II24125), .A1(g14201), .A2(II24123) );
  NAND2_X1 NAND2_723( .ZN(g18109), .A1(II24124), .A2(II24125) );
  NAND2_X1 NAND2_724( .ZN(II24131), .A1(g14107), .A2(g9471) );
  NAND2_X1 NAND2_725( .ZN(II24132), .A1(g14107), .A2(II24131) );
  NAND2_X1 NAND2_726( .ZN(II24133), .A1(g9471), .A2(II24131) );
  NAND2_X1 NAND2_727( .ZN(g18115), .A1(II24132), .A2(II24133) );
  NAND2_X1 NAND2_728( .ZN(II24148), .A1(g7079), .A2(g14408) );
  NAND2_X1 NAND2_729( .ZN(II24149), .A1(g7079), .A2(II24148) );
  NAND2_X1 NAND2_730( .ZN(II24150), .A1(g14408), .A2(II24148) );
  NAND2_X1 NAND2_731( .ZN(g18141), .A1(II24149), .A2(II24150) );
  NAND2_X1 NAND2_732( .ZN(II24156), .A1(g14322), .A2(g9407) );
  NAND2_X1 NAND2_733( .ZN(II24157), .A1(g14322), .A2(II24156) );
  NAND2_X1 NAND2_734( .ZN(II24158), .A1(g9407), .A2(II24156) );
  NAND2_X1 NAND2_735( .ZN(g18147), .A1(II24157), .A2(II24158) );
  NAND2_X1 NAND2_736( .ZN(II24178), .A1(g13873), .A2(g9161) );
  NAND2_X1 NAND2_737( .ZN(II24179), .A1(g13873), .A2(II24178) );
  NAND2_X1 NAND2_738( .ZN(II24180), .A1(g9161), .A2(II24178) );
  NAND2_X1 NAND2_739( .ZN(g18183), .A1(II24179), .A2(II24180) );
  NAND2_X1 NAND2_740( .ZN(II24186), .A1(g6177), .A2(g13958) );
  NAND2_X1 NAND2_741( .ZN(II24187), .A1(g6177), .A2(II24186) );
  NAND2_X1 NAND2_742( .ZN(II24188), .A1(g13958), .A2(II24186) );
  NAND2_X1 NAND2_743( .ZN(g18189), .A1(II24187), .A2(II24188) );
  NAND2_X1 NAND2_744( .ZN(II24194), .A1(g13927), .A2(g15188) );
  NAND2_X1 NAND2_745( .ZN(II24195), .A1(g13927), .A2(II24194) );
  NAND2_X1 NAND2_746( .ZN(II24196), .A1(g15188), .A2(II24194) );
  NAND2_X1 NAND2_747( .ZN(g18195), .A1(II24195), .A2(II24196) );
  NAND2_X1 NAND2_748( .ZN(II24205), .A1(g6568), .A2(g14102) );
  NAND2_X1 NAND2_749( .ZN(II24206), .A1(g6568), .A2(II24205) );
  NAND2_X1 NAND2_750( .ZN(II24207), .A1(g14102), .A2(II24205) );
  NAND2_X1 NAND2_751( .ZN(g18206), .A1(II24206), .A2(II24207) );
  NAND2_X1 NAND2_752( .ZN(II24213), .A1(g14033), .A2(g9711) );
  NAND2_X1 NAND2_753( .ZN(II24214), .A1(g14033), .A2(II24213) );
  NAND2_X1 NAND2_754( .ZN(II24215), .A1(g9711), .A2(II24213) );
  NAND2_X1 NAND2_755( .ZN(g18212), .A1(II24214), .A2(II24215) );
  NAND2_X1 NAND2_756( .ZN(g18218), .A1(g14702), .A2(g9928) );
  NAND2_X1 NAND2_757( .ZN(II24226), .A1(g6427), .A2(g14316) );
  NAND2_X1 NAND2_758( .ZN(II24227), .A1(g6427), .A2(II24226) );
  NAND2_X1 NAND2_759( .ZN(II24228), .A1(g14316), .A2(II24226) );
  NAND2_X1 NAND2_760( .ZN(g18225), .A1(II24227), .A2(II24228) );
  NAND2_X1 NAND2_761( .ZN(II24234), .A1(g14222), .A2(g9613) );
  NAND2_X1 NAND2_762( .ZN(II24235), .A1(g14222), .A2(II24234) );
  NAND2_X1 NAND2_763( .ZN(II24236), .A1(g9613), .A2(II24234) );
  NAND2_X1 NAND2_764( .ZN(g18231), .A1(II24235), .A2(II24236) );
  NAND2_X1 NAND2_765( .ZN(II24251), .A1(g7329), .A2(g14520) );
  NAND2_X1 NAND2_766( .ZN(II24252), .A1(g7329), .A2(II24251) );
  NAND2_X1 NAND2_767( .ZN(II24253), .A1(g14520), .A2(II24251) );
  NAND2_X1 NAND2_768( .ZN(g18257), .A1(II24252), .A2(II24253) );
  NAND2_X1 NAND2_769( .ZN(II24263), .A1(g14342), .A2(g9232) );
  NAND2_X1 NAND2_770( .ZN(II24264), .A1(g14342), .A2(II24263) );
  NAND2_X1 NAND2_771( .ZN(II24265), .A1(g9232), .A2(II24263) );
  NAND2_X1 NAND2_772( .ZN(g18270), .A1(II24264), .A2(II24265) );
  NAND2_X1 NAND2_773( .ZN(II24271), .A1(g6180), .A2(g13922) );
  NAND2_X1 NAND2_774( .ZN(II24272), .A1(g6180), .A2(II24271) );
  NAND2_X1 NAND2_775( .ZN(II24273), .A1(g13922), .A2(II24271) );
  NAND2_X1 NAND2_776( .ZN(g18276), .A1(II24272), .A2(II24273) );
  NAND2_X1 NAND2_777( .ZN(II24278), .A1(g6284), .A2(g13918) );
  NAND2_X1 NAND2_778( .ZN(II24279), .A1(g6284), .A2(II24278) );
  NAND2_X1 NAND2_779( .ZN(II24280), .A1(g13918), .A2(II24278) );
  NAND2_X1 NAND2_780( .ZN(g18277), .A1(II24279), .A2(II24280) );
  NAND2_X1 NAND2_781( .ZN(II24290), .A1(g13895), .A2(g9203) );
  NAND2_X1 NAND2_782( .ZN(II24291), .A1(g13895), .A2(II24290) );
  NAND2_X1 NAND2_783( .ZN(II24292), .A1(g9203), .A2(II24290) );
  NAND2_X1 NAND2_784( .ZN(g18290), .A1(II24291), .A2(II24292) );
  NAND2_X1 NAND2_785( .ZN(II24298), .A1(g6209), .A2(g14028) );
  NAND2_X1 NAND2_786( .ZN(II24299), .A1(g6209), .A2(II24298) );
  NAND2_X1 NAND2_787( .ZN(II24300), .A1(g14028), .A2(II24298) );
  NAND2_X1 NAND2_788( .ZN(g18296), .A1(II24299), .A2(II24300) );
  NAND2_X1 NAND2_789( .ZN(II24306), .A1(g13983), .A2(g15274) );
  NAND2_X1 NAND2_790( .ZN(II24307), .A1(g13983), .A2(II24306) );
  NAND2_X1 NAND2_791( .ZN(II24308), .A1(g15274), .A2(II24306) );
  NAND2_X1 NAND2_792( .ZN(g18302), .A1(II24307), .A2(II24308) );
  NAND2_X1 NAND2_793( .ZN(II24317), .A1(g6832), .A2(g14217) );
  NAND2_X1 NAND2_794( .ZN(II24318), .A1(g6832), .A2(II24317) );
  NAND2_X2 NAND2_795( .ZN(II24319), .A1(g14217), .A2(II24317) );
  NAND2_X2 NAND2_796( .ZN(g18313), .A1(II24318), .A2(II24319) );
  NAND2_X2 NAND2_797( .ZN(II24325), .A1(g14124), .A2(g9857) );
  NAND2_X2 NAND2_798( .ZN(II24326), .A1(g14124), .A2(II24325) );
  NAND2_X1 NAND2_799( .ZN(II24327), .A1(g9857), .A2(II24325) );
  NAND2_X1 NAND2_800( .ZN(g18319), .A1(II24326), .A2(II24327) );
  NAND2_X1 NAND2_801( .ZN(g18325), .A1(g14736), .A2(g10082) );
  NAND2_X1 NAND2_802( .ZN(II24338), .A1(g6632), .A2(g14438) );
  NAND2_X1 NAND2_803( .ZN(II24339), .A1(g6632), .A2(II24338) );
  NAND2_X1 NAND2_804( .ZN(II24340), .A1(g14438), .A2(II24338) );
  NAND2_X1 NAND2_805( .ZN(g18332), .A1(II24339), .A2(II24340) );
  NAND2_X1 NAND2_806( .ZN(II24351), .A1(g14238), .A2(g9356) );
  NAND2_X1 NAND2_807( .ZN(II24352), .A1(g14238), .A2(II24351) );
  NAND2_X1 NAND2_808( .ZN(II24353), .A1(g9356), .A2(II24351) );
  NAND2_X1 NAND2_809( .ZN(g18346), .A1(II24352), .A2(II24353) );
  NAND2_X1 NAND2_810( .ZN(II24361), .A1(g6157), .A2(g14525) );
  NAND2_X1 NAND2_811( .ZN(II24362), .A1(g6157), .A2(II24361) );
  NAND2_X1 NAND2_812( .ZN(II24363), .A1(g14525), .A2(II24361) );
  NAND2_X1 NAND2_813( .ZN(g18354), .A1(II24362), .A2(II24363) );
  NAND2_X1 NAND2_814( .ZN(II24372), .A1(g14454), .A2(g9310) );
  NAND2_X1 NAND2_815( .ZN(II24373), .A1(g14454), .A2(II24372) );
  NAND2_X1 NAND2_816( .ZN(II24374), .A1(g9310), .A2(II24372) );
  NAND2_X1 NAND2_817( .ZN(g18363), .A1(II24373), .A2(II24374) );
  NAND2_X1 NAND2_818( .ZN(II24380), .A1(g6212), .A2(g13978) );
  NAND2_X1 NAND2_819( .ZN(II24381), .A1(g6212), .A2(II24380) );
  NAND2_X1 NAND2_820( .ZN(II24382), .A1(g13978), .A2(II24380) );
  NAND2_X1 NAND2_821( .ZN(g18369), .A1(II24381), .A2(II24382) );
  NAND2_X1 NAND2_822( .ZN(II24387), .A1(g6421), .A2(g13974) );
  NAND2_X1 NAND2_823( .ZN(II24388), .A1(g6421), .A2(II24387) );
  NAND2_X1 NAND2_824( .ZN(II24389), .A1(g13974), .A2(II24387) );
  NAND2_X1 NAND2_825( .ZN(g18370), .A1(II24388), .A2(II24389) );
  NAND2_X1 NAND2_826( .ZN(II24399), .A1(g13936), .A2(g9264) );
  NAND2_X1 NAND2_827( .ZN(II24400), .A1(g13936), .A2(II24399) );
  NAND2_X1 NAND2_828( .ZN(II24401), .A1(g9264), .A2(II24399) );
  NAND2_X1 NAND2_829( .ZN(g18383), .A1(II24400), .A2(II24401) );
  NAND2_X1 NAND2_830( .ZN(II24407), .A1(g6298), .A2(g14119) );
  NAND2_X1 NAND2_831( .ZN(II24408), .A1(g6298), .A2(II24407) );
  NAND2_X1 NAND2_832( .ZN(II24409), .A1(g14119), .A2(II24407) );
  NAND2_X1 NAND2_833( .ZN(g18389), .A1(II24408), .A2(II24409) );
  NAND2_X1 NAND2_834( .ZN(II24415), .A1(g14053), .A2(g15366) );
  NAND2_X1 NAND2_835( .ZN(II24416), .A1(g14053), .A2(II24415) );
  NAND2_X1 NAND2_836( .ZN(II24417), .A1(g15366), .A2(II24415) );
  NAND2_X1 NAND2_837( .ZN(g18395), .A1(II24416), .A2(II24417) );
  NAND2_X1 NAND2_838( .ZN(II24426), .A1(g7134), .A2(g14332) );
  NAND2_X1 NAND2_839( .ZN(II24427), .A1(g7134), .A2(II24426) );
  NAND2_X1 NAND2_840( .ZN(II24428), .A1(g14332), .A2(II24426) );
  NAND2_X1 NAND2_841( .ZN(g18406), .A1(II24427), .A2(II24428) );
  NAND2_X1 NAND2_842( .ZN(II24436), .A1(g14153), .A2(g15022) );
  NAND2_X1 NAND2_843( .ZN(II24437), .A1(g14153), .A2(II24436) );
  NAND2_X1 NAND2_844( .ZN(II24438), .A1(g15022), .A2(II24436) );
  NAND2_X1 NAND2_845( .ZN(g18419), .A1(II24437), .A2(II24438) );
  NAND2_X1 NAND2_846( .ZN(II24443), .A1(g14148), .A2(g9507) );
  NAND2_X1 NAND2_847( .ZN(II24444), .A1(g14148), .A2(II24443) );
  NAND2_X1 NAND2_848( .ZN(II24445), .A1(g9507), .A2(II24443) );
  NAND2_X1 NAND2_849( .ZN(g18424), .A1(II24444), .A2(II24445) );
  NAND2_X1 NAND2_850( .ZN(II24452), .A1(g6142), .A2(g14450) );
  NAND2_X1 NAND2_851( .ZN(II24453), .A1(g6142), .A2(II24452) );
  NAND2_X1 NAND2_852( .ZN(II24454), .A1(g14450), .A2(II24452) );
  NAND2_X1 NAND2_853( .ZN(g18431), .A1(II24453), .A2(II24454) );
  NAND2_X1 NAND2_854( .ZN(II24464), .A1(g14360), .A2(g9453) );
  NAND2_X1 NAND2_855( .ZN(II24465), .A1(g14360), .A2(II24464) );
  NAND2_X1 NAND2_856( .ZN(II24466), .A1(g9453), .A2(II24464) );
  NAND2_X1 NAND2_857( .ZN(g18441), .A1(II24465), .A2(II24466) );
  NAND2_X1 NAND2_858( .ZN(II24474), .A1(g6184), .A2(g14580) );
  NAND2_X1 NAND2_859( .ZN(II24475), .A1(g6184), .A2(II24474) );
  NAND2_X1 NAND2_860( .ZN(II24476), .A1(g14580), .A2(II24474) );
  NAND2_X1 NAND2_861( .ZN(g18449), .A1(II24475), .A2(II24476) );
  NAND2_X1 NAND2_862( .ZN(II24485), .A1(g14541), .A2(g9391) );
  NAND2_X1 NAND2_863( .ZN(II24486), .A1(g14541), .A2(II24485) );
  NAND2_X1 NAND2_864( .ZN(II24487), .A1(g9391), .A2(II24485) );
  NAND2_X1 NAND2_865( .ZN(g18458), .A1(II24486), .A2(II24487) );
  NAND2_X1 NAND2_866( .ZN(II24493), .A1(g6301), .A2(g14048) );
  NAND2_X1 NAND2_867( .ZN(II24494), .A1(g6301), .A2(II24493) );
  NAND2_X1 NAND2_868( .ZN(II24495), .A1(g14048), .A2(II24493) );
  NAND2_X1 NAND2_869( .ZN(g18464), .A1(II24494), .A2(II24495) );
  NAND2_X1 NAND2_870( .ZN(II24500), .A1(g6626), .A2(g14044) );
  NAND2_X1 NAND2_871( .ZN(II24501), .A1(g6626), .A2(II24500) );
  NAND2_X1 NAND2_872( .ZN(II24502), .A1(g14044), .A2(II24500) );
  NAND2_X1 NAND2_873( .ZN(g18465), .A1(II24501), .A2(II24502) );
  NAND2_X1 NAND2_874( .ZN(II24512), .A1(g13992), .A2(g9342) );
  NAND2_X1 NAND2_875( .ZN(II24513), .A1(g13992), .A2(II24512) );
  NAND2_X1 NAND2_876( .ZN(II24514), .A1(g9342), .A2(II24512) );
  NAND2_X1 NAND2_877( .ZN(g18478), .A1(II24513), .A2(II24514) );
  NAND2_X1 NAND2_878( .ZN(II24520), .A1(g6435), .A2(g14234) );
  NAND2_X1 NAND2_879( .ZN(II24521), .A1(g6435), .A2(II24520) );
  NAND2_X1 NAND2_880( .ZN(II24522), .A1(g14234), .A2(II24520) );
  NAND2_X1 NAND2_881( .ZN(g18484), .A1(II24521), .A2(II24522) );
  NAND2_X1 NAND2_882( .ZN(II24530), .A1(g6707), .A2(g14355) );
  NAND2_X1 NAND2_883( .ZN(II24531), .A1(g6707), .A2(II24530) );
  NAND2_X1 NAND2_884( .ZN(II24532), .A1(g14355), .A2(II24530) );
  NAND2_X1 NAND2_885( .ZN(g18491), .A1(II24531), .A2(II24532) );
  NAND2_X1 NAND2_886( .ZN(II24537), .A1(g14268), .A2(g15118) );
  NAND2_X1 NAND2_887( .ZN(II24538), .A1(g14268), .A2(II24537) );
  NAND2_X1 NAND2_888( .ZN(II24539), .A1(g15118), .A2(II24537) );
  NAND2_X1 NAND2_889( .ZN(g18492), .A1(II24538), .A2(II24539) );
  NAND2_X1 NAND2_890( .ZN(II24544), .A1(g14263), .A2(g9649) );
  NAND2_X1 NAND2_891( .ZN(II24545), .A1(g14263), .A2(II24544) );
  NAND2_X1 NAND2_892( .ZN(II24546), .A1(g9649), .A2(II24544) );
  NAND2_X1 NAND2_893( .ZN(g18497), .A1(II24545), .A2(II24546) );
  NAND2_X1 NAND2_894( .ZN(II24553), .A1(g6163), .A2(g14537) );
  NAND2_X1 NAND2_895( .ZN(II24554), .A1(g6163), .A2(II24553) );
  NAND2_X1 NAND2_896( .ZN(II24555), .A1(g14537), .A2(II24553) );
  NAND2_X1 NAND2_897( .ZN(g18504), .A1(II24554), .A2(II24555) );
  NAND2_X1 NAND2_898( .ZN(II24565), .A1(g14472), .A2(g9595) );
  NAND2_X1 NAND2_899( .ZN(II24566), .A1(g14472), .A2(II24565) );
  NAND2_X1 NAND2_900( .ZN(II24567), .A1(g9595), .A2(II24565) );
  NAND2_X1 NAND2_901( .ZN(g18514), .A1(II24566), .A2(II24567) );
  NAND2_X1 NAND2_902( .ZN(II24575), .A1(g6216), .A2(g14614) );
  NAND2_X1 NAND2_903( .ZN(II24576), .A1(g6216), .A2(II24575) );
  NAND2_X1 NAND2_904( .ZN(II24577), .A1(g14614), .A2(II24575) );
  NAND2_X1 NAND2_905( .ZN(g18522), .A1(II24576), .A2(II24577) );
  NAND2_X1 NAND2_906( .ZN(II24586), .A1(g14596), .A2(g9488) );
  NAND2_X1 NAND2_907( .ZN(II24587), .A1(g14596), .A2(II24586) );
  NAND2_X1 NAND2_908( .ZN(II24588), .A1(g9488), .A2(II24586) );
  NAND2_X1 NAND2_909( .ZN(g18531), .A1(II24587), .A2(II24588) );
  NAND2_X1 NAND2_910( .ZN(II24594), .A1(g6438), .A2(g14139) );
  NAND2_X1 NAND2_911( .ZN(II24595), .A1(g6438), .A2(II24594) );
  NAND2_X1 NAND2_912( .ZN(II24596), .A1(g14139), .A2(II24594) );
  NAND2_X1 NAND2_913( .ZN(g18537), .A1(II24595), .A2(II24596) );
  NAND2_X1 NAND2_914( .ZN(II24601), .A1(g6890), .A2(g14135) );
  NAND2_X1 NAND2_915( .ZN(II24602), .A1(g6890), .A2(II24601) );
  NAND2_X1 NAND2_916( .ZN(II24603), .A1(g14135), .A2(II24601) );
  NAND2_X1 NAND2_917( .ZN(g18538), .A1(II24602), .A2(II24603) );
  NAND2_X1 NAND2_918( .ZN(II24611), .A1(g15814), .A2(g15978) );
  NAND2_X1 NAND2_919( .ZN(II24612), .A1(g15814), .A2(II24611) );
  NAND2_X1 NAND2_920( .ZN(II24613), .A1(g15978), .A2(II24611) );
  NAND2_X1 NAND2_921( .ZN(g18542), .A1(II24612), .A2(II24613) );
  NAND2_X1 NAND2_922( .ZN(II24624), .A1(g6136), .A2(g14252) );
  NAND2_X2 NAND2_923( .ZN(II24625), .A1(g6136), .A2(II24624) );
  NAND2_X2 NAND2_924( .ZN(II24626), .A1(g14252), .A2(II24624) );
  NAND2_X1 NAND2_925( .ZN(g18553), .A1(II24625), .A2(II24626) );
  NAND2_X1 NAND2_926( .ZN(II24632), .A1(g7009), .A2(g14467) );
  NAND2_X1 NAND2_927( .ZN(II24633), .A1(g7009), .A2(II24632) );
  NAND2_X1 NAND2_928( .ZN(II24634), .A1(g14467), .A2(II24632) );
  NAND2_X1 NAND2_929( .ZN(g18555), .A1(II24633), .A2(II24634) );
  NAND2_X1 NAND2_930( .ZN(II24639), .A1(g14390), .A2(g15210) );
  NAND2_X1 NAND2_931( .ZN(II24640), .A1(g14390), .A2(II24639) );
  NAND2_X1 NAND2_932( .ZN(II24641), .A1(g15210), .A2(II24639) );
  NAND2_X1 NAND2_933( .ZN(g18556), .A1(II24640), .A2(II24641) );
  NAND2_X1 NAND2_934( .ZN(II24646), .A1(g14385), .A2(g9795) );
  NAND2_X1 NAND2_935( .ZN(II24647), .A1(g14385), .A2(II24646) );
  NAND2_X1 NAND2_936( .ZN(II24648), .A1(g9795), .A2(II24646) );
  NAND2_X1 NAND2_937( .ZN(g18561), .A1(II24647), .A2(II24648) );
  NAND2_X1 NAND2_938( .ZN(II24655), .A1(g6190), .A2(g14592) );
  NAND2_X1 NAND2_939( .ZN(II24656), .A1(g6190), .A2(II24655) );
  NAND2_X1 NAND2_940( .ZN(II24657), .A1(g14592), .A2(II24655) );
  NAND2_X1 NAND2_941( .ZN(g18568), .A1(II24656), .A2(II24657) );
  NAND2_X1 NAND2_942( .ZN(II24667), .A1(g14559), .A2(g9737) );
  NAND2_X1 NAND2_943( .ZN(II24668), .A1(g14559), .A2(II24667) );
  NAND2_X1 NAND2_944( .ZN(II24669), .A1(g9737), .A2(II24667) );
  NAND2_X1 NAND2_945( .ZN(g18578), .A1(II24668), .A2(II24669) );
  NAND2_X1 NAND2_946( .ZN(II24677), .A1(g6305), .A2(g14637) );
  NAND2_X1 NAND2_947( .ZN(II24678), .A1(g6305), .A2(II24677) );
  NAND2_X1 NAND2_948( .ZN(II24679), .A1(g14637), .A2(II24677) );
  NAND2_X1 NAND2_949( .ZN(g18586), .A1(II24678), .A2(II24679) );
  NAND2_X1 NAND2_950( .ZN(II24694), .A1(g6146), .A2(g14374) );
  NAND2_X1 NAND2_951( .ZN(II24695), .A1(g6146), .A2(II24694) );
  NAND2_X1 NAND2_952( .ZN(II24696), .A1(g14374), .A2(II24694) );
  NAND2_X1 NAND2_953( .ZN(g18603), .A1(II24695), .A2(II24696) );
  NAND2_X1 NAND2_954( .ZN(II24702), .A1(g7259), .A2(g14554) );
  NAND2_X1 NAND2_955( .ZN(II24703), .A1(g7259), .A2(II24702) );
  NAND2_X1 NAND2_956( .ZN(II24704), .A1(g14554), .A2(II24702) );
  NAND2_X1 NAND2_957( .ZN(g18605), .A1(II24703), .A2(II24704) );
  NAND2_X1 NAND2_958( .ZN(II24709), .A1(g14502), .A2(g15296) );
  NAND2_X1 NAND2_959( .ZN(II24710), .A1(g14502), .A2(II24709) );
  NAND2_X1 NAND2_960( .ZN(II24711), .A1(g15296), .A2(II24709) );
  NAND2_X1 NAND2_961( .ZN(g18606), .A1(II24710), .A2(II24711) );
  NAND2_X1 NAND2_962( .ZN(II24716), .A1(g14497), .A2(g9941) );
  NAND2_X1 NAND2_963( .ZN(II24717), .A1(g14497), .A2(II24716) );
  NAND2_X1 NAND2_964( .ZN(II24718), .A1(g9941), .A2(II24716) );
  NAND2_X1 NAND2_965( .ZN(g18611), .A1(II24717), .A2(II24718) );
  NAND2_X1 NAND2_966( .ZN(II24725), .A1(g6222), .A2(g14626) );
  NAND2_X1 NAND2_967( .ZN(II24726), .A1(g6222), .A2(II24725) );
  NAND2_X1 NAND2_968( .ZN(II24727), .A1(g14626), .A2(II24725) );
  NAND2_X1 NAND2_969( .ZN(g18618), .A1(II24726), .A2(II24727) );
  NAND2_X1 NAND2_970( .ZN(II24743), .A1(g6167), .A2(g14486) );
  NAND2_X1 NAND2_971( .ZN(II24744), .A1(g6167), .A2(II24743) );
  NAND2_X1 NAND2_972( .ZN(II24745), .A1(g14486), .A2(II24743) );
  NAND2_X1 NAND2_973( .ZN(g18635), .A1(II24744), .A2(II24745) );
  NAND2_X1 NAND2_974( .ZN(II24751), .A1(g7455), .A2(g14609) );
  NAND2_X2 NAND2_975( .ZN(II24752), .A1(g7455), .A2(II24751) );
  NAND2_X1 NAND2_976( .ZN(II24753), .A1(g14609), .A2(II24751) );
  NAND2_X1 NAND2_977( .ZN(g18637), .A1(II24752), .A2(II24753) );
  NAND2_X1 NAND2_978( .ZN(II24763), .A1(g6194), .A2(g14573) );
  NAND2_X1 NAND2_979( .ZN(II24764), .A1(g6194), .A2(II24763) );
  NAND2_X1 NAND2_980( .ZN(II24765), .A1(g14573), .A2(II24763) );
  NAND2_X1 NAND2_981( .ZN(g18644), .A1(II24764), .A2(II24765) );
  NAND2_X1 NAND2_982( .ZN(g18977), .A1(g15797), .A2(g3006) );
  NAND2_X1 NAND2_983( .ZN(II25030), .A1(g8029), .A2(g13507) );
  NAND2_X1 NAND2_984( .ZN(II25031), .A1(g8029), .A2(II25030) );
  NAND2_X1 NAND2_985( .ZN(II25032), .A1(g13507), .A2(II25030) );
  NAND2_X1 NAND2_986( .ZN(g18980), .A1(II25031), .A2(II25032) );
  NAND2_X1 NAND2_987( .ZN(g19067), .A1(g16554), .A2(g16578) );
  NAND2_X1 NAND2_988( .ZN(g19084), .A1(g16586), .A2(g16602) );
  NAND2_X1 NAND2_989( .ZN(g19103), .A1(g18590), .A2(g2924) );
  NAND2_X1 NAND2_990( .ZN(g19121), .A1(g16682), .A2(g16697) );
  NAND2_X1 NAND2_991( .ZN(g19128), .A1(g16708), .A2(g16728) );
  NAND2_X1 NAND2_992( .ZN(g19135), .A1(g16739), .A2(g16770) );
  NAND2_X1 NAND2_993( .ZN(g19138), .A1(g16781), .A2(g16797) );
  NAND2_X1 NAND2_994( .ZN(g19141), .A1(g3088), .A2(g16825) );
  NAND2_X1 NAND2_995( .ZN(g19152), .A1(g5378), .A2(g18884) );
  NAND2_X1 NAND2_996( .ZN(II25532), .A1(g52), .A2(g18179) );
  NAND2_X1 NAND2_997( .ZN(II25533), .A1(g52), .A2(II25532) );
  NAND2_X1 NAND2_998( .ZN(II25534), .A1(g18179), .A2(II25532) );
  NAND2_X1 NAND2_999( .ZN(g19261), .A1(II25533), .A2(II25534) );
  NAND2_X1 NAND2_1000( .ZN(II25539), .A1(g92), .A2(g18174) );
  NAND2_X1 NAND2_1001( .ZN(II25540), .A1(g92), .A2(II25539) );
  NAND2_X1 NAND2_1002( .ZN(II25541), .A1(g18174), .A2(II25539) );
  NAND2_X1 NAND2_1003( .ZN(g19262), .A1(II25540), .A2(II25541) );
  NAND2_X1 NAND2_1004( .ZN(II25560), .A1(g56), .A2(g17724) );
  NAND2_X1 NAND2_1005( .ZN(II25561), .A1(g56), .A2(II25560) );
  NAND2_X1 NAND2_1006( .ZN(II25562), .A1(g17724), .A2(II25560) );
  NAND2_X1 NAND2_1007( .ZN(g19271), .A1(II25561), .A2(II25562) );
  NAND2_X1 NAND2_1008( .ZN(II25571), .A1(g740), .A2(g18286) );
  NAND2_X1 NAND2_1009( .ZN(II25572), .A1(g740), .A2(II25571) );
  NAND2_X1 NAND2_1010( .ZN(II25573), .A1(g18286), .A2(II25571) );
  NAND2_X1 NAND2_1011( .ZN(g19276), .A1(II25572), .A2(II25573) );
  NAND2_X1 NAND2_1012( .ZN(II25578), .A1(g780), .A2(g18281) );
  NAND2_X1 NAND2_1013( .ZN(II25579), .A1(g780), .A2(II25578) );
  NAND2_X1 NAND2_1014( .ZN(II25580), .A1(g18281), .A2(II25578) );
  NAND2_X1 NAND2_1015( .ZN(g19277), .A1(II25579), .A2(II25580) );
  NAND2_X1 NAND2_1016( .ZN(II25595), .A1(g61), .A2(g18074) );
  NAND2_X1 NAND2_1017( .ZN(II25596), .A1(g61), .A2(II25595) );
  NAND2_X1 NAND2_1018( .ZN(II25597), .A1(g18074), .A2(II25595) );
  NAND2_X1 NAND2_1019( .ZN(g19286), .A1(II25596), .A2(II25597) );
  NAND3_X1 NAND3_8( .ZN(g19288), .A1(g14685), .A2(g8580), .A3(g17057) );
  NAND2_X1 NAND2_1020( .ZN(II25605), .A1(g744), .A2(g17825) );
  NAND2_X1 NAND2_1021( .ZN(II25606), .A1(g744), .A2(II25605) );
  NAND2_X1 NAND2_1022( .ZN(II25607), .A1(g17825), .A2(II25605) );
  NAND2_X1 NAND2_1023( .ZN(g19290), .A1(II25606), .A2(II25607) );
  NAND2_X1 NAND2_1024( .ZN(II25616), .A1(g1426), .A2(g18379) );
  NAND2_X1 NAND2_1025( .ZN(II25617), .A1(g1426), .A2(II25616) );
  NAND2_X1 NAND2_1026( .ZN(II25618), .A1(g18379), .A2(II25616) );
  NAND2_X1 NAND2_1027( .ZN(g19295), .A1(II25617), .A2(II25618) );
  NAND2_X1 NAND2_1028( .ZN(II25623), .A1(g1466), .A2(g18374) );
  NAND2_X1 NAND2_1029( .ZN(II25624), .A1(g1466), .A2(II25623) );
  NAND2_X1 NAND2_1030( .ZN(II25625), .A1(g18374), .A2(II25623) );
  NAND2_X1 NAND2_1031( .ZN(g19296), .A1(II25624), .A2(II25625) );
  NAND2_X1 NAND2_1032( .ZN(II25633), .A1(g65), .A2(g17640) );
  NAND2_X1 NAND2_1033( .ZN(II25634), .A1(g65), .A2(II25633) );
  NAND2_X1 NAND2_1034( .ZN(II25635), .A1(g17640), .A2(II25633) );
  NAND2_X1 NAND2_1035( .ZN(g19300), .A1(II25634), .A2(II25635) );
  NAND2_X1 NAND2_1036( .ZN(II25643), .A1(g749), .A2(g18190) );
  NAND2_X1 NAND2_1037( .ZN(II25644), .A1(g749), .A2(II25643) );
  NAND2_X1 NAND2_1038( .ZN(II25645), .A1(g18190), .A2(II25643) );
  NAND2_X1 NAND2_1039( .ZN(g19304), .A1(II25644), .A2(II25645) );
  NAND3_X1 NAND3_9( .ZN(g19306), .A1(g14719), .A2(g8587), .A3(g17092) );
  NAND2_X1 NAND2_1040( .ZN(II25653), .A1(g1430), .A2(g17937) );
  NAND2_X1 NAND2_1041( .ZN(II25654), .A1(g1430), .A2(II25653) );
  NAND2_X1 NAND2_1042( .ZN(II25655), .A1(g17937), .A2(II25653) );
  NAND2_X1 NAND2_1043( .ZN(g19308), .A1(II25654), .A2(II25655) );
  NAND2_X1 NAND2_1044( .ZN(II25664), .A1(g2120), .A2(g18474) );
  NAND2_X1 NAND2_1045( .ZN(II25665), .A1(g2120), .A2(II25664) );
  NAND2_X1 NAND2_1046( .ZN(II25666), .A1(g18474), .A2(II25664) );
  NAND2_X1 NAND2_1047( .ZN(g19313), .A1(II25665), .A2(II25666) );
  NAND2_X1 NAND2_1048( .ZN(II25671), .A1(g2160), .A2(g18469) );
  NAND2_X1 NAND2_1049( .ZN(II25672), .A1(g2160), .A2(II25671) );
  NAND2_X1 NAND2_1050( .ZN(II25673), .A1(g18469), .A2(II25671) );
  NAND2_X1 NAND2_1051( .ZN(g19314), .A1(II25672), .A2(II25673) );
  NAND2_X1 NAND2_1052( .ZN(II25681), .A1(g70), .A2(g17974) );
  NAND2_X1 NAND2_1053( .ZN(II25682), .A1(g70), .A2(II25681) );
  NAND2_X1 NAND2_1054( .ZN(II25683), .A1(g17974), .A2(II25681) );
  NAND2_X1 NAND2_1055( .ZN(g19318), .A1(II25682), .A2(II25683) );
  NAND2_X1 NAND2_1056( .ZN(II25690), .A1(g753), .A2(g17741) );
  NAND2_X1 NAND2_1057( .ZN(II25691), .A1(g753), .A2(II25690) );
  NAND2_X1 NAND2_1058( .ZN(II25692), .A1(g17741), .A2(II25690) );
  NAND2_X1 NAND2_1059( .ZN(g19321), .A1(II25691), .A2(II25692) );
  NAND2_X1 NAND2_1060( .ZN(II25700), .A1(g1435), .A2(g18297) );
  NAND2_X1 NAND2_1061( .ZN(II25701), .A1(g1435), .A2(II25700) );
  NAND2_X1 NAND2_1062( .ZN(II25702), .A1(g18297), .A2(II25700) );
  NAND2_X1 NAND2_1063( .ZN(g19325), .A1(II25701), .A2(II25702) );
  NAND3_X1 NAND3_10( .ZN(g19327), .A1(g14747), .A2(g8594), .A3(g17130) );
  NAND2_X1 NAND2_1064( .ZN(II25710), .A1(g2124), .A2(g18048) );
  NAND2_X1 NAND2_1065( .ZN(II25711), .A1(g2124), .A2(II25710) );
  NAND2_X1 NAND2_1066( .ZN(II25712), .A1(g18048), .A2(II25710) );
  NAND2_X1 NAND2_1067( .ZN(g19329), .A1(II25711), .A2(II25712) );
  NAND2_X1 NAND2_1068( .ZN(II25721), .A1(g74), .A2(g18341) );
  NAND2_X1 NAND2_1069( .ZN(II25722), .A1(g74), .A2(II25721) );
  NAND2_X1 NAND2_1070( .ZN(II25723), .A1(g18341), .A2(II25721) );
  NAND2_X1 NAND2_1071( .ZN(g19334), .A1(II25722), .A2(II25723) );
  NAND2_X1 NAND2_1072( .ZN(II25731), .A1(g758), .A2(g18091) );
  NAND2_X1 NAND2_1073( .ZN(II25732), .A1(g758), .A2(II25731) );
  NAND2_X1 NAND2_1074( .ZN(II25733), .A1(g18091), .A2(II25731) );
  NAND2_X1 NAND2_1075( .ZN(g19345), .A1(II25732), .A2(II25733) );
  NAND2_X1 NAND2_1076( .ZN(II25740), .A1(g1439), .A2(g17842) );
  NAND2_X1 NAND2_1077( .ZN(II25741), .A1(g1439), .A2(II25740) );
  NAND2_X1 NAND2_1078( .ZN(II25742), .A1(g17842), .A2(II25740) );
  NAND2_X1 NAND2_1079( .ZN(g19348), .A1(II25741), .A2(II25742) );
  NAND2_X1 NAND2_1080( .ZN(II25750), .A1(g2129), .A2(g18390) );
  NAND2_X1 NAND2_1081( .ZN(II25751), .A1(g2129), .A2(II25750) );
  NAND2_X1 NAND2_1082( .ZN(II25752), .A1(g18390), .A2(II25750) );
  NAND2_X1 NAND2_1083( .ZN(g19352), .A1(II25751), .A2(II25752) );
  NAND3_X1 NAND3_11( .ZN(g19354), .A1(g14768), .A2(g8605), .A3(g17157) );
  NAND2_X1 NAND2_1084( .ZN(II25761), .A1(g79), .A2(g17882) );
  NAND2_X1 NAND2_1085( .ZN(II25762), .A1(g79), .A2(II25761) );
  NAND2_X1 NAND2_1086( .ZN(II25763), .A1(g17882), .A2(II25761) );
  NAND2_X1 NAND2_1087( .ZN(g19357), .A1(II25762), .A2(II25763) );
  NAND2_X1 NAND2_1088( .ZN(II25771), .A1(g762), .A2(g18436) );
  NAND2_X1 NAND2_1089( .ZN(II25772), .A1(g762), .A2(II25771) );
  NAND2_X1 NAND2_1090( .ZN(II25773), .A1(g18436), .A2(II25771) );
  NAND2_X1 NAND2_1091( .ZN(g19368), .A1(II25772), .A2(II25773) );
  NAND2_X1 NAND2_1092( .ZN(II25781), .A1(g1444), .A2(g18207) );
  NAND2_X2 NAND2_1093( .ZN(II25782), .A1(g1444), .A2(II25781) );
  NAND2_X1 NAND2_1094( .ZN(II25783), .A1(g18207), .A2(II25781) );
  NAND2_X1 NAND2_1095( .ZN(g19379), .A1(II25782), .A2(II25783) );
  NAND2_X1 NAND2_1096( .ZN(II25790), .A1(g2133), .A2(g17954) );
  NAND2_X1 NAND2_1097( .ZN(II25791), .A1(g2133), .A2(II25790) );
  NAND2_X1 NAND2_1098( .ZN(II25792), .A1(g17954), .A2(II25790) );
  NAND2_X1 NAND2_1099( .ZN(g19382), .A1(II25791), .A2(II25792) );
  NAND2_X1 NAND2_1100( .ZN(II25800), .A1(g83), .A2(g18265) );
  NAND2_X1 NAND2_1101( .ZN(II25801), .A1(g83), .A2(II25800) );
  NAND2_X1 NAND2_1102( .ZN(II25802), .A1(g18265), .A2(II25800) );
  NAND2_X1 NAND2_1103( .ZN(g19386), .A1(II25801), .A2(II25802) );
  NAND2_X1 NAND2_1104( .ZN(II25809), .A1(g767), .A2(g17993) );
  NAND2_X1 NAND2_1105( .ZN(II25810), .A1(g767), .A2(II25809) );
  NAND2_X1 NAND2_1106( .ZN(II25811), .A1(g17993), .A2(II25809) );
  NAND2_X1 NAND2_1107( .ZN(g19389), .A1(II25810), .A2(II25811) );
  NAND2_X1 NAND2_1108( .ZN(II25819), .A1(g1448), .A2(g18509) );
  NAND2_X1 NAND2_1109( .ZN(II25820), .A1(g1448), .A2(II25819) );
  NAND2_X1 NAND2_1110( .ZN(II25821), .A1(g18509), .A2(II25819) );
  NAND2_X1 NAND2_1111( .ZN(g19400), .A1(II25820), .A2(II25821) );
  NAND2_X1 NAND2_1112( .ZN(II25829), .A1(g2138), .A2(g18314) );
  NAND2_X1 NAND2_1113( .ZN(II25830), .A1(g2138), .A2(II25829) );
  NAND2_X1 NAND2_1114( .ZN(II25831), .A1(g18314), .A2(II25829) );
  NAND2_X1 NAND2_1115( .ZN(g19411), .A1(II25830), .A2(II25831) );
  NAND2_X1 NAND2_1116( .ZN(II25838), .A1(g88), .A2(g17802) );
  NAND2_X1 NAND2_1117( .ZN(II25839), .A1(g88), .A2(II25838) );
  NAND2_X1 NAND2_1118( .ZN(II25840), .A1(g17802), .A2(II25838) );
  NAND2_X1 NAND2_1119( .ZN(g19414), .A1(II25839), .A2(II25840) );
  NAND2_X1 NAND2_1120( .ZN(II25846), .A1(g771), .A2(g18358) );
  NAND2_X1 NAND2_1121( .ZN(II25847), .A1(g771), .A2(II25846) );
  NAND2_X1 NAND2_1122( .ZN(II25848), .A1(g18358), .A2(II25846) );
  NAND2_X1 NAND2_1123( .ZN(g19416), .A1(II25847), .A2(II25848) );
  NAND2_X1 NAND2_1124( .ZN(II25855), .A1(g1453), .A2(g18110) );
  NAND2_X1 NAND2_1125( .ZN(II25856), .A1(g1453), .A2(II25855) );
  NAND2_X1 NAND2_1126( .ZN(II25857), .A1(g18110), .A2(II25855) );
  NAND2_X1 NAND2_1127( .ZN(g19419), .A1(II25856), .A2(II25857) );
  NAND2_X1 NAND2_1128( .ZN(II25865), .A1(g2142), .A2(g18573) );
  NAND2_X1 NAND2_1129( .ZN(II25866), .A1(g2142), .A2(II25865) );
  NAND2_X1 NAND2_1130( .ZN(II25867), .A1(g18573), .A2(II25865) );
  NAND2_X1 NAND2_1131( .ZN(g19430), .A1(II25866), .A2(II25867) );
  NAND2_X1 NAND2_1132( .ZN(II25880), .A1(g776), .A2(g17914) );
  NAND2_X1 NAND2_1133( .ZN(II25881), .A1(g776), .A2(II25880) );
  NAND2_X1 NAND2_1134( .ZN(II25882), .A1(g17914), .A2(II25880) );
  NAND2_X1 NAND2_1135( .ZN(g19451), .A1(II25881), .A2(II25882) );
  NAND2_X1 NAND2_1136( .ZN(II25888), .A1(g1457), .A2(g18453) );
  NAND2_X1 NAND2_1137( .ZN(II25889), .A1(g1457), .A2(II25888) );
  NAND2_X1 NAND2_1138( .ZN(II25890), .A1(g18453), .A2(II25888) );
  NAND2_X1 NAND2_1139( .ZN(g19453), .A1(II25889), .A2(II25890) );
  NAND2_X1 NAND2_1140( .ZN(II25897), .A1(g2147), .A2(g18226) );
  NAND2_X1 NAND2_1141( .ZN(II25898), .A1(g2147), .A2(II25897) );
  NAND2_X1 NAND2_1142( .ZN(II25899), .A1(g18226), .A2(II25897) );
  NAND2_X1 NAND2_1143( .ZN(g19456), .A1(II25898), .A2(II25899) );
  NAND2_X1 NAND2_1144( .ZN(II25913), .A1(g1462), .A2(g18025) );
  NAND2_X1 NAND2_1145( .ZN(II25914), .A1(g1462), .A2(II25913) );
  NAND2_X1 NAND2_1146( .ZN(II25915), .A1(g18025), .A2(II25913) );
  NAND2_X1 NAND2_1147( .ZN(g19478), .A1(II25914), .A2(II25915) );
  NAND2_X1 NAND2_1148( .ZN(II25921), .A1(g2151), .A2(g18526) );
  NAND2_X1 NAND2_1149( .ZN(II25922), .A1(g2151), .A2(II25921) );
  NAND2_X1 NAND2_1150( .ZN(II25923), .A1(g18526), .A2(II25921) );
  NAND2_X1 NAND2_1151( .ZN(g19480), .A1(II25922), .A2(II25923) );
  NAND2_X1 NAND2_1152( .ZN(II25938), .A1(g2156), .A2(g18142) );
  NAND2_X1 NAND2_1153( .ZN(II25939), .A1(g2156), .A2(II25938) );
  NAND2_X1 NAND2_1154( .ZN(II25940), .A1(g18142), .A2(II25938) );
  NAND2_X1 NAND2_1155( .ZN(g19501), .A1(II25939), .A2(II25940) );
  NAND2_X1 NAND2_1156( .ZN(g19865), .A1(g16607), .A2(g9636) );
  NAND2_X1 NAND2_1157( .ZN(g19896), .A1(g16625), .A2(g9782) );
  NAND2_X1 NAND2_1158( .ZN(g19921), .A1(g16639), .A2(g9928) );
  NAND2_X1 NAND2_1159( .ZN(g19936), .A1(g16650), .A2(g10082) );
  NAND2_X1 NAND2_1160( .ZN(g19954), .A1(g17186), .A2(g92) );
  NAND2_X1 NAND2_1161( .ZN(g19984), .A1(g17197), .A2(g780) );
  NAND2_X1 NAND2_1162( .ZN(g20022), .A1(g17204), .A2(g1466) );
  NAND2_X1 NAND2_1163( .ZN(g20064), .A1(g17209), .A2(g2160) );
  NAND2_X1 NAND2_1164( .ZN(g20473), .A1(g18085), .A2(g646) );
  NAND2_X1 NAND2_1165( .ZN(g20481), .A1(g18201), .A2(g1332) );
  NAND2_X1 NAND2_1166( .ZN(g20487), .A1(g18308), .A2(g2026) );
  NAND2_X1 NAND2_1167( .ZN(g20493), .A1(g18401), .A2(g2720) );
  NAND2_X1 NAND2_1168( .ZN(g20497), .A1(g5410), .A2(g18886) );
  NAND2_X1 NAND2_1169( .ZN(g20522), .A1(g16501), .A2(g16515) );
  NAND2_X1 NAND2_1170( .ZN(g20537), .A1(g18626), .A2(g3036) );
  NAND2_X1 NAND2_1171( .ZN(g20542), .A1(g16523), .A2(g16546) );
  NAND2_X1 NAND2_1172( .ZN(g20633), .A1(g20164), .A2(g3254) );
  NAND2_X1 NAND2_1173( .ZN(g20648), .A1(g20164), .A2(g3254) );
  NAND2_X1 NAND2_1174( .ZN(g20658), .A1(g20198), .A2(g3410) );
  NAND2_X1 NAND2_1175( .ZN(g20672), .A1(g20164), .A2(g3254) );
  NAND2_X1 NAND2_1176( .ZN(g20683), .A1(g20198), .A2(g3410) );
  NAND2_X1 NAND2_1177( .ZN(g20693), .A1(g20228), .A2(g3566) );
  NAND2_X1 NAND2_1178( .ZN(g20700), .A1(g20153), .A2(g2903) );
  NAND2_X1 NAND2_1179( .ZN(g20703), .A1(g20164), .A2(g3254) );
  NAND2_X1 NAND2_1180( .ZN(g20707), .A1(g20198), .A2(g3410) );
  NAND2_X1 NAND2_1181( .ZN(g20718), .A1(g20228), .A2(g3566) );
  NAND2_X1 NAND2_1182( .ZN(g20728), .A1(g20255), .A2(g3722) );
  NAND2_X1 NAND2_1183( .ZN(g20738), .A1(g20198), .A2(g3410) );
  NAND2_X1 NAND2_1184( .ZN(g20742), .A1(g20228), .A2(g3566) );
  NAND2_X1 NAND2_1185( .ZN(g20753), .A1(g20255), .A2(g3722) );
  NAND2_X1 NAND2_1186( .ZN(g20775), .A1(g20228), .A2(g3566) );
  NAND2_X1 NAND2_1187( .ZN(g20779), .A1(g20255), .A2(g3722) );
  NAND2_X1 NAND2_1188( .ZN(g20805), .A1(g20255), .A2(g3722) );
  NAND2_X1 NAND2_1189( .ZN(g20825), .A1(g19219), .A2(g15959) );
  NAND2_X1 NAND2_1190( .ZN(g21659), .A1(g20164), .A2(g6314) );
  NAND2_X1 NAND2_1191( .ZN(II28189), .A1(g14079), .A2(g19444) );
  NAND2_X1 NAND2_1192( .ZN(II28190), .A1(g14079), .A2(II28189) );
  NAND2_X1 NAND2_1193( .ZN(II28191), .A1(g19444), .A2(II28189) );
  NAND2_X1 NAND2_1194( .ZN(g21660), .A1(II28190), .A2(II28191) );
  NAND2_X1 NAND2_1195( .ZN(g21685), .A1(g20164), .A2(g6232) );
  NAND2_X1 NAND2_1196( .ZN(g21686), .A1(g20164), .A2(g6314) );
  NAND2_X1 NAND2_1197( .ZN(g21688), .A1(g20198), .A2(g6519) );
  NAND2_X1 NAND2_1198( .ZN(II28217), .A1(g14194), .A2(g19471) );
  NAND2_X1 NAND2_1199( .ZN(II28218), .A1(g14194), .A2(II28217) );
  NAND2_X1 NAND2_1200( .ZN(II28219), .A1(g19471), .A2(II28217) );
  NAND2_X1 NAND2_1201( .ZN(g21689), .A1(II28218), .A2(II28219) );
  NAND2_X1 NAND2_1202( .ZN(g21714), .A1(g20164), .A2(g6232) );
  NAND2_X1 NAND2_1203( .ZN(g21715), .A1(g20164), .A2(g6314) );
  NAND4_X1 NAND4_1( .ZN(g21720), .A1(g14256), .A2(g15177), .A3(g19871), .A4(g19842) );
  NAND2_X1 NAND2_1204( .ZN(g21721), .A1(g20198), .A2(g6369) );
  NAND2_X1 NAND2_1205( .ZN(g21722), .A1(g20198), .A2(g6519) );
  NAND2_X1 NAND2_1206( .ZN(g21724), .A1(g20228), .A2(g6783) );
  NAND2_X1 NAND2_1207( .ZN(II28247), .A1(g14309), .A2(g19494) );
  NAND2_X1 NAND2_1208( .ZN(II28248), .A1(g14309), .A2(II28247) );
  NAND2_X2 NAND2_1209( .ZN(II28249), .A1(g19494), .A2(II28247) );
  NAND2_X2 NAND2_1210( .ZN(g21725), .A1(II28248), .A2(II28249) );
  NAND2_X1 NAND2_1211( .ZN(g21736), .A1(g20164), .A2(g6232) );
  NAND2_X1 NAND2_1212( .ZN(g21737), .A1(g20164), .A2(g6314) );
  NAND2_X1 NAND2_1213( .ZN(g21740), .A1(g20198), .A2(g6369) );
  NAND2_X1 NAND2_1214( .ZN(g21741), .A1(g20198), .A2(g6519) );
  NAND4_X1 NAND4_2( .ZN(g21746), .A1(g14378), .A2(g15263), .A3(g19902), .A4(g19875) );
  NAND2_X1 NAND2_1215( .ZN(g21747), .A1(g20228), .A2(g6574) );
  NAND2_X1 NAND2_1216( .ZN(g21748), .A1(g20228), .A2(g6783) );
  NAND2_X1 NAND2_1217( .ZN(g21750), .A1(g20255), .A2(g7085) );
  NAND2_X1 NAND2_1218( .ZN(II28271), .A1(g14431), .A2(g19515) );
  NAND2_X1 NAND2_1219( .ZN(II28272), .A1(g14431), .A2(II28271) );
  NAND2_X1 NAND2_1220( .ZN(II28273), .A1(g19515), .A2(II28271) );
  NAND2_X1 NAND2_1221( .ZN(g21751), .A1(II28272), .A2(II28273) );
  NAND2_X1 NAND2_1222( .ZN(g21759), .A1(g20164), .A2(g6232) );
  NAND2_X1 NAND2_1223( .ZN(g21760), .A1(g20198), .A2(g6369) );
  NAND2_X1 NAND2_1224( .ZN(g21761), .A1(g20198), .A2(g6519) );
  NAND2_X1 NAND2_1225( .ZN(g21764), .A1(g20228), .A2(g6574) );
  NAND2_X1 NAND2_1226( .ZN(g21765), .A1(g20228), .A2(g6783) );
  NAND4_X1 NAND4_3( .ZN(g21770), .A1(g14490), .A2(g15355), .A3(g19927), .A4(g19906) );
  NAND2_X1 NAND2_1227( .ZN(g21771), .A1(g20255), .A2(g6838) );
  NAND2_X1 NAND2_1228( .ZN(g21772), .A1(g20255), .A2(g7085) );
  NAND2_X1 NAND2_1229( .ZN(g21775), .A1(g20198), .A2(g6369) );
  NAND2_X1 NAND2_1230( .ZN(g21776), .A1(g20228), .A2(g6574) );
  NAND2_X1 NAND2_1231( .ZN(g21777), .A1(g20228), .A2(g6783) );
  NAND2_X1 NAND2_1232( .ZN(g21780), .A1(g20255), .A2(g6838) );
  NAND2_X1 NAND2_1233( .ZN(g21781), .A1(g20255), .A2(g7085) );
  NAND4_X1 NAND4_4( .ZN(g21786), .A1(g14577), .A2(g15441), .A3(g19942), .A4(g19931) );
  NAND2_X1 NAND2_1234( .ZN(g21790), .A1(g20228), .A2(g6574) );
  NAND2_X1 NAND2_1235( .ZN(g21791), .A1(g20255), .A2(g6838) );
  NAND2_X1 NAND2_1236( .ZN(g21792), .A1(g20255), .A2(g7085) );
  NAND2_X1 NAND2_1237( .ZN(g21804), .A1(g20255), .A2(g6838) );
  NAND3_X1 NAND3_12( .ZN(g21848), .A1(g17807), .A2(g19181), .A3(g19186) );
  NAND3_X1 NAND3_13( .ZN(g21850), .A1(g17979), .A2(g19187), .A3(g19191) );
  NAND3_X1 NAND3_14( .ZN(g21855), .A1(g17919), .A2(g19188), .A3(g19193) );
  NAND3_X1 NAND3_15( .ZN(g21857), .A1(g18079), .A2(g19192), .A3(g19200) );
  NAND3_X1 NAND3_16( .ZN(g21858), .A1(g18096), .A2(g19194), .A3(g19202) );
  NAND3_X1 NAND3_17( .ZN(g21859), .A1(g18030), .A2(g19195), .A3(g19204) );
  NAND3_X1 NAND3_18( .ZN(g21860), .A1(g18270), .A2(g19201), .A3(g19209) );
  NAND3_X1 NAND3_19( .ZN(g21862), .A1(g18195), .A2(g19203), .A3(g19211) );
  NAND3_X1 NAND3_20( .ZN(g21863), .A1(g18212), .A2(g19205), .A3(g19213) );
  NAND3_X1 NAND3_21( .ZN(g21864), .A1(g18147), .A2(g19206), .A3(g19215) );
  NAND3_X1 NAND3_22( .ZN(g21865), .A1(g18424), .A2(g19210), .A3(g19221) );
  NAND3_X1 NAND3_23( .ZN(g21866), .A1(g18363), .A2(g19212), .A3(g19222) );
  NAND3_X1 NAND3_24( .ZN(g21868), .A1(g18302), .A2(g19214), .A3(g19224) );
  NAND3_X1 NAND3_25( .ZN(g21869), .A1(g18319), .A2(g19216), .A3(g19226) );
  NAND3_X1 NAND3_26( .ZN(g21870), .A1(g18497), .A2(g19223), .A3(g19231) );
  NAND3_X1 NAND3_27( .ZN(g21871), .A1(g18458), .A2(g19225), .A3(g19232) );
  NAND3_X1 NAND3_28( .ZN(g21873), .A1(g18395), .A2(g19227), .A3(g19234) );
  NAND3_X1 NAND3_29( .ZN(g21874), .A1(g18561), .A2(g19233), .A3(g19244) );
  NAND3_X1 NAND3_30( .ZN(g21875), .A1(g18531), .A2(g19235), .A3(g19245) );
  NAND3_X1 NAND3_31( .ZN(g21877), .A1(g18611), .A2(g19246), .A3(g19257) );
  NAND3_X1 NAND3_32( .ZN(g21879), .A1(g18419), .A2(g19250), .A3(g19263) );
  NAND3_X1 NAND3_33( .ZN(g21881), .A1(g18492), .A2(g19264), .A3(g19278) );
  NAND3_X1 NAND3_34( .ZN(g21885), .A1(g18556), .A2(g19279), .A3(g19297) );
  NAND3_X1 NAND3_35( .ZN(g21888), .A1(g18606), .A2(g19298), .A3(g19315) );
  NAND2_X1 NAND2_1238( .ZN(g21903), .A1(g20008), .A2(g3013) );
  NAND3_X1 NAND3_36( .ZN(g21976), .A1(g19242), .A2(g21120), .A3(g19275) );
  NAND3_X1 NAND3_37( .ZN(g21983), .A1(g19255), .A2(g21139), .A3(g19294) );
  NAND2_X1 NAND2_1239( .ZN(g21989), .A1(g21048), .A2(g18623) );
  NAND2_X1 NAND2_1240( .ZN(g21991), .A1(g21501), .A2(g21536) );
  NAND3_X1 NAND3_38( .ZN(g21996), .A1(g19268), .A2(g21159), .A3(g19312) );
  NAND2_X2 NAND2_1241( .ZN(g22002), .A1(g21065), .A2(g21711) );
  NAND2_X2 NAND2_1242( .ZN(g22005), .A1(g21540), .A2(g21572) );
  NAND3_X1 NAND3_39( .ZN(g22009), .A1(g19283), .A2(g21179), .A3(g19333) );
  NAND2_X1 NAND2_1243( .ZN(g22016), .A1(g21576), .A2(g21605) );
  NAND2_X1 NAND2_1244( .ZN(g22021), .A1(g21609), .A2(g21634) );
  NAND3_X1 NAND3_40( .ZN(g22050), .A1(g19450), .A2(g21244), .A3(g19503) );
  NAND3_X1 NAND3_41( .ZN(g22069), .A1(g19477), .A2(g21253), .A3(g19522) );
  NAND2_X1 NAND2_1245( .ZN(g22083), .A1(g21774), .A2(g21787) );
  NAND3_X1 NAND3_42( .ZN(g22093), .A1(g19500), .A2(g21261), .A3(g19532) );
  NAND2_X1 NAND2_1246( .ZN(g22108), .A1(g21789), .A2(g21801) );
  NAND3_X1 NAND3_43( .ZN(g22118), .A1(g19521), .A2(g21269), .A3(g19542) );
  NAND2_X1 NAND2_1247( .ZN(g22134), .A1(g21803), .A2(g21809) );
  NAND2_X1 NAND2_1248( .ZN(g22157), .A1(g21811), .A2(g21816) );
  NAND2_X1 NAND2_1249( .ZN(II28726), .A1(g21887), .A2(g13519) );
  NAND2_X1 NAND2_1250( .ZN(II28727), .A1(g21887), .A2(II28726) );
  NAND2_X1 NAND2_1251( .ZN(II28728), .A1(g13519), .A2(II28726) );
  NAND2_X1 NAND2_1252( .ZN(g22188), .A1(II28727), .A2(II28728) );
  NAND2_X1 NAND2_1253( .ZN(II28741), .A1(g21890), .A2(g13530) );
  NAND2_X1 NAND2_1254( .ZN(II28742), .A1(g21890), .A2(II28741) );
  NAND2_X1 NAND2_1255( .ZN(II28743), .A1(g13530), .A2(II28741) );
  NAND2_X1 NAND2_1256( .ZN(g22197), .A1(II28742), .A2(II28743) );
  NAND2_X1 NAND2_1257( .ZN(II28753), .A1(g21893), .A2(g13541) );
  NAND2_X1 NAND2_1258( .ZN(II28754), .A1(g21893), .A2(II28753) );
  NAND2_X1 NAND2_1259( .ZN(II28755), .A1(g13541), .A2(II28753) );
  NAND2_X1 NAND2_1260( .ZN(g22203), .A1(II28754), .A2(II28755) );
  NAND2_X1 NAND2_1261( .ZN(II28765), .A1(g21901), .A2(g13552) );
  NAND2_X1 NAND2_1262( .ZN(II28766), .A1(g21901), .A2(II28765) );
  NAND2_X1 NAND2_1263( .ZN(II28767), .A1(g13552), .A2(II28765) );
  NAND2_X1 NAND2_1264( .ZN(g22209), .A1(II28766), .A2(II28767) );
  NAND3_X1 NAND3_44( .ZN(g22317), .A1(g21152), .A2(g21241), .A3(g21136) );
  NAND3_X1 NAND3_45( .ZN(g22339), .A1(g14442), .A2(g21149), .A3(g10694) );
  NAND3_X1 NAND3_46( .ZN(g22342), .A1(g21172), .A2(g21249), .A3(g21156) );
  NAND3_X1 NAND3_47( .ZN(g22362), .A1(g14529), .A2(g21169), .A3(g10714) );
  NAND3_X1 NAND3_48( .ZN(g22365), .A1(g21192), .A2(g21258), .A3(g21176) );
  NAND3_X1 NAND3_49( .ZN(g22381), .A1(g21211), .A2(g14442), .A3(g10694) );
  NAND3_X1 NAND3_50( .ZN(g22382), .A1(g14584), .A2(g21189), .A3(g10735) );
  NAND3_X1 NAND3_51( .ZN(g22385), .A1(g21207), .A2(g21266), .A3(g21196) );
  NAND3_X1 NAND3_52( .ZN(g22396), .A1(g21219), .A2(g14529), .A3(g10714) );
  NAND3_X1 NAND3_53( .ZN(g22397), .A1(g14618), .A2(g21204), .A3(g10754) );
  NAND3_X1 NAND3_54( .ZN(g22399), .A1(g21230), .A2(g14584), .A3(g10735) );
  NAND3_X1 NAND3_55( .ZN(g22400), .A1(g21235), .A2(g14618), .A3(g10754) );
  NAND2_X1 NAND2_1265( .ZN(g22608), .A1(g20842), .A2(g20885) );
  NAND2_X1 NAND2_1266( .ZN(g22644), .A1(g20850), .A2(g20904) );
  NAND2_X1 NAND2_1267( .ZN(g22668), .A1(g16075), .A2(g21271) );
  NAND2_X1 NAND2_1268( .ZN(g22680), .A1(g20858), .A2(g20928) );
  NAND2_X1 NAND2_1269( .ZN(g22708), .A1(g16113), .A2(g21278) );
  NAND2_X1 NAND2_1270( .ZN(g22720), .A1(g20866), .A2(g20956) );
  NAND2_X1 NAND2_1271( .ZN(g22739), .A1(g16164), .A2(g21285) );
  NAND2_X1 NAND2_1272( .ZN(g22771), .A1(g16223), .A2(g21293) );
  NAND3_X1 NAND3_56( .ZN(g22809), .A1(g21850), .A2(g21848), .A3(g21879) );
  NAND3_X1 NAND3_57( .ZN(g22844), .A1(g21865), .A2(g21860), .A3(g21857) );
  NAND2_X1 NAND2_1273( .ZN(g22845), .A1(g19441), .A2(g20885) );
  NAND2_X1 NAND2_1274( .ZN(g22846), .A1(g8278), .A2(g21660) );
  NAND3_X1 NAND3_58( .ZN(g22850), .A1(g21858), .A2(g21855), .A3(g21881) );
  NAND2_X1 NAND2_1275( .ZN(g22876), .A1(g21238), .A2(g83) );
  NAND3_X1 NAND3_59( .ZN(g22879), .A1(g21870), .A2(g21866), .A3(g21862) );
  NAND2_X1 NAND2_1276( .ZN(g22880), .A1(g19468), .A2(g20904) );
  NAND2_X1 NAND2_1277( .ZN(g22881), .A1(g8287), .A2(g21689) );
  NAND3_X1 NAND3_60( .ZN(g22885), .A1(g21863), .A2(g21859), .A3(g21885) );
  NAND2_X1 NAND2_1278( .ZN(g22911), .A1(g21246), .A2(g771) );
  NAND3_X1 NAND3_61( .ZN(g22914), .A1(g21874), .A2(g21871), .A3(g21868) );
  NAND2_X1 NAND2_1279( .ZN(g22915), .A1(g19491), .A2(g20928) );
  NAND2_X1 NAND2_1280( .ZN(g22916), .A1(g8296), .A2(g21725) );
  NAND3_X1 NAND3_62( .ZN(g22920), .A1(g21869), .A2(g21864), .A3(g21888) );
  NAND2_X1 NAND2_1281( .ZN(g22936), .A1(g21255), .A2(g1457) );
  NAND3_X1 NAND3_63( .ZN(g22939), .A1(g21877), .A2(g21875), .A3(g21873) );
  NAND2_X1 NAND2_1282( .ZN(g22940), .A1(g19512), .A2(g20956) );
  NAND2_X1 NAND2_1283( .ZN(g22941), .A1(g8305), .A2(g21751) );
  NAND2_X1 NAND2_1284( .ZN(g22942), .A1(g21263), .A2(g2151) );
  NAND2_X1 NAND2_1285( .ZN(g22992), .A1(g21636), .A2(g672) );
  NAND2_X1 NAND2_1286( .ZN(g23003), .A1(g21667), .A2(g1358) );
  NAND2_X1 NAND2_1287( .ZN(g23017), .A1(g21696), .A2(g2052) );
  NAND2_X1 NAND2_1288( .ZN(g23033), .A1(g21732), .A2(g2746) );
  NAND2_X1 NAND2_1289( .ZN(g23320), .A1(g23066), .A2(g23051) );
  NAND2_X1 NAND2_1290( .ZN(g23325), .A1(g23080), .A2(g23070) );
  NAND2_X1 NAND2_1291( .ZN(g23331), .A1(g22999), .A2(g22174) );
  NAND2_X1 NAND2_1292( .ZN(g23335), .A1(g23096), .A2(g23083) );
  NAND2_X1 NAND2_1293( .ZN(g23340), .A1(g23013), .A2(g22189) );
  NAND2_X1 NAND2_1294( .ZN(g23344), .A1(g23113), .A2(g23099) );
  NAND2_X1 NAND2_1295( .ZN(g23349), .A1(g23029), .A2(g22198) );
  NAND2_X1 NAND2_1296( .ZN(g23353), .A1(g23046), .A2(g22204) );
  NAND2_X1 NAND2_1297( .ZN(g23360), .A1(g21980), .A2(g21975) );
  NAND2_X1 NAND2_1298( .ZN(g23364), .A1(g21987), .A2(g21981) );
  NAND2_X1 NAND2_1299( .ZN(g23368), .A1(g23135), .A2(g22288) );
  NAND2_X1 NAND2_1300( .ZN(g23372), .A1(g22000), .A2(g21988) );
  NAND2_X1 NAND2_1301( .ZN(g23376), .A1(g18435), .A2(g22812) );
  NAND2_X1 NAND2_1302( .ZN(g23377), .A1(g21968), .A2(g22308) );
  NAND2_X1 NAND2_1303( .ZN(g23381), .A1(g22013), .A2(g22001) );
  NAND2_X1 NAND2_1304( .ZN(g23387), .A1(g18508), .A2(g22852) );
  NAND2_X1 NAND2_1305( .ZN(g23388), .A1(g21971), .A2(g22336) );
  NAND2_X1 NAND2_1306( .ZN(g23394), .A1(g18572), .A2(g22887) );
  NAND2_X1 NAND2_1307( .ZN(g23395), .A1(g21973), .A2(g22361) );
  NAND2_X1 NAND2_1308( .ZN(g23402), .A1(g18622), .A2(g22922) );
  NAND3_X1 NAND3_64( .ZN(g23478), .A1(g22809), .A2(g14442), .A3(g10694) );
  NAND3_X1 NAND3_65( .ZN(g23486), .A1(g22844), .A2(g14442), .A3(g10694) );
  NAND3_X1 NAND3_66( .ZN(g23489), .A1(g22850), .A2(g14529), .A3(g10714) );
  NAND3_X1 NAND3_67( .ZN(g23495), .A1(g10694), .A2(g14442), .A3(g22316) );
  NAND3_X1 NAND3_68( .ZN(g23502), .A1(g22879), .A2(g14529), .A3(g10714) );
  NAND3_X1 NAND3_69( .ZN(g23505), .A1(g22885), .A2(g14584), .A3(g10735) );
  NAND3_X1 NAND3_70( .ZN(g23511), .A1(g10714), .A2(g14529), .A3(g22341) );
  NAND3_X1 NAND3_71( .ZN(g23518), .A1(g22914), .A2(g14584), .A3(g10735) );
  NAND3_X1 NAND3_72( .ZN(g23521), .A1(g22920), .A2(g14618), .A3(g10754) );
  NAND3_X1 NAND3_73( .ZN(g23526), .A1(g10735), .A2(g14584), .A3(g22364) );
  NAND3_X1 NAND3_74( .ZN(g23533), .A1(g22939), .A2(g14618), .A3(g10754) );
  NAND3_X1 NAND3_75( .ZN(g23537), .A1(g10754), .A2(g14618), .A3(g22384) );
  NAND2_X1 NAND2_1309( .ZN(II30790), .A1(g22846), .A2(g14079) );
  NAND2_X1 NAND2_1310( .ZN(II30791), .A1(g22846), .A2(II30790) );
  NAND2_X1 NAND2_1311( .ZN(II30792), .A1(g14079), .A2(II30790) );
  NAND2_X1 NAND2_1312( .ZN(g23660), .A1(II30791), .A2(II30792) );
  NAND2_X1 NAND2_1313( .ZN(II30868), .A1(g22881), .A2(g14194) );
  NAND2_X1 NAND2_1314( .ZN(II30869), .A1(g22881), .A2(II30868) );
  NAND2_X1 NAND2_1315( .ZN(II30870), .A1(g14194), .A2(II30868) );
  NAND2_X1 NAND2_1316( .ZN(g23710), .A1(II30869), .A2(II30870) );
  NAND2_X1 NAND2_1317( .ZN(II30952), .A1(g22916), .A2(g14309) );
  NAND2_X1 NAND2_1318( .ZN(II30953), .A1(g22916), .A2(II30952) );
  NAND2_X1 NAND2_1319( .ZN(II30954), .A1(g14309), .A2(II30952) );
  NAND2_X1 NAND2_1320( .ZN(g23764), .A1(II30953), .A2(II30954) );
  NAND2_X1 NAND2_1321( .ZN(II31035), .A1(g22941), .A2(g14431) );
  NAND2_X1 NAND2_1322( .ZN(II31036), .A1(g22941), .A2(II31035) );
  NAND2_X1 NAND2_1323( .ZN(II31037), .A1(g14431), .A2(II31035) );
  NAND2_X1 NAND2_1324( .ZN(g23819), .A1(II31036), .A2(II31037) );
  NAND2_X1 NAND2_1325( .ZN(g23906), .A1(g22812), .A2(g13958) );
  NAND2_X1 NAND2_1326( .ZN(g23936), .A1(g22812), .A2(g13922) );
  NAND2_X1 NAND2_1327( .ZN(g23937), .A1(g22812), .A2(g13918) );
  NAND2_X1 NAND2_1328( .ZN(g23938), .A1(g22852), .A2(g14028) );
  NAND2_X1 NAND2_1329( .ZN(g23953), .A1(g22812), .A2(g14525) );
  NAND2_X1 NAND2_1330( .ZN(g23968), .A1(g22852), .A2(g13978) );
  NAND2_X1 NAND2_1331( .ZN(g23969), .A1(g22852), .A2(g13974) );
  NAND2_X1 NAND2_1332( .ZN(g23970), .A1(g22887), .A2(g14119) );
  NAND2_X1 NAND2_1333( .ZN(g23973), .A1(g22812), .A2(g14450) );
  NAND2_X1 NAND2_1334( .ZN(g23982), .A1(g22852), .A2(g14580) );
  NAND2_X1 NAND2_1335( .ZN(g23997), .A1(g22887), .A2(g14048) );
  NAND2_X1 NAND2_1336( .ZN(g23998), .A1(g22887), .A2(g14044) );
  NAND2_X1 NAND2_1337( .ZN(g23999), .A1(g22922), .A2(g14234) );
  NAND2_X1 NAND2_1338( .ZN(g24002), .A1(g22812), .A2(g14355) );
  NAND2_X1 NAND2_1339( .ZN(g24003), .A1(g22852), .A2(g14537) );
  NAND2_X1 NAND2_1340( .ZN(g24012), .A1(g22887), .A2(g14614) );
  NAND2_X1 NAND2_1341( .ZN(g24027), .A1(g22922), .A2(g14139) );
  NAND2_X1 NAND2_1342( .ZN(g24028), .A1(g22922), .A2(g14135) );
  NAND2_X1 NAND2_1343( .ZN(g24034), .A1(g22812), .A2(g14252) );
  NAND2_X1 NAND2_1344( .ZN(g24036), .A1(g22852), .A2(g14467) );
  NAND2_X1 NAND2_1345( .ZN(g24037), .A1(g22887), .A2(g14592) );
  NAND2_X1 NAND2_1346( .ZN(g24046), .A1(g22922), .A2(g14637) );
  NAND2_X1 NAND2_1347( .ZN(g24052), .A1(g22812), .A2(g14171) );
  NAND2_X1 NAND2_1348( .ZN(g24054), .A1(g22852), .A2(g14374) );
  NAND2_X1 NAND2_1349( .ZN(g24056), .A1(g22887), .A2(g14554) );
  NAND2_X1 NAND2_1350( .ZN(g24057), .A1(g22922), .A2(g14626) );
  NAND2_X1 NAND2_1351( .ZN(g24058), .A1(g22812), .A2(g14086) );
  NAND2_X1 NAND2_1352( .ZN(g24065), .A1(g22852), .A2(g14286) );
  NAND2_X1 NAND2_1353( .ZN(g24067), .A1(g22887), .A2(g14486) );
  NAND2_X1 NAND2_1354( .ZN(g24069), .A1(g22922), .A2(g14609) );
  NAND2_X1 NAND2_1355( .ZN(g24070), .A1(g22812), .A2(g14011) );
  NAND2_X1 NAND2_1356( .ZN(g24071), .A1(g22852), .A2(g14201) );
  NAND2_X1 NAND2_1357( .ZN(g24078), .A1(g22887), .A2(g14408) );
  NAND2_X1 NAND2_1358( .ZN(g24080), .A1(g22922), .A2(g14573) );
  NAND2_X1 NAND2_1359( .ZN(g24081), .A1(g22852), .A2(g14102) );
  NAND2_X1 NAND2_1360( .ZN(g24082), .A1(g22887), .A2(g14316) );
  NAND2_X1 NAND2_1361( .ZN(g24089), .A1(g22922), .A2(g14520) );
  NAND2_X1 NAND2_1362( .ZN(g24090), .A1(g22887), .A2(g14217) );
  NAND2_X1 NAND2_1363( .ZN(g24091), .A1(g22922), .A2(g14438) );
  NAND2_X1 NAND2_1364( .ZN(g24093), .A1(g22922), .A2(g14332) );
  NAND2_X1 NAND2_1365( .ZN(g24100), .A1(g20885), .A2(g22175) );
  NAND2_X1 NAND2_1366( .ZN(g24109), .A1(g20904), .A2(g22190) );
  NAND2_X1 NAND2_1367( .ZN(g24126), .A1(g20928), .A2(g22199) );
  NAND2_X1 NAND2_1368( .ZN(g24145), .A1(g20956), .A2(g22205) );
  NAND2_X1 NAND2_1369( .ZN(g24442), .A1(g23644), .A2(g3306) );
  NAND2_X1 NAND2_1370( .ZN(g24443), .A1(g23644), .A2(g3306) );
  NAND2_X1 NAND2_1371( .ZN(g24444), .A1(g23694), .A2(g3462) );
  NAND2_X1 NAND2_1372( .ZN(g24447), .A1(g23644), .A2(g3306) );
  NAND2_X1 NAND2_1373( .ZN(g24448), .A1(g23923), .A2(g3338) );
  NAND2_X1 NAND2_1374( .ZN(g24449), .A1(g23694), .A2(g3462) );
  NAND2_X1 NAND2_1375( .ZN(g24450), .A1(g23748), .A2(g3618) );
  NAND2_X2 NAND2_1376( .ZN(g24451), .A1(g23644), .A2(g3306) );
  NAND2_X2 NAND2_1377( .ZN(g24452), .A1(g23923), .A2(g3338) );
  NAND2_X2 NAND2_1378( .ZN(g24453), .A1(g23694), .A2(g3462) );
  NAND2_X1 NAND2_1379( .ZN(g24454), .A1(g23955), .A2(g3494) );
  NAND2_X1 NAND2_1380( .ZN(g24455), .A1(g23748), .A2(g3618) );
  NAND2_X1 NAND2_1381( .ZN(g24456), .A1(g23803), .A2(g3774) );
  NAND2_X1 NAND2_1382( .ZN(g24457), .A1(g23923), .A2(g3338) );
  NAND2_X1 NAND2_1383( .ZN(g24458), .A1(g23694), .A2(g3462) );
  NAND2_X1 NAND2_1384( .ZN(g24459), .A1(g23955), .A2(g3494) );
  NAND2_X1 NAND2_1385( .ZN(g24460), .A1(g23748), .A2(g3618) );
  NAND2_X1 NAND2_1386( .ZN(g24461), .A1(g23984), .A2(g3650) );
  NAND2_X1 NAND2_1387( .ZN(g24462), .A1(g23803), .A2(g3774) );
  NAND2_X1 NAND2_1388( .ZN(g24463), .A1(g23923), .A2(g3338) );
  NAND2_X1 NAND2_1389( .ZN(g24464), .A1(g23955), .A2(g3494) );
  NAND2_X1 NAND2_1390( .ZN(g24465), .A1(g23748), .A2(g3618) );
  NAND2_X1 NAND2_1391( .ZN(g24466), .A1(g23984), .A2(g3650) );
  NAND2_X1 NAND2_1392( .ZN(g24467), .A1(g23803), .A2(g3774) );
  NAND2_X1 NAND2_1393( .ZN(g24468), .A1(g24014), .A2(g3806) );
  NAND2_X1 NAND2_1394( .ZN(g24469), .A1(g23955), .A2(g3494) );
  NAND2_X1 NAND2_1395( .ZN(g24470), .A1(g23984), .A2(g3650) );
  NAND2_X1 NAND2_1396( .ZN(g24471), .A1(g23803), .A2(g3774) );
  NAND2_X1 NAND2_1397( .ZN(g24472), .A1(g24014), .A2(g3806) );
  NAND2_X1 NAND2_1398( .ZN(g24474), .A1(g23984), .A2(g3650) );
  NAND2_X1 NAND2_1399( .ZN(g24475), .A1(g24014), .A2(g3806) );
  NAND2_X1 NAND2_1400( .ZN(g24477), .A1(g24014), .A2(g3806) );
  NAND2_X1 NAND2_1401( .ZN(g24616), .A1(g499), .A2(g23376) );
  NAND2_X1 NAND2_1402( .ZN(g24627), .A1(g1186), .A2(g23387) );
  NAND2_X1 NAND2_1403( .ZN(g24641), .A1(g1880), .A2(g23394) );
  NAND2_X1 NAND2_1404( .ZN(g24660), .A1(g2574), .A2(g23402) );
  NAND2_X1 NAND2_1405( .ZN(II32265), .A1(g17903), .A2(g23936) );
  NAND2_X1 NAND2_1406( .ZN(II32266), .A1(g17903), .A2(II32265) );
  NAND2_X1 NAND2_1407( .ZN(II32267), .A1(g23936), .A2(II32265) );
  NAND2_X1 NAND2_1408( .ZN(g24753), .A1(II32266), .A2(II32267) );
  NAND2_X1 NAND2_1409( .ZN(II32284), .A1(g17815), .A2(g23953) );
  NAND2_X1 NAND2_1410( .ZN(II32285), .A1(g17815), .A2(II32284) );
  NAND2_X1 NAND2_1411( .ZN(II32286), .A1(g23953), .A2(II32284) );
  NAND2_X1 NAND2_1412( .ZN(g24766), .A1(II32285), .A2(II32286) );
  NAND2_X1 NAND2_1413( .ZN(II32295), .A1(g18014), .A2(g23968) );
  NAND2_X1 NAND2_1414( .ZN(II32296), .A1(g18014), .A2(II32295) );
  NAND2_X1 NAND2_1415( .ZN(II32297), .A1(g23968), .A2(II32295) );
  NAND2_X1 NAND2_1416( .ZN(g24771), .A1(II32296), .A2(II32297) );
  NAND2_X1 NAND2_1417( .ZN(II32308), .A1(g17903), .A2(g23973) );
  NAND2_X1 NAND2_1418( .ZN(II32309), .A1(g17903), .A2(II32308) );
  NAND2_X1 NAND2_1419( .ZN(II32310), .A1(g23973), .A2(II32308) );
  NAND2_X1 NAND2_1420( .ZN(g24778), .A1(II32309), .A2(II32310) );
  NAND2_X1 NAND2_1421( .ZN(II32323), .A1(g17927), .A2(g23982) );
  NAND2_X1 NAND2_1422( .ZN(II32324), .A1(g17927), .A2(II32323) );
  NAND2_X1 NAND2_1423( .ZN(II32325), .A1(g23982), .A2(II32323) );
  NAND2_X1 NAND2_1424( .ZN(g24787), .A1(II32324), .A2(II32325) );
  NAND2_X1 NAND2_1425( .ZN(II32333), .A1(g18131), .A2(g23997) );
  NAND2_X1 NAND2_1426( .ZN(II32334), .A1(g18131), .A2(II32333) );
  NAND2_X1 NAND2_1427( .ZN(II32335), .A1(g23997), .A2(II32333) );
  NAND2_X1 NAND2_1428( .ZN(g24791), .A1(II32334), .A2(II32335) );
  NAND2_X1 NAND2_1429( .ZN(II32345), .A1(g17815), .A2(g24002) );
  NAND2_X1 NAND2_1430( .ZN(II32346), .A1(g17815), .A2(II32345) );
  NAND2_X1 NAND2_1431( .ZN(II32347), .A1(g24002), .A2(II32345) );
  NAND2_X1 NAND2_1432( .ZN(g24797), .A1(II32346), .A2(II32347) );
  NAND2_X1 NAND2_1433( .ZN(II32355), .A1(g18014), .A2(g24003) );
  NAND2_X1 NAND2_1434( .ZN(II32356), .A1(g18014), .A2(II32355) );
  NAND2_X1 NAND2_1435( .ZN(II32357), .A1(g24003), .A2(II32355) );
  NAND2_X1 NAND2_1436( .ZN(g24801), .A1(II32356), .A2(II32357) );
  NAND2_X1 NAND2_1437( .ZN(II32368), .A1(g18038), .A2(g24012) );
  NAND2_X1 NAND2_1438( .ZN(II32369), .A1(g18038), .A2(II32368) );
  NAND2_X1 NAND2_1439( .ZN(II32370), .A1(g24012), .A2(II32368) );
  NAND2_X1 NAND2_1440( .ZN(g24808), .A1(II32369), .A2(II32370) );
  NAND2_X1 NAND2_1441( .ZN(II32378), .A1(g18247), .A2(g24027) );
  NAND2_X1 NAND2_1442( .ZN(II32379), .A1(g18247), .A2(II32378) );
  NAND2_X1 NAND2_1443( .ZN(II32380), .A1(g24027), .A2(II32378) );
  NAND2_X1 NAND2_1444( .ZN(g24812), .A1(II32379), .A2(II32380) );
  NAND2_X1 NAND2_1445( .ZN(g24814), .A1(g24239), .A2(g24244) );
  NAND2_X1 NAND2_1446( .ZN(II32391), .A1(g17903), .A2(g24034) );
  NAND2_X1 NAND2_1447( .ZN(II32392), .A1(g17903), .A2(II32391) );
  NAND2_X1 NAND2_1448( .ZN(II32393), .A1(g24034), .A2(II32391) );
  NAND2_X1 NAND2_1449( .ZN(g24817), .A1(II32392), .A2(II32393) );
  NAND2_X1 NAND2_1450( .ZN(II32400), .A1(g17927), .A2(g24036) );
  NAND2_X1 NAND2_1451( .ZN(II32401), .A1(g17927), .A2(II32400) );
  NAND2_X1 NAND2_1452( .ZN(II32402), .A1(g24036), .A2(II32400) );
  NAND2_X1 NAND2_1453( .ZN(g24820), .A1(II32401), .A2(II32402) );
  NAND2_X1 NAND2_1454( .ZN(II32409), .A1(g18131), .A2(g24037) );
  NAND2_X1 NAND2_1455( .ZN(II32410), .A1(g18131), .A2(II32409) );
  NAND2_X1 NAND2_1456( .ZN(II32411), .A1(g24037), .A2(II32409) );
  NAND2_X1 NAND2_1457( .ZN(g24823), .A1(II32410), .A2(II32411) );
  NAND2_X1 NAND2_1458( .ZN(II32422), .A1(g18155), .A2(g24046) );
  NAND2_X1 NAND2_1459( .ZN(II32423), .A1(g18155), .A2(II32422) );
  NAND2_X1 NAND2_1460( .ZN(II32424), .A1(g24046), .A2(II32422) );
  NAND2_X1 NAND2_1461( .ZN(g24830), .A1(II32423), .A2(II32424) );
  NAND2_X1 NAND2_1462( .ZN(II32430), .A1(g17815), .A2(g24052) );
  NAND2_X1 NAND2_1463( .ZN(II32431), .A1(g17815), .A2(II32430) );
  NAND2_X1 NAND2_1464( .ZN(II32432), .A1(g24052), .A2(II32430) );
  NAND2_X1 NAND2_1465( .ZN(g24832), .A1(II32431), .A2(II32432) );
  NAND2_X1 NAND2_1466( .ZN(g24833), .A1(g24245), .A2(g24252) );
  NAND2_X1 NAND2_1467( .ZN(II32443), .A1(g18014), .A2(g24054) );
  NAND2_X1 NAND2_1468( .ZN(II32444), .A1(g18014), .A2(II32443) );
  NAND2_X1 NAND2_1469( .ZN(II32445), .A1(g24054), .A2(II32443) );
  NAND2_X1 NAND2_1470( .ZN(g24837), .A1(II32444), .A2(II32445) );
  NAND2_X1 NAND2_1471( .ZN(II32451), .A1(g18038), .A2(g24056) );
  NAND2_X1 NAND2_1472( .ZN(II32452), .A1(g18038), .A2(II32451) );
  NAND2_X1 NAND2_1473( .ZN(II32453), .A1(g24056), .A2(II32451) );
  NAND2_X1 NAND2_1474( .ZN(g24839), .A1(II32452), .A2(II32453) );
  NAND2_X1 NAND2_1475( .ZN(II32460), .A1(g18247), .A2(g24057) );
  NAND2_X1 NAND2_1476( .ZN(II32461), .A1(g18247), .A2(II32460) );
  NAND2_X1 NAND2_1477( .ZN(II32462), .A1(g24057), .A2(II32460) );
  NAND2_X1 NAND2_1478( .ZN(g24842), .A1(II32461), .A2(II32462) );
  NAND2_X1 NAND2_1479( .ZN(II32468), .A1(g17903), .A2(g24058) );
  NAND2_X1 NAND2_1480( .ZN(II32469), .A1(g17903), .A2(II32468) );
  NAND2_X1 NAND2_1481( .ZN(II32470), .A1(g24058), .A2(II32468) );
  NAND2_X1 NAND2_1482( .ZN(g24844), .A1(II32469), .A2(II32470) );
  NAND2_X1 NAND2_1483( .ZN(II32478), .A1(g17927), .A2(g24065) );
  NAND2_X1 NAND2_1484( .ZN(II32479), .A1(g17927), .A2(II32478) );
  NAND2_X1 NAND2_1485( .ZN(II32480), .A1(g24065), .A2(II32478) );
  NAND2_X1 NAND2_1486( .ZN(g24848), .A1(II32479), .A2(II32480) );
  NAND2_X1 NAND2_1487( .ZN(g24849), .A1(g24254), .A2(g24257) );
  NAND2_X1 NAND2_1488( .ZN(II32490), .A1(g18131), .A2(g24067) );
  NAND2_X1 NAND2_1489( .ZN(II32491), .A1(g18131), .A2(II32490) );
  NAND2_X2 NAND2_1490( .ZN(II32492), .A1(g24067), .A2(II32490) );
  NAND2_X2 NAND2_1491( .ZN(g24852), .A1(II32491), .A2(II32492) );
  NAND2_X2 NAND2_1492( .ZN(II32498), .A1(g18155), .A2(g24069) );
  NAND2_X1 NAND2_1493( .ZN(II32499), .A1(g18155), .A2(II32498) );
  NAND2_X1 NAND2_1494( .ZN(II32500), .A1(g24069), .A2(II32498) );
  NAND2_X1 NAND2_1495( .ZN(g24854), .A1(II32499), .A2(II32500) );
  NAND2_X1 NAND2_1496( .ZN(II32509), .A1(g17815), .A2(g24070) );
  NAND2_X1 NAND2_1497( .ZN(II32510), .A1(g17815), .A2(II32509) );
  NAND2_X1 NAND2_1498( .ZN(II32511), .A1(g24070), .A2(II32509) );
  NAND2_X1 NAND2_1499( .ZN(g24857), .A1(II32510), .A2(II32511) );
  NAND2_X1 NAND2_1500( .ZN(II32518), .A1(g18014), .A2(g24071) );
  NAND2_X1 NAND2_1501( .ZN(II32519), .A1(g18014), .A2(II32518) );
  NAND2_X1 NAND2_1502( .ZN(II32520), .A1(g24071), .A2(II32518) );
  NAND2_X1 NAND2_1503( .ZN(g24860), .A1(II32519), .A2(II32520) );
  NAND2_X1 NAND2_1504( .ZN(II32526), .A1(g18038), .A2(g24078) );
  NAND2_X1 NAND2_1505( .ZN(II32527), .A1(g18038), .A2(II32526) );
  NAND2_X1 NAND2_1506( .ZN(II32528), .A1(g24078), .A2(II32526) );
  NAND2_X1 NAND2_1507( .ZN(g24862), .A1(II32527), .A2(II32528) );
  NAND2_X1 NAND2_1508( .ZN(g24863), .A1(g24258), .A2(g23319) );
  NAND2_X1 NAND2_1509( .ZN(II32538), .A1(g18247), .A2(g24080) );
  NAND2_X1 NAND2_1510( .ZN(II32539), .A1(g18247), .A2(II32538) );
  NAND2_X1 NAND2_1511( .ZN(II32540), .A1(g24080), .A2(II32538) );
  NAND2_X1 NAND2_1512( .ZN(g24866), .A1(II32539), .A2(II32540) );
  NAND2_X1 NAND2_1513( .ZN(II32546), .A1(g17903), .A2(g23906) );
  NAND2_X1 NAND2_1514( .ZN(II32547), .A1(g17903), .A2(II32546) );
  NAND2_X1 NAND2_1515( .ZN(II32548), .A1(g23906), .A2(II32546) );
  NAND2_X1 NAND2_1516( .ZN(g24868), .A1(II32547), .A2(II32548) );
  NAND2_X1 NAND2_1517( .ZN(II32559), .A1(g17927), .A2(g24081) );
  NAND2_X1 NAND2_1518( .ZN(II32560), .A1(g17927), .A2(II32559) );
  NAND2_X1 NAND2_1519( .ZN(II32561), .A1(g24081), .A2(II32559) );
  NAND2_X1 NAND2_1520( .ZN(g24873), .A1(II32560), .A2(II32561) );
  NAND2_X1 NAND2_1521( .ZN(II32567), .A1(g18131), .A2(g24082) );
  NAND2_X1 NAND2_1522( .ZN(II32568), .A1(g18131), .A2(II32567) );
  NAND2_X1 NAND2_1523( .ZN(II32569), .A1(g24082), .A2(II32567) );
  NAND2_X1 NAND2_1524( .ZN(g24875), .A1(II32568), .A2(II32569) );
  NAND2_X1 NAND2_1525( .ZN(II32575), .A1(g18155), .A2(g24089) );
  NAND2_X1 NAND2_1526( .ZN(II32576), .A1(g18155), .A2(II32575) );
  NAND2_X1 NAND2_1527( .ZN(II32577), .A1(g24089), .A2(II32575) );
  NAND2_X1 NAND2_1528( .ZN(g24877), .A1(II32576), .A2(II32577) );
  NAND2_X1 NAND2_1529( .ZN(II32586), .A1(g17815), .A2(g23937) );
  NAND2_X1 NAND2_1530( .ZN(II32587), .A1(g17815), .A2(II32586) );
  NAND2_X1 NAND2_1531( .ZN(II32588), .A1(g23937), .A2(II32586) );
  NAND2_X1 NAND2_1532( .ZN(g24880), .A1(II32587), .A2(II32588) );
  NAND2_X1 NAND2_1533( .ZN(II32595), .A1(g18014), .A2(g23938) );
  NAND2_X1 NAND2_1534( .ZN(II32596), .A1(g18014), .A2(II32595) );
  NAND2_X1 NAND2_1535( .ZN(II32597), .A1(g23938), .A2(II32595) );
  NAND2_X1 NAND2_1536( .ZN(g24883), .A1(II32596), .A2(II32597) );
  NAND2_X1 NAND2_1537( .ZN(II32607), .A1(g18038), .A2(g24090) );
  NAND2_X1 NAND2_1538( .ZN(II32608), .A1(g18038), .A2(II32607) );
  NAND2_X1 NAND2_1539( .ZN(II32609), .A1(g24090), .A2(II32607) );
  NAND2_X1 NAND2_1540( .ZN(g24887), .A1(II32608), .A2(II32609) );
  NAND2_X1 NAND2_1541( .ZN(II32615), .A1(g18247), .A2(g24091) );
  NAND2_X1 NAND2_1542( .ZN(II32616), .A1(g18247), .A2(II32615) );
  NAND2_X1 NAND2_1543( .ZN(II32617), .A1(g24091), .A2(II32615) );
  NAND2_X1 NAND2_1544( .ZN(g24889), .A1(II32616), .A2(II32617) );
  NAND2_X1 NAND2_1545( .ZN(II32624), .A1(g17927), .A2(g23969) );
  NAND2_X1 NAND2_1546( .ZN(II32625), .A1(g17927), .A2(II32624) );
  NAND2_X1 NAND2_1547( .ZN(II32626), .A1(g23969), .A2(II32624) );
  NAND2_X1 NAND2_1548( .ZN(g24897), .A1(II32625), .A2(II32626) );
  NAND2_X1 NAND2_1549( .ZN(II32633), .A1(g18131), .A2(g23970) );
  NAND2_X2 NAND2_1550( .ZN(II32634), .A1(g18131), .A2(II32633) );
  NAND2_X1 NAND2_1551( .ZN(II32635), .A1(g23970), .A2(II32633) );
  NAND2_X1 NAND2_1552( .ZN(g24900), .A1(II32634), .A2(II32635) );
  NAND2_X1 NAND2_1553( .ZN(II32645), .A1(g18155), .A2(g24093) );
  NAND2_X1 NAND2_1554( .ZN(II32646), .A1(g18155), .A2(II32645) );
  NAND2_X1 NAND2_1555( .ZN(II32647), .A1(g24093), .A2(II32645) );
  NAND2_X1 NAND2_1556( .ZN(g24904), .A1(II32646), .A2(II32647) );
  NAND2_X1 NAND2_1557( .ZN(II32659), .A1(g18038), .A2(g23998) );
  NAND2_X1 NAND2_1558( .ZN(II32660), .A1(g18038), .A2(II32659) );
  NAND2_X1 NAND2_1559( .ZN(II32661), .A1(g23998), .A2(II32659) );
  NAND2_X1 NAND2_1560( .ZN(g24920), .A1(II32660), .A2(II32661) );
  NAND2_X1 NAND2_1561( .ZN(II32668), .A1(g18247), .A2(g23999) );
  NAND2_X1 NAND2_1562( .ZN(II32669), .A1(g18247), .A2(II32668) );
  NAND2_X1 NAND2_1563( .ZN(II32670), .A1(g23999), .A2(II32668) );
  NAND2_X1 NAND2_1564( .ZN(g24923), .A1(II32669), .A2(II32670) );
  NAND2_X1 NAND2_1565( .ZN(II32677), .A1(g23823), .A2(g14165) );
  NAND2_X1 NAND2_1566( .ZN(II32678), .A1(g23823), .A2(II32677) );
  NAND2_X1 NAND2_1567( .ZN(II32679), .A1(g14165), .A2(II32677) );
  NAND2_X1 NAND2_1568( .ZN(g24928), .A1(II32678), .A2(II32679) );
  NAND2_X1 NAND2_1569( .ZN(II32686), .A1(g18155), .A2(g24028) );
  NAND2_X1 NAND2_1570( .ZN(II32687), .A1(g18155), .A2(II32686) );
  NAND2_X1 NAND2_1571( .ZN(II32688), .A1(g24028), .A2(II32686) );
  NAND2_X1 NAND2_1572( .ZN(g24937), .A1(II32687), .A2(II32688) );
  NAND2_X1 NAND2_1573( .ZN(II32695), .A1(g23858), .A2(g14280) );
  NAND2_X1 NAND2_1574( .ZN(II32696), .A1(g23858), .A2(II32695) );
  NAND2_X1 NAND2_1575( .ZN(II32697), .A1(g14280), .A2(II32695) );
  NAND2_X1 NAND2_1576( .ZN(g24940), .A1(II32696), .A2(II32697) );
  NAND2_X1 NAND2_1577( .ZN(II32708), .A1(g23892), .A2(g14402) );
  NAND2_X1 NAND2_1578( .ZN(II32709), .A1(g23892), .A2(II32708) );
  NAND2_X1 NAND2_1579( .ZN(II32710), .A1(g14402), .A2(II32708) );
  NAND2_X1 NAND2_1580( .ZN(g24951), .A1(II32709), .A2(II32710) );
  NAND2_X1 NAND2_1581( .ZN(II32724), .A1(g23913), .A2(g14514) );
  NAND2_X1 NAND2_1582( .ZN(II32725), .A1(g23913), .A2(II32724) );
  NAND2_X1 NAND2_1583( .ZN(II32726), .A1(g14514), .A2(II32724) );
  NAND2_X1 NAND2_1584( .ZN(g24963), .A1(II32725), .A2(II32726) );
  NAND2_X1 NAND2_1585( .ZN(g24975), .A1(g23497), .A2(g74) );
  NAND2_X1 NAND2_1586( .ZN(g24986), .A1(g23513), .A2(g762) );
  NAND2_X1 NAND2_1587( .ZN(g24997), .A1(g23528), .A2(g1448) );
  NAND2_X1 NAND2_1588( .ZN(g25004), .A1(g23644), .A2(g6448) );
  NAND2_X1 NAND2_1589( .ZN(g25005), .A1(g23539), .A2(g2142) );
  NAND2_X1 NAND2_1590( .ZN(g25008), .A1(g23644), .A2(g5438) );
  NAND2_X1 NAND2_1591( .ZN(g25009), .A1(g23644), .A2(g6448) );
  NAND2_X1 NAND2_1592( .ZN(g25010), .A1(g23694), .A2(g6713) );
  NAND2_X1 NAND2_1593( .ZN(g25011), .A1(g23644), .A2(g5438) );
  NAND2_X1 NAND2_1594( .ZN(g25012), .A1(g23644), .A2(g6448) );
  NAND2_X1 NAND2_1595( .ZN(g25013), .A1(g23923), .A2(g6643) );
  NAND2_X1 NAND2_1596( .ZN(g25014), .A1(g23694), .A2(g5473) );
  NAND2_X1 NAND2_1597( .ZN(g25015), .A1(g23694), .A2(g6713) );
  NAND2_X1 NAND2_1598( .ZN(g25016), .A1(g23748), .A2(g7015) );
  NAND2_X1 NAND2_1599( .ZN(g25017), .A1(g23644), .A2(g5438) );
  NAND2_X1 NAND2_1600( .ZN(g25018), .A1(g23644), .A2(g6448) );
  NAND2_X1 NAND2_1601( .ZN(g25019), .A1(g23923), .A2(g6486) );
  NAND2_X1 NAND2_1602( .ZN(g25020), .A1(g23923), .A2(g6643) );
  NAND2_X1 NAND2_1603( .ZN(g25021), .A1(g23694), .A2(g5473) );
  NAND2_X1 NAND2_1604( .ZN(g25022), .A1(g23694), .A2(g6713) );
  NAND2_X1 NAND2_1605( .ZN(g25023), .A1(g23955), .A2(g6945) );
  NAND2_X1 NAND2_1606( .ZN(g25024), .A1(g23748), .A2(g5512) );
  NAND2_X1 NAND2_1607( .ZN(g25025), .A1(g23748), .A2(g7015) );
  NAND2_X2 NAND2_1608( .ZN(g25026), .A1(g23803), .A2(g7265) );
  NAND2_X1 NAND2_1609( .ZN(g25028), .A1(g23644), .A2(g5438) );
  NAND2_X1 NAND2_1610( .ZN(g25029), .A1(g23923), .A2(g6486) );
  NAND2_X1 NAND2_1611( .ZN(g25030), .A1(g23923), .A2(g6643) );
  NAND2_X1 NAND2_1612( .ZN(g25031), .A1(g23694), .A2(g5473) );
  NAND2_X1 NAND2_1613( .ZN(g25032), .A1(g23694), .A2(g6713) );
  NAND2_X1 NAND2_1614( .ZN(g25033), .A1(g23955), .A2(g6751) );
  NAND2_X1 NAND2_1615( .ZN(g25034), .A1(g23955), .A2(g6945) );
  NAND2_X1 NAND2_1616( .ZN(g25035), .A1(g23748), .A2(g5512) );
  NAND2_X1 NAND2_1617( .ZN(g25036), .A1(g23748), .A2(g7015) );
  NAND2_X1 NAND2_1618( .ZN(g25037), .A1(g23984), .A2(g7195) );
  NAND2_X1 NAND2_1619( .ZN(g25038), .A1(g23803), .A2(g5556) );
  NAND2_X1 NAND2_1620( .ZN(g25039), .A1(g23803), .A2(g7265) );
  NAND2_X1 NAND2_1621( .ZN(g25040), .A1(g23923), .A2(g6486) );
  NAND2_X1 NAND2_1622( .ZN(g25041), .A1(g23923), .A2(g6643) );
  NAND2_X1 NAND2_1623( .ZN(g25043), .A1(g23694), .A2(g5473) );
  NAND2_X1 NAND2_1624( .ZN(g25044), .A1(g23955), .A2(g6751) );
  NAND2_X1 NAND2_1625( .ZN(g25045), .A1(g23955), .A2(g6945) );
  NAND2_X1 NAND2_1626( .ZN(g25046), .A1(g23748), .A2(g5512) );
  NAND2_X1 NAND2_1627( .ZN(g25047), .A1(g23748), .A2(g7015) );
  NAND2_X1 NAND2_1628( .ZN(g25048), .A1(g23984), .A2(g7053) );
  NAND2_X1 NAND2_1629( .ZN(g25049), .A1(g23984), .A2(g7195) );
  NAND2_X1 NAND2_1630( .ZN(g25050), .A1(g23803), .A2(g5556) );
  NAND2_X1 NAND2_1631( .ZN(g25051), .A1(g23803), .A2(g7265) );
  NAND2_X1 NAND2_1632( .ZN(g25052), .A1(g24014), .A2(g7391) );
  NAND2_X1 NAND2_1633( .ZN(g25053), .A1(g23923), .A2(g6486) );
  NAND2_X1 NAND2_1634( .ZN(g25054), .A1(g23955), .A2(g6751) );
  NAND2_X1 NAND2_1635( .ZN(g25055), .A1(g23955), .A2(g6945) );
  NAND2_X1 NAND2_1636( .ZN(g25057), .A1(g23748), .A2(g5512) );
  NAND2_X1 NAND2_1637( .ZN(g25058), .A1(g23984), .A2(g7053) );
  NAND2_X1 NAND2_1638( .ZN(g25059), .A1(g23984), .A2(g7195) );
  NAND2_X1 NAND2_1639( .ZN(g25060), .A1(g23803), .A2(g5556) );
  NAND2_X1 NAND2_1640( .ZN(g25061), .A1(g23803), .A2(g7265) );
  NAND2_X1 NAND2_1641( .ZN(g25062), .A1(g24014), .A2(g7303) );
  NAND2_X1 NAND2_1642( .ZN(g25063), .A1(g24014), .A2(g7391) );
  NAND2_X1 NAND2_1643( .ZN(g25064), .A1(g23955), .A2(g6751) );
  NAND2_X1 NAND2_1644( .ZN(g25065), .A1(g23984), .A2(g7053) );
  NAND2_X1 NAND2_1645( .ZN(g25066), .A1(g23984), .A2(g7195) );
  NAND2_X1 NAND2_1646( .ZN(g25068), .A1(g23803), .A2(g5556) );
  NAND2_X1 NAND2_1647( .ZN(g25069), .A1(g24014), .A2(g7303) );
  NAND2_X1 NAND2_1648( .ZN(g25070), .A1(g24014), .A2(g7391) );
  NAND2_X1 NAND2_1649( .ZN(g25071), .A1(g23984), .A2(g7053) );
  NAND2_X1 NAND2_1650( .ZN(g25072), .A1(g24014), .A2(g7303) );
  NAND2_X1 NAND2_1651( .ZN(g25073), .A1(g24014), .A2(g7391) );
  NAND2_X1 NAND2_1652( .ZN(g25074), .A1(g24014), .A2(g7303) );
  NAND2_X1 NAND2_1653( .ZN(g25088), .A1(g23950), .A2(g679) );
  NAND2_X1 NAND2_1654( .ZN(g25096), .A1(g23979), .A2(g1365) );
  NAND2_X1 NAND2_1655( .ZN(g25106), .A1(g24009), .A2(g2059) );
  NAND2_X1 NAND2_1656( .ZN(g25112), .A1(g24043), .A2(g2753) );
  NAND2_X1 NAND2_1657( .ZN(g25200), .A1(g24965), .A2(g3306) );
  NAND2_X1 NAND2_1658( .ZN(g25203), .A1(g24978), .A2(g3462) );
  NAND2_X1 NAND2_1659( .ZN(g25205), .A1(g24989), .A2(g3618) );
  NAND2_X1 NAND2_1660( .ZN(g25210), .A1(g25000), .A2(g3774) );
  NAND4_X1 NAND4_5( .ZN(g25312), .A1(g21211), .A2(g14442), .A3(g10694), .A4(g24590) );
  NAND4_X1 NAND4_6( .ZN(g25320), .A1(g21219), .A2(g14529), .A3(g10714), .A4(g24595) );
  NAND4_X1 NAND4_7( .ZN(g25331), .A1(g21230), .A2(g14584), .A3(g10735), .A4(g24603) );
  NAND4_X1 NAND4_8( .ZN(g25340), .A1(g21235), .A2(g14618), .A3(g10754), .A4(g24610) );
  NAND2_X2 NAND2_1661( .ZN(g25927), .A1(g24965), .A2(g6448) );
  NAND2_X1 NAND2_1662( .ZN(g25928), .A1(g24965), .A2(g5438) );
  NAND2_X1 NAND2_1663( .ZN(g25929), .A1(g24978), .A2(g6713) );
  NAND2_X1 NAND2_1664( .ZN(g25930), .A1(g24978), .A2(g5473) );
  NAND2_X1 NAND2_1665( .ZN(g25931), .A1(g24989), .A2(g7015) );
  NAND2_X1 NAND2_1666( .ZN(g25933), .A1(g24989), .A2(g5512) );
  NAND2_X1 NAND2_1667( .ZN(g25934), .A1(g25000), .A2(g7265) );
  NAND2_X1 NAND2_1668( .ZN(g25936), .A1(g25000), .A2(g5556) );
  NAND2_X1 NAND2_1669( .ZN(g25954), .A1(g22806), .A2(g24517) );
  NAND2_X1 NAND2_1670( .ZN(g25958), .A1(g22847), .A2(g24530) );
  NAND2_X1 NAND2_1671( .ZN(g25964), .A1(g22882), .A2(g24543) );
  NAND2_X1 NAND2_1672( .ZN(g25969), .A1(g22917), .A2(g24555) );
  NAND3_X1 NAND3_76( .ZN(g26059), .A1(g25422), .A2(g25379), .A3(g25274) );
  NAND3_X1 NAND3_77( .ZN(g26066), .A1(g25431), .A2(g25395), .A3(g25283) );
  NAND3_X1 NAND3_78( .ZN(g26073), .A1(g25438), .A2(g25405), .A3(g25291) );
  NAND3_X1 NAND3_79( .ZN(g26079), .A1(g25445), .A2(g25413), .A3(g25301) );
  NAND2_X1 NAND2_1673( .ZN(g26106), .A1(g23644), .A2(g25354) );
  NAND4_X1 NAND4_9( .ZN(g26119), .A1(g8278), .A2(g14657), .A3(g25422), .A4(g25379) );
  NAND2_X1 NAND2_1674( .ZN(g26120), .A1(g23694), .A2(g25369) );
  NAND4_X1 NAND4_10( .ZN(g26129), .A1(g8287), .A2(g14691), .A3(g25431), .A4(g25395) );
  NAND2_X1 NAND2_1675( .ZN(g26130), .A1(g23748), .A2(g25386) );
  NAND4_X1 NAND4_11( .ZN(g26143), .A1(g8296), .A2(g14725), .A3(g25438), .A4(g25405) );
  NAND2_X1 NAND2_1676( .ZN(g26144), .A1(g23803), .A2(g25402) );
  NAND4_X1 NAND4_12( .ZN(g26148), .A1(g8305), .A2(g14753), .A3(g25445), .A4(g25413) );
  NAND2_X1 NAND2_1677( .ZN(g26356), .A1(g16539), .A2(g25183) );
  NAND2_X1 NAND2_1678( .ZN(g26399), .A1(g16571), .A2(g25186) );
  NAND2_X1 NAND2_1679( .ZN(g26440), .A1(g16595), .A2(g25190) );
  NAND2_X1 NAND2_1680( .ZN(g26458), .A1(g25343), .A2(g65) );
  NAND2_X1 NAND2_1681( .ZN(g26472), .A1(g16615), .A2(g25195) );
  NAND2_X1 NAND2_1682( .ZN(g26482), .A1(g25357), .A2(g753) );
  NAND2_X1 NAND2_1683( .ZN(g26498), .A1(g25372), .A2(g1439) );
  NAND2_X1 NAND2_1684( .ZN(g26513), .A1(g25389), .A2(g2133) );
  NAND2_X1 NAND2_1685( .ZN(g26772), .A1(g26320), .A2(g3306) );
  NAND2_X1 NAND2_1686( .ZN(g26779), .A1(g26367), .A2(g3462) );
  NAND2_X1 NAND2_1687( .ZN(g26785), .A1(g26410), .A2(g3618) );
  NAND2_X1 NAND2_1688( .ZN(g26792), .A1(g26451), .A2(g3774) );
  NAND2_X1 NAND2_1689( .ZN(II35020), .A1(g26110), .A2(g26099) );
  NAND2_X1 NAND2_1690( .ZN(II35021), .A1(g26110), .A2(II35020) );
  NAND2_X1 NAND2_1691( .ZN(II35022), .A1(g26099), .A2(II35020) );
  NAND2_X1 NAND2_1692( .ZN(g26859), .A1(II35021), .A2(II35022) );
  NAND2_X1 NAND2_1693( .ZN(II35034), .A1(g26087), .A2(g26154) );
  NAND2_X1 NAND2_1694( .ZN(II35035), .A1(g26087), .A2(II35034) );
  NAND2_X1 NAND2_1695( .ZN(II35036), .A1(g26154), .A2(II35034) );
  NAND2_X1 NAND2_1696( .ZN(g26865), .A1(II35035), .A2(II35036) );
  NAND2_X1 NAND2_1697( .ZN(II35042), .A1(g26151), .A2(g26145) );
  NAND2_X1 NAND2_1698( .ZN(II35043), .A1(g26151), .A2(II35042) );
  NAND2_X1 NAND2_1699( .ZN(II35044), .A1(g26145), .A2(II35042) );
  NAND2_X1 NAND2_1700( .ZN(g26867), .A1(II35043), .A2(II35044) );
  NAND2_X1 NAND2_1701( .ZN(II35057), .A1(g26137), .A2(g26126) );
  NAND2_X1 NAND2_1702( .ZN(II35058), .A1(g26137), .A2(II35057) );
  NAND2_X1 NAND2_1703( .ZN(II35059), .A1(g26126), .A2(II35057) );
  NAND2_X1 NAND2_1704( .ZN(g26874), .A1(II35058), .A2(II35059) );
  NAND4_X1 NAND4_13( .ZN(g26892), .A1(g25699), .A2(g26283), .A3(g25569), .A4(g25631) );
  NAND3_X1 NAND3_80( .ZN(g26902), .A1(g25631), .A2(g26283), .A3(g25569) );
  NAND4_X1 NAND4_14( .ZN(g26906), .A1(g25772), .A2(g26327), .A3(g25648), .A4(g25708) );
  NAND2_X1 NAND2_1705( .ZN(g26911), .A1(g25569), .A2(g26283) );
  NAND3_X1 NAND3_81( .ZN(g26915), .A1(g25708), .A2(g26327), .A3(g25648) );
  NAND4_X1 NAND4_15( .ZN(g26918), .A1(g25826), .A2(g26374), .A3(g25725), .A4(g25781) );
  NAND2_X2 NAND2_1706( .ZN(g26925), .A1(g25648), .A2(g26327) );
  NAND3_X1 NAND3_82( .ZN(g26928), .A1(g25781), .A2(g26374), .A3(g25725) );
  NAND4_X1 NAND4_16( .ZN(g26931), .A1(g25861), .A2(g26417), .A3(g25798), .A4(g25835) );
  NAND2_X1 NAND2_1707( .ZN(II35123), .A1(g26107), .A2(g26096) );
  NAND2_X1 NAND2_1708( .ZN(II35124), .A1(g26107), .A2(II35123) );
  NAND2_X1 NAND2_1709( .ZN(II35125), .A1(g26096), .A2(II35123) );
  NAND2_X1 NAND2_1710( .ZN(g26934), .A1(II35124), .A2(II35125) );
  NAND2_X1 NAND2_1711( .ZN(g26938), .A1(g25725), .A2(g26374) );
  NAND3_X2 NAND3_83( .ZN(g26941), .A1(g25835), .A2(g26417), .A3(g25798) );
  NAND2_X1 NAND2_1712( .ZN(g26947), .A1(g25798), .A2(g26417) );
  NAND2_X1 NAND2_1713( .ZN(g27117), .A1(g26320), .A2(g6448) );
  NAND2_X1 NAND2_1714( .ZN(g27118), .A1(g26320), .A2(g5438) );
  NAND2_X1 NAND2_1715( .ZN(g27119), .A1(g26367), .A2(g6713) );
  NAND2_X1 NAND2_1716( .ZN(g27121), .A1(g26367), .A2(g5473) );
  NAND2_X1 NAND2_1717( .ZN(g27122), .A1(g26410), .A2(g7015) );
  NAND2_X1 NAND2_1718( .ZN(g27124), .A1(g26410), .A2(g5512) );
  NAND2_X1 NAND2_1719( .ZN(g27125), .A1(g26451), .A2(g7265) );
  NAND2_X1 NAND2_1720( .ZN(g27130), .A1(g26451), .A2(g5556) );
  NAND2_X1 NAND2_1721( .ZN(II35701), .A1(g26867), .A2(g26874) );
  NAND2_X1 NAND2_1722( .ZN(II35702), .A1(g26867), .A2(II35701) );
  NAND2_X1 NAND2_1723( .ZN(II35703), .A1(g26874), .A2(II35701) );
  NAND2_X1 NAND2_1724( .ZN(g27379), .A1(II35702), .A2(II35703) );
  NAND2_X1 NAND2_1725( .ZN(II35714), .A1(g26859), .A2(g26865) );
  NAND2_X1 NAND2_1726( .ZN(II35715), .A1(g26859), .A2(II35714) );
  NAND2_X1 NAND2_1727( .ZN(II35716), .A1(g26865), .A2(II35714) );
  NAND2_X1 NAND2_1728( .ZN(g27382), .A1(II35715), .A2(II35716) );
  NAND2_X1 NAND2_1729( .ZN(g27390), .A1(g26989), .A2(g6448) );
  NAND2_X1 NAND2_1730( .ZN(g27395), .A1(g26989), .A2(g5438) );
  NAND2_X1 NAND2_1731( .ZN(g27400), .A1(g27012), .A2(g6713) );
  NAND2_X1 NAND2_1732( .ZN(g27408), .A1(g27012), .A2(g5473) );
  NAND2_X1 NAND2_1733( .ZN(g27413), .A1(g27038), .A2(g7015) );
  NAND2_X1 NAND2_1734( .ZN(g27426), .A1(g27038), .A2(g5512) );
  NAND2_X1 NAND2_1735( .ZN(g27431), .A1(g27066), .A2(g7265) );
  NAND2_X1 NAND2_1736( .ZN(g27447), .A1(g27066), .A2(g5556) );
  NAND2_X1 NAND2_1737( .ZN(II35904), .A1(g27051), .A2(g14831) );
  NAND2_X1 NAND2_1738( .ZN(II35905), .A1(g27051), .A2(II35904) );
  NAND2_X1 NAND2_1739( .ZN(II35906), .A1(g14831), .A2(II35904) );
  NAND2_X1 NAND2_1740( .ZN(g27528), .A1(II35905), .A2(II35906) );
  NAND2_X1 NAND2_1741( .ZN(II35944), .A1(g27078), .A2(g14904) );
  NAND2_X1 NAND2_1742( .ZN(II35945), .A1(g27078), .A2(II35944) );
  NAND2_X1 NAND2_1743( .ZN(II35946), .A1(g14904), .A2(II35944) );
  NAND2_X1 NAND2_1744( .ZN(g27550), .A1(II35945), .A2(II35946) );
  NAND2_X1 NAND2_1745( .ZN(II35974), .A1(g27094), .A2(g14985) );
  NAND2_X1 NAND2_1746( .ZN(II35975), .A1(g27094), .A2(II35974) );
  NAND2_X1 NAND2_1747( .ZN(II35976), .A1(g14985), .A2(II35974) );
  NAND2_X1 NAND2_1748( .ZN(g27566), .A1(II35975), .A2(II35976) );
  NAND2_X1 NAND2_1749( .ZN(g27571), .A1(g26869), .A2(g56) );
  NAND2_X1 NAND2_1750( .ZN(II35992), .A1(g27106), .A2(g15074) );
  NAND2_X1 NAND2_1751( .ZN(II35993), .A1(g27106), .A2(II35992) );
  NAND2_X1 NAND2_1752( .ZN(II35994), .A1(g15074), .A2(II35992) );
  NAND2_X1 NAND2_1753( .ZN(g27576), .A1(II35993), .A2(II35994) );
  NAND2_X1 NAND2_1754( .ZN(g27580), .A1(g26878), .A2(g744) );
  NAND2_X1 NAND2_1755( .ZN(g27583), .A1(g26887), .A2(g1430) );
  NAND2_X1 NAND2_1756( .ZN(g27587), .A1(g26897), .A2(g2124) );
  NAND2_X1 NAND2_1757( .ZN(g27626), .A1(g26989), .A2(g3306) );
  NAND2_X1 NAND2_1758( .ZN(g27627), .A1(g27012), .A2(g3462) );
  NAND2_X1 NAND2_1759( .ZN(g27628), .A1(g27038), .A2(g3618) );
  NAND2_X1 NAND2_1760( .ZN(g27630), .A1(g27066), .A2(g3774) );
  NAND2_X1 NAND2_1761( .ZN(g27738), .A1(g25367), .A2(g27415) );
  NAND2_X2 NAND2_1762( .ZN(g27743), .A1(g25384), .A2(g27436) );
  NAND2_X1 NAND2_1763( .ZN(g27751), .A1(g25400), .A2(g27455) );
  NAND2_X1 NAND2_1764( .ZN(g27756), .A1(g25410), .A2(g27471) );
  NAND2_X1 NAND2_1765( .ZN(II36256), .A1(g27527), .A2(g15859) );
  NAND2_X1 NAND2_1766( .ZN(II36257), .A1(g27527), .A2(II36256) );
  NAND2_X1 NAND2_1767( .ZN(II36258), .A1(g15859), .A2(II36256) );
  NAND2_X1 NAND2_1768( .ZN(g27801), .A1(II36257), .A2(II36258) );
  NAND2_X1 NAND2_1769( .ZN(II36270), .A1(g27549), .A2(g15890) );
  NAND2_X1 NAND2_1770( .ZN(II36271), .A1(g27549), .A2(II36270) );
  NAND2_X1 NAND2_1771( .ZN(II36272), .A1(g15890), .A2(II36270) );
  NAND2_X1 NAND2_1772( .ZN(g27809), .A1(II36271), .A2(II36272) );
  NAND2_X1 NAND2_1773( .ZN(II36289), .A1(g27565), .A2(g15923) );
  NAND2_X1 NAND2_1774( .ZN(II36290), .A1(g27565), .A2(II36289) );
  NAND2_X1 NAND2_1775( .ZN(II36291), .A1(g15923), .A2(II36289) );
  NAND2_X1 NAND2_1776( .ZN(g27830), .A1(II36290), .A2(II36291) );
  NAND2_X1 NAND2_1777( .ZN(II36300), .A1(g27382), .A2(g27379) );
  NAND2_X1 NAND2_1778( .ZN(II36301), .A1(g27382), .A2(II36300) );
  NAND2_X1 NAND2_1779( .ZN(II36302), .A1(g27379), .A2(II36300) );
  NAND2_X1 NAND2_1780( .ZN(g27838), .A1(II36301), .A2(II36302) );
  NAND2_X1 NAND2_1781( .ZN(II36314), .A1(g27575), .A2(g15952) );
  NAND2_X1 NAND2_1782( .ZN(II36315), .A1(g27575), .A2(II36314) );
  NAND2_X1 NAND2_1783( .ZN(II36316), .A1(g15952), .A2(II36314) );
  NAND2_X1 NAND2_1784( .ZN(g27846), .A1(II36315), .A2(II36316) );
  NAND2_X1 NAND2_1785( .ZN(II36591), .A1(g27529), .A2(g14885) );
  NAND2_X1 NAND2_1786( .ZN(II36592), .A1(g27529), .A2(II36591) );
  NAND2_X1 NAND2_1787( .ZN(II36593), .A1(g14885), .A2(II36591) );
  NAND2_X1 NAND2_1788( .ZN(g28046), .A1(II36592), .A2(II36593) );
  NAND2_X1 NAND2_1789( .ZN(II36666), .A1(g27551), .A2(g14966) );
  NAND2_X1 NAND2_1790( .ZN(II36667), .A1(g27551), .A2(II36666) );
  NAND2_X1 NAND2_1791( .ZN(II36668), .A1(g14966), .A2(II36666) );
  NAND2_X1 NAND2_1792( .ZN(g28075), .A1(II36667), .A2(II36668) );
  NAND2_X1 NAND2_1793( .ZN(II36731), .A1(g27567), .A2(g15055) );
  NAND2_X1 NAND2_1794( .ZN(II36732), .A1(g27567), .A2(II36731) );
  NAND2_X1 NAND2_1795( .ZN(II36733), .A1(g15055), .A2(II36731) );
  NAND2_X1 NAND2_1796( .ZN(g28100), .A1(II36732), .A2(II36733) );
  NAND2_X1 NAND2_1797( .ZN(II36779), .A1(g27577), .A2(g15151) );
  NAND2_X1 NAND2_1798( .ZN(II36780), .A1(g27577), .A2(II36779) );
  NAND2_X1 NAND2_1799( .ZN(II36781), .A1(g15151), .A2(II36779) );
  NAND2_X1 NAND2_1800( .ZN(g28118), .A1(II36780), .A2(II36781) );
  NAND2_X1 NAND2_1801( .ZN(II37295), .A1(g27827), .A2(g27814) );
  NAND2_X1 NAND2_1802( .ZN(II37296), .A1(g27827), .A2(II37295) );
  NAND2_X1 NAND2_1803( .ZN(II37297), .A1(g27814), .A2(II37295) );
  NAND2_X1 NAND2_1804( .ZN(g28384), .A1(II37296), .A2(II37297) );
  NAND2_X1 NAND2_1805( .ZN(II37303), .A1(g27802), .A2(g27900) );
  NAND2_X1 NAND2_1806( .ZN(II37304), .A1(g27802), .A2(II37303) );
  NAND2_X1 NAND2_1807( .ZN(II37305), .A1(g27900), .A2(II37303) );
  NAND2_X1 NAND2_1808( .ZN(g28386), .A1(II37304), .A2(II37305) );
  NAND2_X1 NAND2_1809( .ZN(II37311), .A1(g27897), .A2(g27883) );
  NAND2_X1 NAND2_1810( .ZN(II37312), .A1(g27897), .A2(II37311) );
  NAND2_X1 NAND2_1811( .ZN(II37313), .A1(g27883), .A2(II37311) );
  NAND2_X1 NAND2_1812( .ZN(g28388), .A1(II37312), .A2(II37313) );
  NAND2_X1 NAND2_1813( .ZN(II37322), .A1(g27865), .A2(g27855) );
  NAND2_X1 NAND2_1814( .ZN(II37323), .A1(g27865), .A2(II37322) );
  NAND2_X1 NAND2_1815( .ZN(II37324), .A1(g27855), .A2(II37322) );
  NAND2_X1 NAND2_1816( .ZN(g28391), .A1(II37323), .A2(II37324) );
  NAND2_X2 NAND2_1817( .ZN(II37356), .A1(g27824), .A2(g27811) );
  NAND2_X1 NAND2_1818( .ZN(II37357), .A1(g27824), .A2(II37356) );
  NAND2_X1 NAND2_1819( .ZN(II37358), .A1(g27811), .A2(II37356) );
  NAND2_X1 NAND2_1820( .ZN(g28415), .A1(II37357), .A2(II37358) );
  NAND2_X1 NAND2_1821( .ZN(II37813), .A1(g28388), .A2(g28391) );
  NAND2_X1 NAND2_1822( .ZN(II37814), .A1(g28388), .A2(II37813) );
  NAND2_X1 NAND2_1823( .ZN(II37815), .A1(g28391), .A2(II37813) );
  NAND2_X1 NAND2_1824( .ZN(g28842), .A1(II37814), .A2(II37815) );
  NAND2_X1 NAND2_1825( .ZN(II37822), .A1(g28384), .A2(g28386) );
  NAND2_X1 NAND2_1826( .ZN(II37823), .A1(g28384), .A2(II37822) );
  NAND2_X1 NAND2_1827( .ZN(II37824), .A1(g28386), .A2(II37822) );
  NAND2_X1 NAND2_1828( .ZN(g28845), .A1(II37823), .A2(II37824) );
  NAND2_X1 NAND2_1829( .ZN(g28978), .A1(g9150), .A2(g28512) );
  NAND2_X1 NAND2_1830( .ZN(g29001), .A1(g9161), .A2(g28512) );
  NAND2_X1 NAND2_1831( .ZN(g29008), .A1(g9174), .A2(g28540) );
  NAND2_X1 NAND2_1832( .ZN(g29026), .A1(g9187), .A2(g28512) );
  NAND2_X1 NAND2_1833( .ZN(g29030), .A1(g9203), .A2(g28540) );
  NAND2_X1 NAND2_1834( .ZN(g29038), .A1(g9216), .A2(g28567) );
  NAND2_X1 NAND2_1835( .ZN(g29045), .A1(g9232), .A2(g28512) );
  NAND2_X1 NAND2_1836( .ZN(g29049), .A1(g9248), .A2(g28540) );
  NAND2_X1 NAND2_1837( .ZN(g29053), .A1(g9264), .A2(g28567) );
  NAND2_X1 NAND2_1838( .ZN(g29060), .A1(g9277), .A2(g28595) );
  NAND2_X1 NAND2_1839( .ZN(g29062), .A1(g9310), .A2(g28540) );
  NAND2_X1 NAND2_1840( .ZN(g29068), .A1(g9326), .A2(g28567) );
  NAND2_X1 NAND2_1841( .ZN(g29072), .A1(g9342), .A2(g28595) );
  NAND2_X1 NAND2_1842( .ZN(g29076), .A1(g9391), .A2(g28567) );
  NAND2_X1 NAND2_1843( .ZN(g29080), .A1(g9407), .A2(g28595) );
  NAND2_X1 NAND2_1844( .ZN(g29087), .A1(g9488), .A2(g28595) );
  NAND2_X1 NAND2_1845( .ZN(g29088), .A1(g9507), .A2(g28512) );
  NAND2_X1 NAND2_1846( .ZN(g29096), .A1(g9649), .A2(g28540) );
  NAND2_X1 NAND2_1847( .ZN(g29103), .A1(g9795), .A2(g28567) );
  NAND2_X1 NAND2_1848( .ZN(g29107), .A1(g9941), .A2(g28595) );
  NAND2_X1 NAND2_1849( .ZN(II38378), .A1(g28845), .A2(g28842) );
  NAND2_X1 NAND2_1850( .ZN(II38379), .A1(g28845), .A2(II38378) );
  NAND2_X1 NAND2_1851( .ZN(II38380), .A1(g28842), .A2(II38378) );
  NAND2_X1 NAND2_1852( .ZN(g29265), .A1(II38379), .A2(II38380) );
  NAND2_X1 NAND2_1853( .ZN(II38810), .A1(g29303), .A2(g15904) );
  NAND2_X1 NAND2_1854( .ZN(II38811), .A1(g29303), .A2(II38810) );
  NAND2_X1 NAND2_1855( .ZN(II38812), .A1(g15904), .A2(II38810) );
  NAND2_X1 NAND2_1856( .ZN(g29498), .A1(II38811), .A2(II38812) );
  NAND2_X1 NAND2_1857( .ZN(II38820), .A1(g29313), .A2(g15933) );
  NAND2_X1 NAND2_1858( .ZN(II38821), .A1(g29313), .A2(II38820) );
  NAND2_X1 NAND2_1859( .ZN(II38822), .A1(g15933), .A2(II38820) );
  NAND2_X1 NAND2_1860( .ZN(g29500), .A1(II38821), .A2(II38822) );
  NAND2_X1 NAND2_1861( .ZN(II38831), .A1(g29324), .A2(g15962) );
  NAND2_X1 NAND2_1862( .ZN(II38832), .A1(g29324), .A2(II38831) );
  NAND2_X1 NAND2_1863( .ZN(II38833), .A1(g15962), .A2(II38831) );
  NAND2_X1 NAND2_1864( .ZN(g29503), .A1(II38832), .A2(II38833) );
  NAND2_X1 NAND2_1865( .ZN(II38841), .A1(g29333), .A2(g15981) );
  NAND2_X1 NAND2_1866( .ZN(II38842), .A1(g29333), .A2(II38841) );
  NAND2_X1 NAND2_1867( .ZN(II38843), .A1(g15981), .A2(II38841) );
  NAND2_X1 NAND2_1868( .ZN(g29505), .A1(II38842), .A2(II38843) );
  NAND2_X1 NAND2_1869( .ZN(II39323), .A1(g29721), .A2(g29713) );
  NAND2_X1 NAND2_1870( .ZN(II39324), .A1(g29721), .A2(II39323) );
  NAND2_X1 NAND2_1871( .ZN(II39325), .A1(g29713), .A2(II39323) );
  NAND2_X1 NAND2_1872( .ZN(g29911), .A1(II39324), .A2(II39325) );
  NAND2_X1 NAND2_1873( .ZN(II39331), .A1(g29705), .A2(g29751) );
  NAND2_X1 NAND2_1874( .ZN(II39332), .A1(g29705), .A2(II39331) );
  NAND2_X1 NAND2_1875( .ZN(II39333), .A1(g29751), .A2(II39331) );
  NAND2_X2 NAND2_1876( .ZN(g29913), .A1(II39332), .A2(II39333) );
  NAND2_X2 NAND2_1877( .ZN(II39339), .A1(g29748), .A2(g29741) );
  NAND2_X2 NAND2_1878( .ZN(II39340), .A1(g29748), .A2(II39339) );
  NAND2_X1 NAND2_1879( .ZN(II39341), .A1(g29741), .A2(II39339) );
  NAND2_X1 NAND2_1880( .ZN(g29915), .A1(II39340), .A2(II39341) );
  NAND2_X1 NAND2_1881( .ZN(II39347), .A1(g29732), .A2(g29728) );
  NAND2_X1 NAND2_1882( .ZN(II39348), .A1(g29732), .A2(II39347) );
  NAND2_X1 NAND2_1883( .ZN(II39349), .A1(g29728), .A2(II39347) );
  NAND2_X1 NAND2_1884( .ZN(g29917), .A1(II39348), .A2(II39349) );
  NAND2_X1 NAND2_1885( .ZN(II39359), .A1(g29766), .A2(g15880) );
  NAND2_X1 NAND2_1886( .ZN(II39360), .A1(g29766), .A2(II39359) );
  NAND2_X1 NAND2_1887( .ZN(II39361), .A1(g15880), .A2(II39359) );
  NAND2_X1 NAND2_1888( .ZN(g29923), .A1(II39360), .A2(II39361) );
  NAND2_X1 NAND2_1889( .ZN(II39367), .A1(g29767), .A2(g15913) );
  NAND2_X1 NAND2_1890( .ZN(II39368), .A1(g29767), .A2(II39367) );
  NAND2_X1 NAND2_1891( .ZN(II39369), .A1(g15913), .A2(II39367) );
  NAND2_X1 NAND2_1892( .ZN(g29925), .A1(II39368), .A2(II39369) );
  NAND2_X1 NAND2_1893( .ZN(II39375), .A1(g29768), .A2(g15942) );
  NAND2_X1 NAND2_1894( .ZN(II39376), .A1(g29768), .A2(II39375) );
  NAND2_X1 NAND2_1895( .ZN(II39377), .A1(g15942), .A2(II39375) );
  NAND2_X1 NAND2_1896( .ZN(g29927), .A1(II39376), .A2(II39377) );
  NAND2_X1 NAND2_1897( .ZN(II39384), .A1(g29718), .A2(g29710) );
  NAND2_X1 NAND2_1898( .ZN(II39385), .A1(g29718), .A2(II39384) );
  NAND2_X1 NAND2_1899( .ZN(II39386), .A1(g29710), .A2(II39384) );
  NAND2_X1 NAND2_1900( .ZN(g29930), .A1(II39385), .A2(II39386) );
  NAND2_X1 NAND2_1901( .ZN(II39391), .A1(g29769), .A2(g15971) );
  NAND2_X1 NAND2_1902( .ZN(II39392), .A1(g29769), .A2(II39391) );
  NAND2_X1 NAND2_1903( .ZN(II39393), .A1(g15971), .A2(II39391) );
  NAND2_X1 NAND2_1904( .ZN(g29931), .A1(II39392), .A2(II39393) );
  NAND2_X1 NAND2_1905( .ZN(II39532), .A1(g29915), .A2(g29917) );
  NAND2_X1 NAND2_1906( .ZN(II39533), .A1(g29915), .A2(II39532) );
  NAND2_X1 NAND2_1907( .ZN(II39534), .A1(g29917), .A2(II39532) );
  NAND2_X1 NAND2_1908( .ZN(g30034), .A1(II39533), .A2(II39534) );
  NAND2_X1 NAND2_1909( .ZN(II39539), .A1(g29911), .A2(g29913) );
  NAND2_X1 NAND2_1910( .ZN(II39540), .A1(g29911), .A2(II39539) );
  NAND2_X1 NAND2_1911( .ZN(II39541), .A1(g29913), .A2(II39539) );
  NAND2_X1 NAND2_1912( .ZN(g30035), .A1(II39540), .A2(II39541) );
  NAND2_X1 NAND2_1913( .ZN(II39689), .A1(g30035), .A2(g30034) );
  NAND2_X1 NAND2_1914( .ZN(II39690), .A1(g30035), .A2(II39689) );
  NAND2_X1 NAND2_1915( .ZN(II39691), .A1(g30034), .A2(II39689) );
  NAND2_X1 NAND2_1916( .ZN(g30228), .A1(II39690), .A2(II39691) );
  NAND2_X1 NAND2_1917( .ZN(II40558), .A1(g30605), .A2(g30597) );
  NAND2_X1 NAND2_1918( .ZN(II40559), .A1(g30605), .A2(II40558) );
  NAND2_X1 NAND2_1919( .ZN(II40560), .A1(g30597), .A2(II40558) );
  NAND2_X1 NAND2_1920( .ZN(g30768), .A1(II40559), .A2(II40560) );
  NAND2_X1 NAND2_1921( .ZN(II40571), .A1(g30588), .A2(g30632) );
  NAND2_X1 NAND2_1922( .ZN(II40572), .A1(g30588), .A2(II40571) );
  NAND2_X1 NAND2_1923( .ZN(II40573), .A1(g30632), .A2(II40571) );
  NAND2_X1 NAND2_1924( .ZN(g30771), .A1(II40572), .A2(II40573) );
  NAND2_X1 NAND2_1925( .ZN(II40587), .A1(g30629), .A2(g30622) );
  NAND2_X1 NAND2_1926( .ZN(II40588), .A1(g30629), .A2(II40587) );
  NAND2_X1 NAND2_1927( .ZN(II40589), .A1(g30622), .A2(II40587) );
  NAND2_X1 NAND2_1928( .ZN(g30775), .A1(II40588), .A2(II40589) );
  NAND2_X1 NAND2_1929( .ZN(II40603), .A1(g30614), .A2(g30610) );
  NAND2_X1 NAND2_1930( .ZN(II40604), .A1(g30614), .A2(II40603) );
  NAND2_X1 NAND2_1931( .ZN(II40605), .A1(g30610), .A2(II40603) );
  NAND2_X2 NAND2_1932( .ZN(g30779), .A1(II40604), .A2(II40605) );
  NAND2_X1 NAND2_1933( .ZN(II40627), .A1(g30602), .A2(g30594) );
  NAND2_X1 NAND2_1934( .ZN(II40628), .A1(g30602), .A2(II40627) );
  NAND2_X1 NAND2_1935( .ZN(II40629), .A1(g30594), .A2(II40627) );
  NAND2_X1 NAND2_1936( .ZN(g30791), .A1(II40628), .A2(II40629) );
  NAND2_X1 NAND2_1937( .ZN(II41010), .A1(g30775), .A2(g30779) );
  NAND2_X1 NAND2_1938( .ZN(II41011), .A1(g30775), .A2(II41010) );
  NAND2_X1 NAND2_1939( .ZN(II41012), .A1(g30779), .A2(II41010) );
  NAND2_X1 NAND2_1940( .ZN(g30926), .A1(II41011), .A2(II41012) );
  NAND2_X1 NAND2_1941( .ZN(II41017), .A1(g30768), .A2(g30771) );
  NAND2_X1 NAND2_1942( .ZN(II41018), .A1(g30768), .A2(II41017) );
  NAND2_X1 NAND2_1943( .ZN(II41019), .A1(g30771), .A2(II41017) );
  NAND2_X1 NAND2_1944( .ZN(g30927), .A1(II41018), .A2(II41019) );
  NAND2_X1 NAND2_1945( .ZN(II41064), .A1(g30927), .A2(g30926) );
  NAND2_X1 NAND2_1946( .ZN(II41065), .A1(g30927), .A2(II41064) );
  NAND2_X1 NAND2_1947( .ZN(II41066), .A1(g30926), .A2(II41064) );
  NAND2_X1 NAND2_1948( .ZN(g30952), .A1(II41065), .A2(II41066) );
  NOR3_X1 NOR3_0( .ZN(g7528), .A1(g3151), .A2(g3142), .A3(g3147) );
  NOR2_X1 NOR2_0( .ZN(g7575), .A1(g2984), .A2(g2985) );
  NOR2_X1 NOR2_1( .ZN(g7795), .A1(g2992), .A2(g2991) );
  NOR3_X1 NOR4_0_A( .ZN(extra0), .A1(g3198), .A2(g8120), .A3(g3194) );
  NOR2_X1 NOR4_0( .ZN(g8430), .A1(extra0), .A2(g3191) );
  NOR3_X1 NOR3_1( .ZN(g10784), .A1(g5630), .A2(g5649), .A3(g5676) );
  NOR3_X1 NOR3_2( .ZN(g10789), .A1(g5650), .A2(g5677), .A3(g5709) );
  NOR3_X1 NOR3_3( .ZN(g10793), .A1(g5658), .A2(g5687), .A3(g5728) );
  NOR3_X1 NOR3_4( .ZN(g10797), .A1(g5678), .A2(g5710), .A3(g5757) );
  NOR3_X1 NOR3_5( .ZN(g10801), .A1(g5688), .A2(g5729), .A3(g5767) );
  NOR3_X1 NOR3_6( .ZN(g10805), .A1(g5696), .A2(g5739), .A3(g5786) );
  NOR3_X1 NOR3_7( .ZN(g10810), .A1(g5711), .A2(g5758), .A3(g5807) );
  NOR3_X1 NOR3_8( .ZN(g10814), .A1(g5730), .A2(g5768), .A3(g5816) );
  NOR3_X2 NOR3_9( .ZN(g10818), .A1(g5740), .A2(g5787), .A3(g5826) );
  NOR3_X2 NOR3_10( .ZN(g10822), .A1(g5748), .A2(g5797), .A3(g5845) );
  NOR3_X2 NOR3_11( .ZN(g10831), .A1(g5769), .A2(g5817), .A3(g5863) );
  NOR3_X2 NOR3_12( .ZN(g10835), .A1(g5788), .A2(g5827), .A3(g5872) );
  NOR3_X1 NOR3_13( .ZN(g10839), .A1(g5798), .A2(g5846), .A3(g5882) );
  NOR3_X1 NOR3_14( .ZN(g10851), .A1(g5828), .A2(g5873), .A3(g5910) );
  NOR3_X1 NOR3_15( .ZN(g10855), .A1(g5847), .A2(g5883), .A3(g5919) );
  NOR3_X1 NOR3_16( .ZN(g10872), .A1(g5884), .A2(g5920), .A3(g5949) );
  NOR3_X1 NOR3_17( .ZN(g11600), .A1(g9049), .A2(g9064), .A3(g9078) );
  NOR3_X1 NOR4_1_A( .ZN(extra1), .A1(g8183), .A2(g11332), .A3(g7928) );
  NOR2_X1 NOR4_1( .ZN(g11622), .A1(extra1), .A2(g11069) );
  NOR3_X1 NOR3_18( .ZN(g11624), .A1(g9062), .A2(g9075), .A3(g9091) );
  NOR3_X1 NOR3_19( .ZN(g11627), .A1(g9063), .A2(g9077), .A3(g9093) );
  NOR3_X1 NOR3_20( .ZN(g11630), .A1(g9066), .A2(g9081), .A3(g9097) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(g11481), .A2(g8045), .A3(g7928) );
  NOR2_X1 NOR4_2( .ZN(g11643), .A1(extra2), .A2(g11069) );
  NOR3_X1 NOR3_21( .ZN(g11644), .A1(g9076), .A2(g9092), .A3(g9102) );
  NOR3_X1 NOR3_22( .ZN(g11647), .A1(g9079), .A2(g9094), .A3(g9103) );
  NOR3_X1 NOR3_23( .ZN(g11650), .A1(g9080), .A2(g9096), .A3(g9105) );
  NOR3_X1 NOR3_24( .ZN(g11653), .A1(g9083), .A2(g9100), .A3(g9109) );
  NOR3_X1 NOR4_3_A( .ZN(extra3), .A1(g8183), .A2(g8045), .A3(g7928) );
  NOR2_X1 NOR4_3( .ZN(g11660), .A1(extra3), .A2(g11069) );
  NOR3_X1 NOR3_25( .ZN(g11663), .A1(g9095), .A2(g9104), .A3(g9112) );
  NOR3_X1 NOR3_26( .ZN(g11666), .A1(g9098), .A2(g9106), .A3(g9113) );
  NOR3_X1 NOR3_27( .ZN(g11669), .A1(g9099), .A2(g9108), .A3(g9115) );
  NOR3_X1 NOR3_28( .ZN(g11675), .A1(g9107), .A2(g9114), .A3(g9120) );
  NOR3_X1 NOR3_29( .ZN(g11678), .A1(g9110), .A2(g9116), .A3(g9121) );
  NOR3_X1 NOR3_30( .ZN(g11681), .A1(g9111), .A2(g9118), .A3(g9123) );
  NOR3_X1 NOR3_31( .ZN(g11687), .A1(g9117), .A2(g9122), .A3(g9126) );
  NOR3_X1 NOR3_32( .ZN(g11690), .A1(g9119), .A2(g9124), .A3(g9127) );
  NOR3_X1 NOR3_33( .ZN(g11697), .A1(g9125), .A2(g9131), .A3(g9133) );
  NOR3_X1 NOR3_34( .ZN(g11703), .A1(g9132), .A2(g9137), .A3(g9139) );
  NOR3_X1 NOR3_35( .ZN(g11711), .A1(g9138), .A2(g9143), .A3(g9145) );
  NOR3_X1 NOR3_36( .ZN(g11744), .A1(g9241), .A2(g9301), .A3(g9364) );
  NOR3_X1 NOR3_37( .ZN(g11759), .A1(g9302), .A2(g9365), .A3(g9438) );
  NOR3_X1 NOR3_38( .ZN(g11760), .A1(g9319), .A2(g9382), .A3(g9461) );
  NOR3_X1 NOR3_39( .ZN(g11767), .A1(g9366), .A2(g9439), .A3(g9518) );
  NOR3_X1 NOR3_40( .ZN(g11768), .A1(g9367), .A2(g9441), .A3(g9521) );
  NOR3_X1 NOR3_41( .ZN(g11772), .A1(g9383), .A2(g9462), .A3(g9580) );
  NOR3_X1 NOR3_42( .ZN(g11773), .A1(g9400), .A2(g9479), .A3(g9603) );
  NOR3_X1 NOR3_43( .ZN(g11780), .A1(g9440), .A2(g9519), .A3(g9630) );
  NOR3_X1 NOR3_44( .ZN(g11781), .A1(g9442), .A2(g9522), .A3(g9633) );
  NOR3_X1 NOR3_45( .ZN(g11784), .A1(g9463), .A2(g9581), .A3(g9660) );
  NOR3_X1 NOR3_46( .ZN(g11785), .A1(g9464), .A2(g9583), .A3(g9663) );
  NOR3_X1 NOR3_47( .ZN(g11789), .A1(g9480), .A2(g9604), .A3(g9722) );
  NOR3_X1 NOR3_48( .ZN(g11790), .A1(g9497), .A2(g9621), .A3(g9745) );
  NOR3_X1 NOR3_49( .ZN(g11799), .A1(g9520), .A2(g9631), .A3(g9759) );
  NOR3_X1 NOR3_50( .ZN(g11800), .A1(g9523), .A2(g9634), .A3(g9762) );
  NOR3_X1 NOR3_51( .ZN(g11806), .A1(g9582), .A2(g9661), .A3(g9776) );
  NOR3_X1 NOR3_52( .ZN(g11807), .A1(g9584), .A2(g9664), .A3(g9779) );
  NOR3_X1 NOR3_53( .ZN(g11810), .A1(g9605), .A2(g9723), .A3(g9806) );
  NOR3_X1 NOR3_54( .ZN(g11811), .A1(g9606), .A2(g9725), .A3(g9809) );
  NOR3_X1 NOR3_55( .ZN(g11815), .A1(g9622), .A2(g9746), .A3(g9868) );
  NOR3_X1 NOR3_56( .ZN(g11822), .A1(g9632), .A2(g9760), .A3(g9888) );
  NOR3_X1 NOR3_57( .ZN(g11823), .A1(g9635), .A2(g9763), .A3(g9891) );
  NOR3_X1 NOR3_58( .ZN(g11828), .A1(g9639), .A2(g9764), .A3(g9892) );
  NOR3_X1 NOR3_59( .ZN(g11830), .A1(g9647), .A2(g9773), .A3(g9901) );
  NOR3_X1 NOR3_60( .ZN(g11831), .A1(g9648), .A2(g9775), .A3(g9904) );
  NOR3_X1 NOR3_61( .ZN(g11832), .A1(g9662), .A2(g9777), .A3(g9905) );
  NOR3_X1 NOR3_62( .ZN(g11833), .A1(g9665), .A2(g9780), .A3(g9908) );
  NOR3_X1 NOR3_63( .ZN(g11839), .A1(g9724), .A2(g9807), .A3(g9922) );
  NOR3_X1 NOR3_64( .ZN(g11840), .A1(g9726), .A2(g9810), .A3(g9925) );
  NOR3_X1 NOR3_65( .ZN(g11843), .A1(g9747), .A2(g9869), .A3(g9952) );
  NOR3_X1 NOR3_66( .ZN(g11844), .A1(g9748), .A2(g9871), .A3(g9955) );
  NOR3_X1 NOR3_67( .ZN(g11855), .A1(g9761), .A2(g9889), .A3(g10009) );
  NOR3_X1 NOR3_68( .ZN(g11860), .A1(g9765), .A2(g9893), .A3(g10012) );
  NOR3_X1 NOR3_69( .ZN(g11861), .A1(g9766), .A2(g9894), .A3(g10013) );
  NOR3_X1 NOR3_70( .ZN(g11863), .A1(g9774), .A2(g9902), .A3(g10035) );
  NOR3_X1 NOR3_71( .ZN(g11864), .A1(g9778), .A2(g9906), .A3(g10042) );
  NOR3_X1 NOR3_72( .ZN(g11865), .A1(g9781), .A2(g9909), .A3(g10045) );
  NOR3_X1 NOR3_73( .ZN(g11870), .A1(g9785), .A2(g9910), .A3(g10046) );
  NOR3_X1 NOR3_74( .ZN(g11872), .A1(g9793), .A2(g9919), .A3(g10055) );
  NOR3_X1 NOR3_75( .ZN(g11873), .A1(g9794), .A2(g9921), .A3(g10058) );
  NOR3_X1 NOR3_76( .ZN(g11874), .A1(g9808), .A2(g9923), .A3(g10059) );
  NOR3_X1 NOR3_77( .ZN(g11875), .A1(g9811), .A2(g9926), .A3(g10062) );
  NOR3_X2 NOR3_78( .ZN(g11881), .A1(g9870), .A2(g9953), .A3(g10076) );
  NOR3_X2 NOR3_79( .ZN(g11882), .A1(g9872), .A2(g9956), .A3(g10079) );
  NOR3_X1 NOR3_80( .ZN(g11889), .A1(g9887), .A2(g10007), .A3(g10101) );
  NOR3_X1 NOR3_81( .ZN(g11890), .A1(g9890), .A2(g10010), .A3(g10103) );
  NOR3_X1 NOR3_82( .ZN(g11896), .A1(g9903), .A2(g10036), .A3(g10112) );
  NOR3_X1 NOR3_83( .ZN(g11897), .A1(g9907), .A2(g10043), .A3(g10118) );
  NOR3_X1 NOR3_84( .ZN(g11902), .A1(g9911), .A2(g10047), .A3(g10121) );
  NOR3_X1 NOR3_85( .ZN(g11903), .A1(g9912), .A2(g10048), .A3(g10122) );
  NOR3_X1 NOR3_86( .ZN(g11905), .A1(g9920), .A2(g10056), .A3(g10144) );
  NOR3_X1 NOR3_87( .ZN(g11906), .A1(g9924), .A2(g10060), .A3(g10151) );
  NOR3_X1 NOR3_88( .ZN(g11907), .A1(g9927), .A2(g10063), .A3(g10154) );
  NOR3_X1 NOR3_89( .ZN(g11912), .A1(g9931), .A2(g10064), .A3(g10155) );
  NOR3_X1 NOR3_90( .ZN(g11914), .A1(g9939), .A2(g10073), .A3(g10164) );
  NOR3_X1 NOR3_91( .ZN(g11915), .A1(g9940), .A2(g10075), .A3(g10167) );
  NOR3_X1 NOR3_92( .ZN(g11916), .A1(g9954), .A2(g10077), .A3(g10168) );
  NOR3_X1 NOR3_93( .ZN(g11917), .A1(g9957), .A2(g10080), .A3(g10171) );
  NOR3_X1 NOR3_94( .ZN(g11928), .A1(g10008), .A2(g10102), .A3(g10192) );
  NOR3_X1 NOR3_95( .ZN(g11934), .A1(g10011), .A2(g10104), .A3(g10193) );
  NOR3_X1 NOR3_96( .ZN(g11935), .A1(g10014), .A2(g10106), .A3(g10196) );
  NOR3_X1 NOR3_97( .ZN(g11938), .A1(g10037), .A2(g10113), .A3(g10201) );
  NOR3_X1 NOR3_98( .ZN(g11939), .A1(g10041), .A2(g10116), .A3(g10206) );
  NOR3_X1 NOR3_99( .ZN(g11940), .A1(g10044), .A2(g10119), .A3(g10208) );
  NOR3_X1 NOR3_100( .ZN(g11946), .A1(g10057), .A2(g10145), .A3(g10217) );
  NOR3_X1 NOR3_101( .ZN(g11947), .A1(g10061), .A2(g10152), .A3(g10223) );
  NOR3_X1 NOR3_102( .ZN(g11952), .A1(g10065), .A2(g10156), .A3(g10226) );
  NOR3_X1 NOR3_103( .ZN(g11953), .A1(g10066), .A2(g10157), .A3(g10227) );
  NOR3_X1 NOR3_104( .ZN(g11955), .A1(g10074), .A2(g10165), .A3(g10249) );
  NOR3_X1 NOR3_105( .ZN(g11956), .A1(g10078), .A2(g10169), .A3(g10256) );
  NOR3_X1 NOR3_106( .ZN(g11957), .A1(g10081), .A2(g10172), .A3(g10259) );
  NOR3_X1 NOR3_107( .ZN(g11962), .A1(g10085), .A2(g10173), .A3(g10260) );
  NOR3_X1 NOR3_108( .ZN(g11964), .A1(g10093), .A2(g10182), .A3(g10269) );
  NOR3_X1 NOR3_109( .ZN(g11965), .A1(g10094), .A2(g10184), .A3(g10272) );
  NOR3_X1 NOR3_110( .ZN(g11974), .A1(g10105), .A2(g10194), .A3(g10279) );
  NOR3_X1 NOR3_111( .ZN(g11975), .A1(g10107), .A2(g10197), .A3(g10282) );
  NOR3_X1 NOR3_112( .ZN(g11979), .A1(g10114), .A2(g10202), .A3(g10288) );
  NOR3_X1 NOR3_113( .ZN(g11980), .A1(g10115), .A2(g10204), .A3(g10291) );
  NOR3_X1 NOR3_114( .ZN(g11981), .A1(g10117), .A2(g10207), .A3(g10294) );
  NOR3_X1 NOR3_115( .ZN(g11987), .A1(g10120), .A2(g10209), .A3(g10295) );
  NOR3_X1 NOR3_116( .ZN(g11988), .A1(g10123), .A2(g10211), .A3(g10298) );
  NOR3_X1 NOR3_117( .ZN(g11991), .A1(g10146), .A2(g10218), .A3(g10303) );
  NOR3_X1 NOR3_118( .ZN(g11992), .A1(g10150), .A2(g10221), .A3(g10308) );
  NOR3_X1 NOR3_119( .ZN(g11993), .A1(g10153), .A2(g10224), .A3(g10310) );
  NOR3_X1 NOR3_120( .ZN(g11999), .A1(g10166), .A2(g10250), .A3(g10319) );
  NOR3_X1 NOR3_121( .ZN(g12000), .A1(g10170), .A2(g10257), .A3(g10325) );
  NOR3_X1 NOR3_122( .ZN(g12005), .A1(g10174), .A2(g10261), .A3(g10328) );
  NOR3_X1 NOR3_123( .ZN(g12006), .A1(g10175), .A2(g10262), .A3(g10329) );
  NOR3_X1 NOR3_124( .ZN(g12008), .A1(g10183), .A2(g10270), .A3(g10351) );
  NOR3_X1 NOR3_125( .ZN(g12026), .A1(g10195), .A2(g10280), .A3(g10360) );
  NOR3_X1 NOR3_126( .ZN(g12033), .A1(g10199), .A2(g10284), .A3(g10362) );
  NOR3_X1 NOR3_127( .ZN(g12034), .A1(g10200), .A2(g10286), .A3(g10365) );
  NOR3_X1 NOR3_128( .ZN(g12035), .A1(g10203), .A2(g10289), .A3(g10367) );
  NOR3_X1 NOR3_129( .ZN(g12036), .A1(g10205), .A2(g10292), .A3(g10370) );
  NOR3_X1 NOR3_130( .ZN(g12043), .A1(g10210), .A2(g10296), .A3(g10372) );
  NOR3_X1 NOR3_131( .ZN(g12044), .A1(g10212), .A2(g10299), .A3(g10375) );
  NOR3_X1 NOR3_132( .ZN(g12048), .A1(g10219), .A2(g10304), .A3(g10381) );
  NOR3_X1 NOR3_133( .ZN(g12049), .A1(g10220), .A2(g10306), .A3(g10384) );
  NOR3_X1 NOR3_134( .ZN(g12050), .A1(g10222), .A2(g10309), .A3(g10387) );
  NOR3_X1 NOR3_135( .ZN(g12056), .A1(g10225), .A2(g10311), .A3(g10388) );
  NOR3_X1 NOR3_136( .ZN(g12057), .A1(g10228), .A2(g10313), .A3(g10391) );
  NOR3_X1 NOR3_137( .ZN(g12060), .A1(g10251), .A2(g10320), .A3(g10396) );
  NOR3_X1 NOR3_138( .ZN(g12061), .A1(g10255), .A2(g10323), .A3(g10401) );
  NOR3_X1 NOR3_139( .ZN(g12062), .A1(g10258), .A2(g10326), .A3(g10403) );
  NOR3_X1 NOR3_140( .ZN(g12068), .A1(g10271), .A2(g10352), .A3(g10412) );
  NOR3_X1 NOR3_141( .ZN(g12079), .A1(g10281), .A2(g10361), .A3(g10422) );
  NOR3_X1 NOR3_142( .ZN(g12080), .A1(g10285), .A2(g10363), .A3(g10430) );
  NOR3_X1 NOR3_143( .ZN(g12081), .A1(g10287), .A2(g10366), .A3(g10433) );
  NOR3_X1 NOR3_144( .ZN(g12082), .A1(g10290), .A2(g10368), .A3(g10435) );
  NOR3_X1 NOR3_145( .ZN(g12083), .A1(g10293), .A2(g10371), .A3(g10438) );
  NOR3_X1 NOR3_146( .ZN(g12090), .A1(g10297), .A2(g10373), .A3(g10439) );
  NOR3_X1 NOR3_147( .ZN(g12097), .A1(g10301), .A2(g10377), .A3(g10441) );
  NOR3_X1 NOR3_148( .ZN(g12098), .A1(g10302), .A2(g10379), .A3(g10444) );
  NOR3_X2 NOR3_149( .ZN(g12099), .A1(g10305), .A2(g10382), .A3(g10446) );
  NOR3_X2 NOR3_150( .ZN(g12100), .A1(g10307), .A2(g10385), .A3(g10449) );
  NOR3_X1 NOR3_151( .ZN(g12107), .A1(g10312), .A2(g10389), .A3(g10451) );
  NOR3_X1 NOR3_152( .ZN(g12108), .A1(g10314), .A2(g10392), .A3(g10454) );
  NOR3_X1 NOR3_153( .ZN(g12112), .A1(g10321), .A2(g10397), .A3(g10460) );
  NOR3_X1 NOR3_154( .ZN(g12113), .A1(g10322), .A2(g10399), .A3(g10463) );
  NOR3_X1 NOR3_155( .ZN(g12114), .A1(g10324), .A2(g10402), .A3(g10466) );
  NOR3_X1 NOR3_156( .ZN(g12120), .A1(g10327), .A2(g10404), .A3(g10467) );
  NOR3_X1 NOR3_157( .ZN(g12121), .A1(g10330), .A2(g10406), .A3(g10470) );
  NOR3_X1 NOR3_158( .ZN(g12124), .A1(g10353), .A2(g10413), .A3(g10475) );
  NOR3_X1 NOR3_159( .ZN(g12145), .A1(g10364), .A2(g10431), .A3(g10492) );
  NOR3_X1 NOR3_160( .ZN(g12146), .A1(g10369), .A2(g10436), .A3(g10496) );
  NOR3_X1 NOR3_161( .ZN(g12151), .A1(g10374), .A2(g10440), .A3(g10498) );
  NOR3_X1 NOR3_162( .ZN(g12152), .A1(g10378), .A2(g10442), .A3(g10506) );
  NOR3_X1 NOR3_163( .ZN(g12153), .A1(g10380), .A2(g10445), .A3(g10509) );
  NOR3_X1 NOR3_164( .ZN(g12154), .A1(g10383), .A2(g10447), .A3(g10511) );
  NOR3_X1 NOR3_165( .ZN(g12155), .A1(g10386), .A2(g10450), .A3(g10514) );
  NOR3_X1 NOR3_166( .ZN(g12162), .A1(g10390), .A2(g10452), .A3(g10515) );
  NOR3_X1 NOR3_167( .ZN(g12169), .A1(g10394), .A2(g10456), .A3(g10517) );
  NOR3_X1 NOR3_168( .ZN(g12170), .A1(g10395), .A2(g10458), .A3(g10520) );
  NOR3_X1 NOR3_169( .ZN(g12171), .A1(g10398), .A2(g10461), .A3(g10522) );
  NOR3_X1 NOR3_170( .ZN(g12172), .A1(g10400), .A2(g10464), .A3(g10525) );
  NOR3_X1 NOR3_171( .ZN(g12179), .A1(g10405), .A2(g10468), .A3(g10527) );
  NOR3_X1 NOR3_172( .ZN(g12180), .A1(g10407), .A2(g10471), .A3(g10530) );
  NOR3_X1 NOR3_173( .ZN(g12184), .A1(g10414), .A2(g10476), .A3(g10536) );
  NOR3_X1 NOR3_174( .ZN(g12185), .A1(g10415), .A2(g10478), .A3(g10539) );
  NOR3_X1 NOR3_175( .ZN(g12192), .A1(g10423), .A2(g10485), .A3(g10548) );
  NOR3_X1 NOR3_176( .ZN(g12193), .A1(g10432), .A2(g10493), .A3(g10555) );
  NOR3_X1 NOR3_177( .ZN(g12194), .A1(g10434), .A2(g10494), .A3(g10556) );
  NOR3_X1 NOR3_178( .ZN(g12195), .A1(g10437), .A2(g10497), .A3(g10558) );
  NOR3_X1 NOR3_179( .ZN(g12207), .A1(g10443), .A2(g10507), .A3(g10566) );
  NOR3_X1 NOR3_180( .ZN(g12208), .A1(g10448), .A2(g10512), .A3(g10570) );
  NOR3_X1 NOR3_181( .ZN(g12213), .A1(g10453), .A2(g10516), .A3(g10572) );
  NOR3_X1 NOR3_182( .ZN(g12214), .A1(g10457), .A2(g10518), .A3(g10580) );
  NOR3_X1 NOR3_183( .ZN(g12215), .A1(g10459), .A2(g10521), .A3(g10583) );
  NOR3_X1 NOR3_184( .ZN(g12216), .A1(g10462), .A2(g10523), .A3(g10585) );
  NOR3_X1 NOR3_185( .ZN(g12217), .A1(g10465), .A2(g10526), .A3(g10588) );
  NOR3_X1 NOR3_186( .ZN(g12224), .A1(g10469), .A2(g10528), .A3(g10589) );
  NOR3_X1 NOR3_187( .ZN(g12231), .A1(g10473), .A2(g10532), .A3(g10591) );
  NOR3_X1 NOR3_188( .ZN(g12232), .A1(g10474), .A2(g10534), .A3(g10594) );
  NOR3_X1 NOR3_189( .ZN(g12233), .A1(g10477), .A2(g10537), .A3(g10596) );
  NOR3_X1 NOR3_190( .ZN(g12234), .A1(g10479), .A2(g10540), .A3(g10599) );
  NOR3_X1 NOR3_191( .ZN(g12245), .A1(g10495), .A2(g10557), .A3(g10604) );
  NOR3_X1 NOR3_192( .ZN(g12247), .A1(g10499), .A2(g10559), .A3(g10605) );
  NOR3_X1 NOR3_193( .ZN(g12248), .A1(g10508), .A2(g10567), .A3(g10612) );
  NOR3_X1 NOR3_194( .ZN(g12249), .A1(g10510), .A2(g10568), .A3(g10613) );
  NOR3_X1 NOR3_195( .ZN(g12250), .A1(g10513), .A2(g10571), .A3(g10615) );
  NOR3_X1 NOR3_196( .ZN(g12262), .A1(g10519), .A2(g10581), .A3(g10623) );
  NOR3_X1 NOR3_197( .ZN(g12263), .A1(g10524), .A2(g10586), .A3(g10627) );
  NOR3_X1 NOR3_198( .ZN(g12268), .A1(g10529), .A2(g10590), .A3(g10629) );
  NOR3_X1 NOR3_199( .ZN(g12269), .A1(g10533), .A2(g10592), .A3(g10637) );
  NOR3_X1 NOR3_200( .ZN(g12270), .A1(g10535), .A2(g10595), .A3(g10640) );
  NOR3_X1 NOR3_201( .ZN(g12271), .A1(g10538), .A2(g10597), .A3(g10642) );
  NOR3_X1 NOR3_202( .ZN(g12272), .A1(g10541), .A2(g10600), .A3(g10645) );
  NOR3_X1 NOR3_203( .ZN(g12288), .A1(g10569), .A2(g10614), .A3(g10651) );
  NOR3_X1 NOR3_204( .ZN(g12290), .A1(g10573), .A2(g10616), .A3(g10652) );
  NOR3_X1 NOR3_205( .ZN(g12291), .A1(g10582), .A2(g10624), .A3(g10659) );
  NOR3_X1 NOR3_206( .ZN(g12292), .A1(g10584), .A2(g10625), .A3(g10660) );
  NOR3_X1 NOR3_207( .ZN(g12293), .A1(g10587), .A2(g10628), .A3(g10662) );
  NOR3_X1 NOR3_208( .ZN(g12305), .A1(g10593), .A2(g10638), .A3(g10670) );
  NOR3_X1 NOR3_209( .ZN(g12306), .A1(g10598), .A2(g10643), .A3(g10674) );
  NOR3_X1 NOR3_210( .ZN(g12324), .A1(g10626), .A2(g10661), .A3(g10681) );
  NOR3_X1 NOR3_211( .ZN(g12326), .A1(g10630), .A2(g10663), .A3(g10682) );
  NOR3_X1 NOR3_212( .ZN(g12327), .A1(g10639), .A2(g10671), .A3(g10689) );
  NOR3_X1 NOR3_213( .ZN(g12328), .A1(g10641), .A2(g10672), .A3(g10690) );
  NOR3_X1 NOR3_214( .ZN(g12329), .A1(g10644), .A2(g10675), .A3(g10692) );
  NOR3_X1 NOR3_215( .ZN(g12339), .A1(g10650), .A2(g10678), .A3(g10704) );
  NOR3_X1 NOR3_216( .ZN(g12352), .A1(g10673), .A2(g10691), .A3(g10710) );
  NOR3_X1 NOR3_217( .ZN(g12369), .A1(g10680), .A2(g10707), .A3(g10724) );
  NOR3_X1 NOR3_218( .ZN(g12388), .A1(g10709), .A2(g10727), .A3(g10745) );
  NOR3_X1 NOR3_219( .ZN(g12418), .A1(g10729), .A2(g10748), .A3(g10764) );
  NOR2_X1 NOR2_2( .ZN(g12431), .A1(g8580), .A2(g10730) );
  NOR2_X1 NOR2_3( .ZN(g12436), .A1(g8587), .A2(g10749) );
  NOR2_X1 NOR2_4( .ZN(g12441), .A1(g8594), .A2(g10767) );
  NOR2_X1 NOR2_5( .ZN(g12446), .A1(g8605), .A2(g10773) );
  NOR2_X1 NOR2_6( .ZN(g12451), .A1(g499), .A2(g8983) );
  NOR3_X1 NOR3_220( .ZN(g12457), .A1(g9009), .A2(g9033), .A3(g9048) );
  NOR3_X1 NOR3_221( .ZN(g12467), .A1(g9034), .A2(g9056), .A3(g9065) );
  NOR3_X1 NOR3_222( .ZN(g12482), .A1(g9057), .A2(g9073), .A3(g9082) );
  NOR3_X1 NOR3_223( .ZN(g12487), .A1(g10108), .A2(g10198), .A3(g10283) );
  NOR3_X1 NOR3_224( .ZN(g12499), .A1(g9074), .A2(g9090), .A3(g9101) );
  NOR3_X1 NOR3_225( .ZN(g12507), .A1(g10213), .A2(g10300), .A3(g10376) );
  NOR3_X1 NOR3_226( .ZN(g12524), .A1(g10315), .A2(g10393), .A3(g10455) );
  NOR3_X1 NOR3_227( .ZN(g12539), .A1(g10408), .A2(g10472), .A3(g10531) );
  NOR3_X1 NOR3_228( .ZN(g12698), .A1(g11347), .A2(g11420), .A3(g8327) );
  NOR3_X1 NOR3_229( .ZN(g12747), .A1(g11421), .A2(g8328), .A3(g8385) );
  NOR3_X1 NOR3_230( .ZN(g12755), .A1(g11431), .A2(g8339), .A3(g8394) );
  NOR2_X1 NOR2_7( .ZN(g12780), .A1(g9187), .A2(g9161) );
  NOR3_X1 NOR3_231( .ZN(g12781), .A1(g8329), .A2(g8386), .A3(g8431) );
  NOR3_X1 NOR3_232( .ZN(g12789), .A1(g8340), .A2(g8395), .A3(g8437) );
  NOR3_X1 NOR3_233( .ZN(g12797), .A1(g8350), .A2(g8406), .A3(g8446) );
  NOR3_X1 NOR3_234( .ZN(g12814), .A1(g8387), .A2(g8432), .A3(g8463) );
  NOR2_X1 NOR2_8( .ZN(g12819), .A1(g9248), .A2(g9203) );
  NOR3_X1 NOR3_235( .ZN(g12820), .A1(g8396), .A2(g8438), .A3(g8466) );
  NOR3_X1 NOR3_236( .ZN(g12828), .A1(g8407), .A2(g8447), .A3(g8472) );
  NOR3_X1 NOR3_237( .ZN(g12836), .A1(g8417), .A2(g8458), .A3(g8481) );
  NOR3_X1 NOR3_238( .ZN(g12849), .A1(g8433), .A2(g8464), .A3(g8485) );
  NOR3_X1 NOR3_239( .ZN(g12852), .A1(g8439), .A2(g8467), .A3(g8488) );
  NOR2_X1 NOR2_9( .ZN(g12857), .A1(g9326), .A2(g9264) );
  NOR3_X1 NOR3_240( .ZN(g12858), .A1(g8448), .A2(g8473), .A3(g8491) );
  NOR3_X1 NOR3_241( .ZN(g12866), .A1(g8459), .A2(g8482), .A3(g8497) );
  NOR3_X1 NOR3_242( .ZN(g12880), .A1(g8465), .A2(g8486), .A3(g8502) );
  NOR2_X1 NOR2_10( .ZN(g12883), .A1(g10038), .A2(g6284) );
  NOR3_X1 NOR3_243( .ZN(g12890), .A1(g8468), .A2(g8489), .A3(g8505) );
  NOR3_X1 NOR3_244( .ZN(g12893), .A1(g8474), .A2(g8492), .A3(g8508) );
  NOR2_X1 NOR2_11( .ZN(g12898), .A1(g9407), .A2(g9342) );
  NOR3_X1 NOR3_245( .ZN(g12899), .A1(g8483), .A2(g8498), .A3(g8511) );
  NOR3_X1 NOR3_246( .ZN(g12912), .A1(g8484), .A2(g8500), .A3(g8515) );
  NOR3_X1 NOR3_247( .ZN(g12913), .A1(g8487), .A2(g8503), .A3(g8518) );
  NOR3_X1 NOR3_248( .ZN(g12920), .A1(g8490), .A2(g8506), .A3(g8521) );
  NOR2_X1 NOR2_12( .ZN(g12923), .A1(g10147), .A2(g6421) );
  NOR3_X1 NOR3_249( .ZN(g12930), .A1(g8493), .A2(g8509), .A3(g8524) );
  NOR3_X1 NOR3_250( .ZN(g12933), .A1(g8499), .A2(g8512), .A3(g8527) );
  NOR3_X1 NOR3_251( .ZN(g12939), .A1(g8501), .A2(g8516), .A3(g8531) );
  NOR3_X1 NOR3_252( .ZN(g12941), .A1(g8504), .A2(g8519), .A3(g8534) );
  NOR3_X1 NOR3_253( .ZN(g12942), .A1(g8507), .A2(g8522), .A3(g8537) );
  NOR3_X1 NOR3_254( .ZN(g12949), .A1(g8510), .A2(g8525), .A3(g8540) );
  NOR2_X1 NOR2_13( .ZN(g12952), .A1(g10252), .A2(g6626) );
  NOR3_X1 NOR3_255( .ZN(g12959), .A1(g8513), .A2(g8528), .A3(g8543) );
  NOR3_X2 NOR3_256( .ZN(g12967), .A1(g8517), .A2(g8532), .A3(g8546) );
  NOR3_X2 NOR3_257( .ZN(g12968), .A1(g8520), .A2(g8535), .A3(g8548) );
  NOR3_X1 NOR3_258( .ZN(g12970), .A1(g8523), .A2(g8538), .A3(g8551) );
  NOR3_X1 NOR3_259( .ZN(g12971), .A1(g8526), .A2(g8541), .A3(g8554) );
  NOR3_X1 NOR3_260( .ZN(g12978), .A1(g8529), .A2(g8544), .A3(g8557) );
  NOR2_X1 NOR2_14( .ZN(g12981), .A1(g10354), .A2(g6890) );
  NOR3_X1 NOR3_261( .ZN(g12991), .A1(g8536), .A2(g8549), .A3(g8559) );
  NOR3_X1 NOR3_262( .ZN(g12992), .A1(g8539), .A2(g8552), .A3(g8561) );
  NOR3_X1 NOR3_263( .ZN(g12994), .A1(g8542), .A2(g8555), .A3(g8564) );
  NOR3_X1 NOR3_264( .ZN(g12995), .A1(g8545), .A2(g8558), .A3(g8567) );
  NOR3_X1 NOR3_265( .ZN(g13001), .A1(g8553), .A2(g8562), .A3(g8570) );
  NOR3_X1 NOR3_266( .ZN(g13002), .A1(g8556), .A2(g8565), .A3(g8572) );
  NOR3_X1 NOR3_267( .ZN(g13022), .A1(g8566), .A2(g8573), .A3(g8576) );
  NOR3_X1 NOR4_4_A( .ZN(extra4), .A1(g11481), .A2(g8045), .A3(g7928) );
  NOR2_X1 NOR4_4( .ZN(g13024), .A1(extra4), .A2(g7880) );
  NOR3_X1 NOR3_268( .ZN(g13111), .A1(g8601), .A2(g8612), .A3(g8621) );
  NOR3_X1 NOR3_269( .ZN(g13124), .A1(g8613), .A2(g8625), .A3(g8631) );
  NOR3_X1 NOR3_270( .ZN(g13135), .A1(g8626), .A2(g8635), .A3(g8650) );
  NOR3_X1 NOR3_271( .ZN(g13143), .A1(g8636), .A2(g8654), .A3(g8666) );
  NOR3_X1 NOR3_272( .ZN(g13149), .A1(g8676), .A2(g8687), .A3(g8703) );
  NOR3_X1 NOR3_273( .ZN(g13155), .A1(g8688), .A2(g8705), .A3(g8722) );
  NOR3_X1 NOR3_274( .ZN(g13160), .A1(g8704), .A2(g8717), .A3(g8751) );
  NOR3_X1 NOR3_275( .ZN(g13164), .A1(g8706), .A2(g8724), .A3(g8760) );
  NOR3_X1 NOR3_276( .ZN(g13171), .A1(g8723), .A2(g8755), .A3(g8774) );
  NOR3_X1 NOR3_277( .ZN(g13175), .A1(g8725), .A2(g8762), .A3(g8783) );
  NOR3_X1 NOR3_278( .ZN(g13182), .A1(g8761), .A2(g8778), .A3(g8797) );
  NOR3_X1 NOR3_279( .ZN(g13194), .A1(g8784), .A2(g8801), .A3(g8816) );
  NOR3_X1 NOR3_280( .ZN(g13228), .A1(g8841), .A2(g8861), .A3(g8892) );
  NOR3_X1 NOR3_281( .ZN(g13251), .A1(g8868), .A2(g8899), .A3(g8932) );
  NOR3_X1 NOR3_282( .ZN(g13274), .A1(g8906), .A2(g8939), .A3(g8972) );
  NOR3_X1 NOR4_5_A( .ZN(extra5), .A1(g11481), .A2(g11332), .A3(g11190) );
  NOR2_X1 NOR4_5( .ZN(g13286), .A1(extra5), .A2(g7880) );
  NOR3_X1 NOR3_283( .ZN(g13299), .A1(g8946), .A2(g8979), .A3(g9004) );
  NOR3_X1 NOR4_6_A( .ZN(extra6), .A1(g11481), .A2(g11332), .A3(g11190) );
  NOR2_X1 NOR4_6( .ZN(g13310), .A1(extra6), .A2(g11069) );
  NOR3_X1 NOR4_7_A( .ZN(extra7), .A1(g8183), .A2(g11332), .A3(g11190) );
  NOR2_X1 NOR4_7( .ZN(g13313), .A1(extra7), .A2(g7880) );
  NOR3_X1 NOR4_8_A( .ZN(extra8), .A1(g8183), .A2(g11332), .A3(g11190) );
  NOR2_X1 NOR4_8( .ZN(g13331), .A1(extra8), .A2(g11069) );
  NOR3_X1 NOR4_9_A( .ZN(extra9), .A1(g11481), .A2(g8045), .A3(g11190) );
  NOR2_X1 NOR4_9( .ZN(g13332), .A1(extra9), .A2(g7880) );
  NOR3_X1 NOR4_10_A( .ZN(extra10), .A1(g11481), .A2(g8045), .A3(g11190) );
  NOR2_X1 NOR4_10( .ZN(g13353), .A1(extra10), .A2(g11069) );
  NOR3_X1 NOR4_11_A( .ZN(extra11), .A1(g8183), .A2(g8045), .A3(g11190) );
  NOR2_X1 NOR4_11( .ZN(g13354), .A1(extra11), .A2(g7880) );
  NOR3_X1 NOR4_12_A( .ZN(extra12), .A1(g8183), .A2(g8045), .A3(g11190) );
  NOR2_X1 NOR4_12( .ZN(g13374), .A1(extra12), .A2(g11069) );
  NOR3_X1 NOR4_13_A( .ZN(extra13), .A1(g11481), .A2(g11332), .A3(g7928) );
  NOR2_X1 NOR4_13( .ZN(g13375), .A1(extra13), .A2(g7880) );
  NOR3_X1 NOR3_284( .ZN(g13378), .A1(g9026), .A2(g9047), .A3(g9061) );
  NOR3_X1 NOR4_14_A( .ZN(extra14), .A1(g11481), .A2(g11332), .A3(g7928) );
  NOR2_X1 NOR4_14( .ZN(g13401), .A1(extra14), .A2(g11069) );
  NOR3_X1 NOR4_15_A( .ZN(extra15), .A1(g8183), .A2(g11332), .A3(g7928) );
  NOR2_X1 NOR4_15( .ZN(g13404), .A1(extra15), .A2(g7880) );
  NOR2_X1 NOR2_15( .ZN(g15661), .A1(g11737), .A2(g7345) );
  NOR2_X1 NOR2_16( .ZN(g15797), .A1(g13305), .A2(g7143) );
  NOR2_X1 NOR2_17( .ZN(g15873), .A1(g11617), .A2(g7562) );
  NOR2_X1 NOR2_18( .ZN(g15959), .A1(g2814), .A2(g13082) );
  NOR2_X1 NOR2_19( .ZN(g15978), .A1(g11737), .A2(g7152) );
  NOR3_X1 NOR3_285( .ZN(g16020), .A1(g6200), .A2(g12457), .A3(g10952) );
  NOR3_X1 NOR3_286( .ZN(g16036), .A1(g6289), .A2(g12467), .A3(g10952) );
  NOR3_X1 NOR3_287( .ZN(g16058), .A1(g6426), .A2(g12482), .A3(g10952) );
  NOR3_X1 NOR3_288( .ZN(g16082), .A1(g10952), .A2(g6140), .A3(g12487) );
  NOR3_X1 NOR3_289( .ZN(g16094), .A1(g6631), .A2(g12499), .A3(g10952) );
  NOR3_X1 NOR3_290( .ZN(g16120), .A1(g10952), .A2(g6161), .A3(g12507) );
  NOR3_X1 NOR3_291( .ZN(g16171), .A1(g10952), .A2(g6188), .A3(g12524) );
  NOR3_X1 NOR3_292( .ZN(g16230), .A1(g10952), .A2(g6220), .A3(g12539) );
  NOR2_X1 NOR2_20( .ZN(g16498), .A1(g14158), .A2(g14347) );
  NOR2_X1 NOR2_21( .ZN(g16520), .A1(g14273), .A2(g14459) );
  NOR2_X1 NOR2_22( .ZN(g16551), .A1(g14395), .A2(g14546) );
  NOR3_X1 NOR3_293( .ZN(g16567), .A1(g15904), .A2(g15880), .A3(g15859) );
  NOR3_X1 NOR3_294( .ZN(g16570), .A1(g15904), .A2(g15880), .A3(g14630) );
  NOR2_X1 NOR2_23( .ZN(g16583), .A1(g14507), .A2(g14601) );
  NOR3_X1 NOR3_295( .ZN(g16591), .A1(g15933), .A2(g15913), .A3(g15890) );
  NOR3_X1 NOR3_296( .ZN(g16594), .A1(g15933), .A2(g15913), .A3(g14650) );
  NOR3_X1 NOR3_297( .ZN(g16611), .A1(g15962), .A2(g15942), .A3(g15923) );
  NOR3_X1 NOR3_298( .ZN(g16614), .A1(g15962), .A2(g15942), .A3(g14677) );
  NOR3_X1 NOR3_299( .ZN(g16629), .A1(g15981), .A2(g15971), .A3(g15952) );
  NOR3_X1 NOR3_300( .ZN(g16632), .A1(g15981), .A2(g15971), .A3(g14711) );
  NOR3_X1 NOR3_301( .ZN(g16643), .A1(g15904), .A2(g14642), .A3(g15859) );
  NOR2_X1 NOR2_24( .ZN(g16654), .A1(g14690), .A2(g12477) );
  NOR3_X1 NOR3_302( .ZN(g16655), .A1(g15933), .A2(g14669), .A3(g15890) );
  NOR2_X1 NOR2_25( .ZN(g16671), .A1(g14724), .A2(g12494) );
  NOR3_X1 NOR3_303( .ZN(g16672), .A1(g15962), .A2(g14703), .A3(g15923) );
  NOR2_X1 NOR2_26( .ZN(g16679), .A1(g14797), .A2(g14895) );
  NOR2_X1 NOR2_27( .ZN(g16692), .A1(g14752), .A2(g12514) );
  NOR3_X1 NOR3_304( .ZN(g16693), .A1(g15981), .A2(g14737), .A3(g15952) );
  NOR2_X1 NOR2_28( .ZN(g16705), .A1(g14849), .A2(g14976) );
  NOR2_X1 NOR2_29( .ZN(g16718), .A1(g14773), .A2(g12531) );
  NOR2_X1 NOR2_30( .ZN(g16736), .A1(g14922), .A2(g15065) );
  NOR2_X1 NOR2_31( .ZN(g16778), .A1(g15003), .A2(g15161) );
  NOR2_X1 NOR2_32( .ZN(g16802), .A1(g13469), .A2(g3897) );
  NOR2_X1 NOR2_33( .ZN(g16803), .A1(g15593), .A2(g12908) );
  NOR2_X1 NOR2_34( .ZN(g16823), .A1(g5362), .A2(g13469) );
  NOR2_X1 NOR2_35( .ZN(g16824), .A1(g15658), .A2(g12938) );
  NOR2_X1 NOR2_36( .ZN(g16829), .A1(g14956), .A2(g12564) );
  NOR2_X1 NOR2_37( .ZN(g16835), .A1(g15717), .A2(g12966) );
  NOR2_X1 NOR2_38( .ZN(g16841), .A1(g15021), .A2(g12607) );
  NOR2_X1 NOR2_39( .ZN(g16844), .A1(g15754), .A2(g12989) );
  NOR2_X1 NOR2_40( .ZN(g16845), .A1(g15755), .A2(g12990) );
  NOR2_X1 NOR2_41( .ZN(g16847), .A1(g15095), .A2(g12650) );
  NOR2_X2 NOR2_42( .ZN(g16851), .A1(g15781), .A2(g13000) );
  NOR2_X1 NOR2_43( .ZN(g16853), .A1(g15801), .A2(g13009) );
  NOR2_X1 NOR2_44( .ZN(g16854), .A1(g15802), .A2(g13010) );
  NOR2_X1 NOR2_45( .ZN(g16857), .A1(g15817), .A2(g13023) );
  NOR2_X1 NOR2_46( .ZN(g16860), .A1(g15828), .A2(g13031) );
  NOR2_X1 NOR2_47( .ZN(g16861), .A1(g15829), .A2(g13032) );
  NOR2_X1 NOR2_48( .ZN(g16866), .A1(g15840), .A2(g13042) );
  NOR2_X1 NOR2_49( .ZN(g16880), .A1(g15852), .A2(g13056) );
  NOR3_X1 NOR3_305( .ZN(g17012), .A1(g14657), .A2(g14642), .A3(g15859) );
  NOR3_X1 NOR3_306( .ZN(g17025), .A1(g15904), .A2(g15880), .A3(g15859) );
  NOR3_X1 NOR3_307( .ZN(g17042), .A1(g14691), .A2(g14669), .A3(g15890) );
  NOR3_X1 NOR3_308( .ZN(g17051), .A1(g14657), .A2(g15880), .A3(g14630) );
  NOR3_X1 NOR3_309( .ZN(g17059), .A1(g15933), .A2(g15913), .A3(g15890) );
  NOR3_X2 NOR3_310( .ZN(g17076), .A1(g14725), .A2(g14703), .A3(g15923) );
  NOR3_X1 NOR3_311( .ZN(g17086), .A1(g14691), .A2(g15913), .A3(g14650) );
  NOR3_X1 NOR3_312( .ZN(g17094), .A1(g15962), .A2(g15942), .A3(g15923) );
  NOR3_X1 NOR3_313( .ZN(g17111), .A1(g14753), .A2(g14737), .A3(g15952) );
  NOR3_X1 NOR3_314( .ZN(g17124), .A1(g14725), .A2(g15942), .A3(g14677) );
  NOR3_X1 NOR3_315( .ZN(g17132), .A1(g15981), .A2(g15971), .A3(g15952) );
  NOR3_X1 NOR3_316( .ZN(g17151), .A1(g14753), .A2(g15971), .A3(g14711) );
  NOR2_X1 NOR2_50( .ZN(g17186), .A1(g7949), .A2(g14144) );
  NOR2_X1 NOR2_51( .ZN(g17197), .A1(g8000), .A2(g14259) );
  NOR2_X1 NOR2_52( .ZN(g17204), .A1(g8075), .A2(g14381) );
  NOR2_X1 NOR2_53( .ZN(g17209), .A1(g8160), .A2(g14493) );
  NOR2_X1 NOR2_54( .ZN(g17213), .A1(g4326), .A2(g14442) );
  NOR2_X1 NOR2_55( .ZN(g17215), .A1(g15904), .A2(g14642) );
  NOR2_X1 NOR2_56( .ZN(g17216), .A1(g4495), .A2(g14529) );
  NOR2_X1 NOR2_57( .ZN(g17218), .A1(g15933), .A2(g14669) );
  NOR2_X1 NOR2_58( .ZN(g17219), .A1(g4671), .A2(g14584) );
  NOR2_X1 NOR2_59( .ZN(g17220), .A1(g15962), .A2(g14703) );
  NOR2_X1 NOR2_60( .ZN(g17221), .A1(g4848), .A2(g14618) );
  NOR2_X1 NOR2_61( .ZN(g17222), .A1(g15998), .A2(g16003) );
  NOR2_X1 NOR2_62( .ZN(g17223), .A1(g15981), .A2(g14737) );
  NOR2_X1 NOR2_63( .ZN(g17224), .A1(g16004), .A2(g16009) );
  NOR2_X1 NOR2_64( .ZN(g17225), .A1(g16008), .A2(g16015) );
  NOR2_X1 NOR2_65( .ZN(g17226), .A1(g16010), .A2(g16017) );
  NOR2_X1 NOR2_66( .ZN(g17228), .A1(g16016), .A2(g16029) );
  NOR2_X1 NOR2_67( .ZN(g17229), .A1(g16019), .A2(g16032) );
  NOR2_X1 NOR2_68( .ZN(g17234), .A1(g16028), .A2(g16045) );
  NOR2_X1 NOR2_69( .ZN(g17235), .A1(g16030), .A2(g16047) );
  NOR2_X1 NOR2_70( .ZN(g17236), .A1(g16033), .A2(g16051) );
  NOR2_X1 NOR2_71( .ZN(g17246), .A1(g16046), .A2(g16066) );
  NOR2_X1 NOR2_72( .ZN(g17247), .A1(g16050), .A2(g16070) );
  NOR2_X1 NOR2_73( .ZN(g17248), .A1(g16052), .A2(g16072) );
  NOR2_X1 NOR2_74( .ZN(g17269), .A1(g16067), .A2(g16100) );
  NOR2_X1 NOR2_75( .ZN(g17270), .A1(g16071), .A2(g16104) );
  NOR2_X1 NOR2_76( .ZN(g17271), .A1(g16073), .A2(g16106) );
  NOR2_X1 NOR2_77( .ZN(g17302), .A1(g16103), .A2(g16135) );
  NOR2_X1 NOR2_78( .ZN(g17303), .A1(g16105), .A2(g16137) );
  NOR2_X1 NOR2_79( .ZN(g17340), .A1(g16136), .A2(g16183) );
  NOR2_X1 NOR2_80( .ZN(g17341), .A1(g16138), .A2(g16185) );
  NOR2_X1 NOR2_81( .ZN(g17383), .A1(g16184), .A2(g16238) );
  NOR2_X1 NOR2_82( .ZN(g17429), .A1(g16239), .A2(g16288) );
  NOR2_X1 NOR2_83( .ZN(g17507), .A1(g16298), .A2(g13318) );
  NOR2_X1 NOR2_84( .ZN(g17896), .A1(g14352), .A2(g16020) );
  NOR2_X1 NOR2_85( .ZN(g18007), .A1(g14464), .A2(g16036) );
  NOR2_X1 NOR2_86( .ZN(g18085), .A1(g16085), .A2(g6363) );
  NOR2_X1 NOR2_87( .ZN(g18124), .A1(g14551), .A2(g16058) );
  NOR2_X1 NOR2_88( .ZN(g18201), .A1(g16123), .A2(g6568) );
  NOR2_X1 NOR2_89( .ZN(g18240), .A1(g14606), .A2(g16094) );
  NOR2_X2 NOR2_90( .ZN(g18308), .A1(g16174), .A2(g6832) );
  NOR2_X2 NOR2_91( .ZN(g18352), .A1(g16082), .A2(g14249) );
  NOR2_X2 NOR2_92( .ZN(g18401), .A1(g16233), .A2(g7134) );
  NOR2_X2 NOR2_93( .ZN(g18430), .A1(g16020), .A2(g14352) );
  NOR2_X1 NOR2_94( .ZN(g18447), .A1(g16120), .A2(g14371) );
  NOR2_X1 NOR2_95( .ZN(g18503), .A1(g16036), .A2(g14464) );
  NOR2_X1 NOR2_96( .ZN(g18520), .A1(g16171), .A2(g14483) );
  NOR2_X1 NOR2_97( .ZN(g18548), .A1(g14249), .A2(g16082) );
  NOR2_X1 NOR2_98( .ZN(g18567), .A1(g16058), .A2(g14551) );
  NOR2_X1 NOR2_99( .ZN(g18584), .A1(g16230), .A2(g14570) );
  NOR2_X1 NOR2_100( .ZN(g18590), .A1(g16439), .A2(g7522) );
  NOR2_X1 NOR2_101( .ZN(g18598), .A1(g14371), .A2(g16120) );
  NOR2_X2 NOR2_102( .ZN(g18617), .A1(g16094), .A2(g14606) );
  NOR2_X2 NOR2_103( .ZN(g18623), .A1(g15902), .A2(g2814) );
  NOR2_X1 NOR2_104( .ZN(g18626), .A1(g16463), .A2(g7549) );
  NOR2_X1 NOR2_105( .ZN(g18630), .A1(g14483), .A2(g16171) );
  NOR2_X1 NOR2_106( .ZN(g18639), .A1(g14570), .A2(g16230) );
  NOR2_X1 NOR2_107( .ZN(g18669), .A1(g13623), .A2(g13634) );
  NOR2_X1 NOR2_108( .ZN(g18678), .A1(g13625), .A2(g11771) );
  NOR2_X1 NOR2_109( .ZN(g18707), .A1(g13636), .A2(g11788) );
  NOR2_X1 NOR2_110( .ZN(g18719), .A1(g13643), .A2(g13656) );
  NOR2_X1 NOR2_111( .ZN(g18726), .A1(g13645), .A2(g11805) );
  NOR2_X1 NOR2_112( .ZN(g18743), .A1(g13648), .A2(g11814) );
  NOR2_X1 NOR2_113( .ZN(g18754), .A1(g13655), .A2(g11816) );
  NOR2_X1 NOR2_114( .ZN(g18755), .A1(g13871), .A2(g12274) );
  NOR2_X1 NOR2_115( .ZN(g18763), .A1(g13671), .A2(g11838) );
  NOR2_X1 NOR2_116( .ZN(g18780), .A1(g13674), .A2(g11847) );
  NOR2_X1 NOR2_117( .ZN(g18781), .A1(g13675), .A2(g11851) );
  NOR2_X1 NOR2_118( .ZN(g18782), .A1(g13676), .A2(g13705) );
  NOR2_X1 NOR2_119( .ZN(g18794), .A1(g13701), .A2(g11880) );
  NOR2_X1 NOR2_120( .ZN(g18803), .A1(g13704), .A2(g11885) );
  NOR2_X1 NOR2_121( .ZN(g18804), .A1(g13905), .A2(g12331) );
  NOR2_X1 NOR2_122( .ZN(g18820), .A1(g13738), .A2(g11922) );
  NOR2_X1 NOR2_123( .ZN(g18821), .A1(g13740), .A2(g11926) );
  NOR2_X1 NOR2_124( .ZN(g18835), .A1(g13788), .A2(g11966) );
  NOR2_X1 NOR2_125( .ZN(g18836), .A1(g13789), .A2(g11967) );
  NOR2_X1 NOR2_126( .ZN(g18837), .A1(g13998), .A2(g12376) );
  NOR2_X1 NOR2_127( .ZN(g18852), .A1(g13815), .A2(g12012) );
  NOR2_X1 NOR2_128( .ZN(g18866), .A1(g13834), .A2(g12069) );
  NOR2_X1 NOR2_129( .ZN(g18867), .A1(g13835), .A2(g12070) );
  NOR2_X1 NOR2_130( .ZN(g18868), .A1(g14143), .A2(g12419) );
  NOR2_X1 NOR2_131( .ZN(g18883), .A1(g13846), .A2(g12128) );
  NOR2_X1 NOR2_132( .ZN(g18885), .A1(g13847), .A2(g12129) );
  NOR2_X1 NOR2_133( .ZN(g18906), .A1(g13855), .A2(g12186) );
  NOR2_X1 NOR2_134( .ZN(g18907), .A1(g14336), .A2(g12429) );
  NOR2_X1 NOR2_135( .ZN(g18942), .A1(g13870), .A2(g12273) );
  NOR2_X1 NOR2_136( .ZN(g18957), .A1(g13884), .A2(g12307) );
  NOR2_X1 NOR2_137( .ZN(g18968), .A1(g13904), .A2(g12330) );
  NOR2_X1 NOR2_138( .ZN(g18975), .A1(g13944), .A2(g12353) );
  NOR2_X1 NOR2_139( .ZN(g19144), .A1(g17268), .A2(g14884) );
  NOR2_X1 NOR2_140( .ZN(g19149), .A1(g17339), .A2(g15020) );
  NOR2_X1 NOR2_141( .ZN(g19153), .A1(g17381), .A2(g15093) );
  NOR2_X1 NOR2_142( .ZN(g19154), .A1(g17382), .A2(g15094) );
  NOR2_X1 NOR2_143( .ZN(g19157), .A1(g17428), .A2(g15171) );
  NOR2_X1 NOR2_144( .ZN(g19160), .A1(g17446), .A2(g15178) );
  NOR2_X1 NOR2_145( .ZN(g19162), .A1(g17485), .A2(g15243) );
  NOR2_X1 NOR2_146( .ZN(g19163), .A1(g17486), .A2(g15244) );
  NOR2_X1 NOR2_147( .ZN(g19165), .A1(g17526), .A2(g15264) );
  NOR2_X1 NOR2_148( .ZN(g19167), .A1(g17556), .A2(g15320) );
  NOR2_X1 NOR2_149( .ZN(g19171), .A1(g17616), .A2(g15356) );
  NOR2_X1 NOR2_150( .ZN(g19172), .A1(g17635), .A2(g15388) );
  NOR2_X1 NOR2_151( .ZN(g19173), .A1(g17636), .A2(g15389) );
  NOR2_X1 NOR2_152( .ZN(g19177), .A1(g17713), .A2(g15442) );
  NOR2_X1 NOR2_153( .ZN(g19178), .A1(g17718), .A2(g15452) );
  NOR2_X1 NOR2_154( .ZN(g19179), .A1(g17719), .A2(g15453) );
  NOR2_X1 NOR2_155( .ZN(g19184), .A1(g17798), .A2(g15520) );
  NOR2_X1 NOR2_156( .ZN(g19219), .A1(g18165), .A2(g15753) );
  NOR2_X1 NOR2_157( .ZN(g20008), .A1(g18977), .A2(g7338) );
  NOR2_X1 NOR2_158( .ZN(g20054), .A1(g19001), .A2(g16867) );
  NOR2_X1 NOR2_159( .ZN(g20095), .A1(g16507), .A2(g16895) );
  NOR2_X1 NOR2_160( .ZN(g20120), .A1(g16529), .A2(g16924) );
  NOR2_X1 NOR2_161( .ZN(g20150), .A1(g16560), .A2(g16954) );
  NOR2_X1 NOR2_162( .ZN(g20153), .A1(g16536), .A2(g7583) );
  NOR2_X1 NOR2_163( .ZN(g20299), .A1(g16665), .A2(g16884) );
  NOR2_X1 NOR2_164( .ZN(g20310), .A1(g16850), .A2(g13654) );
  NOR2_X1 NOR2_165( .ZN(g20314), .A1(g13646), .A2(g16855) );
  NOR2_X1 NOR2_166( .ZN(g20318), .A1(g16686), .A2(g16913) );
  NOR2_X1 NOR2_167( .ZN(g20333), .A1(g13672), .A2(g16859) );
  NOR2_X1 NOR2_168( .ZN(g20337), .A1(g16712), .A2(g16943) );
  NOR2_X1 NOR2_169( .ZN(g20343), .A1(g16856), .A2(g13703) );
  NOR2_X1 NOR2_170( .ZN(g20353), .A1(g13702), .A2(g16864) );
  NOR2_X1 NOR2_171( .ZN(g20357), .A1(g16743), .A2(g16974) );
  NOR2_X1 NOR2_172( .ZN(g20375), .A1(g13739), .A2(g16879) );
  NOR2_X1 NOR2_173( .ZN(g20376), .A1(g16865), .A2(g13787) );
  NOR2_X1 NOR2_174( .ZN(g20417), .A1(g16907), .A2(g13833) );
  NOR2_X1 NOR2_175( .ZN(g20682), .A1(g19160), .A2(g10024) );
  NOR2_X1 NOR2_176( .ZN(g20717), .A1(g19165), .A2(g10133) );
  NOR2_X1 NOR2_177( .ZN(g20752), .A1(g19171), .A2(g10238) );
  NOR2_X1 NOR2_178( .ZN(g20789), .A1(g19177), .A2(g10340) );
  NOR2_X1 NOR2_179( .ZN(g20841), .A1(g14767), .A2(g19552) );
  NOR2_X1 NOR2_180( .ZN(g20874), .A1(g17301), .A2(g19594) );
  NOR2_X1 NOR2_181( .ZN(g20875), .A1(g19584), .A2(g17352) );
  NOR2_X1 NOR2_182( .ZN(g20876), .A1(g19585), .A2(g17353) );
  NOR2_X1 NOR2_183( .ZN(g20877), .A1(g3919), .A2(g19830) );
  NOR2_X1 NOR2_184( .ZN(g20878), .A1(g19600), .A2(g17395) );
  NOR2_X1 NOR2_185( .ZN(g20879), .A1(g19601), .A2(g17396) );
  NOR2_X1 NOR2_186( .ZN(g20880), .A1(g19602), .A2(g17397) );
  NOR2_X1 NOR2_187( .ZN(g20881), .A1(g19603), .A2(g17398) );
  NOR2_X1 NOR2_188( .ZN(g20882), .A1(g19614), .A2(g17408) );
  NOR2_X1 NOR2_189( .ZN(g20883), .A1(g19615), .A2(g17409) );
  NOR2_X1 NOR2_190( .ZN(g20884), .A1(g5394), .A2(g19830) );
  NOR2_X1 NOR2_191( .ZN(g20891), .A1(g19626), .A2(g17447) );
  NOR2_X1 NOR2_192( .ZN(g20892), .A1(g19627), .A2(g17448) );
  NOR2_X1 NOR2_193( .ZN(g20893), .A1(g19628), .A2(g17449) );
  NOR2_X1 NOR2_194( .ZN(g20894), .A1(g19629), .A2(g17450) );
  NOR2_X1 NOR2_195( .ZN(g20895), .A1(g19633), .A2(g17461) );
  NOR2_X1 NOR2_196( .ZN(g20896), .A1(g19634), .A2(g17462) );
  NOR2_X1 NOR2_197( .ZN(g20897), .A1(g19635), .A2(g17463) );
  NOR2_X1 NOR2_198( .ZN(g20898), .A1(g19636), .A2(g17464) );
  NOR2_X1 NOR2_199( .ZN(g20899), .A1(g19647), .A2(g17474) );
  NOR2_X1 NOR2_200( .ZN(g20900), .A1(g19648), .A2(g17475) );
  NOR2_X1 NOR2_201( .ZN(g20901), .A1(g19660), .A2(g17508) );
  NOR2_X1 NOR2_202( .ZN(g20902), .A1(g19661), .A2(g17509) );
  NOR2_X1 NOR2_203( .ZN(g20903), .A1(g19662), .A2(g17510) );
  NOR2_X1 NOR2_204( .ZN(g20910), .A1(g19666), .A2(g17527) );
  NOR2_X1 NOR2_205( .ZN(g20911), .A1(g19667), .A2(g17528) );
  NOR2_X1 NOR2_206( .ZN(g20912), .A1(g19668), .A2(g17529) );
  NOR2_X1 NOR2_207( .ZN(g20913), .A1(g19669), .A2(g17530) );
  NOR2_X1 NOR2_208( .ZN(g20914), .A1(g19673), .A2(g17541) );
  NOR2_X2 NOR2_209( .ZN(g20915), .A1(g19674), .A2(g17542) );
  NOR2_X2 NOR2_210( .ZN(g20916), .A1(g19675), .A2(g17543) );
  NOR2_X2 NOR2_211( .ZN(g20917), .A1(g19676), .A2(g17544) );
  NOR2_X2 NOR2_212( .ZN(g20918), .A1(g19687), .A2(g17554) );
  NOR2_X2 NOR2_213( .ZN(g20919), .A1(g19688), .A2(g17555) );
  NOR2_X2 NOR2_214( .ZN(g20920), .A1(g19691), .A2(g19726) );
  NOR2_X2 NOR2_215( .ZN(g20921), .A1(g19697), .A2(g17576) );
  NOR2_X2 NOR2_216( .ZN(g20922), .A1(g19698), .A2(g17577) );
  NOR2_X2 NOR2_217( .ZN(g20923), .A1(g19699), .A2(g17578) );
  NOR2_X2 NOR2_218( .ZN(g20924), .A1(g19700), .A2(g15257) );
  NOR2_X1 NOR2_219( .ZN(g20925), .A1(g19708), .A2(g17598) );
  NOR2_X1 NOR2_220( .ZN(g20926), .A1(g19709), .A2(g17599) );
  NOR2_X1 NOR2_221( .ZN(g20927), .A1(g19710), .A2(g17600) );
  NOR2_X1 NOR2_222( .ZN(g20934), .A1(g19714), .A2(g17617) );
  NOR2_X1 NOR2_223( .ZN(g20935), .A1(g19715), .A2(g17618) );
  NOR2_X1 NOR2_224( .ZN(g20936), .A1(g19716), .A2(g17619) );
  NOR2_X1 NOR2_225( .ZN(g20937), .A1(g19717), .A2(g17620) );
  NOR2_X1 NOR2_226( .ZN(g20938), .A1(g19721), .A2(g17631) );
  NOR2_X1 NOR2_227( .ZN(g20939), .A1(g19722), .A2(g17632) );
  NOR2_X1 NOR2_228( .ZN(g20940), .A1(g19723), .A2(g17633) );
  NOR2_X1 NOR2_229( .ZN(g20941), .A1(g19724), .A2(g17634) );
  NOR2_X1 NOR2_230( .ZN(g20944), .A1(g19731), .A2(g17652) );
  NOR2_X1 NOR2_231( .ZN(g20945), .A1(g19732), .A2(g17653) );
  NOR2_X1 NOR2_232( .ZN(g20946), .A1(g19733), .A2(g17654) );
  NOR2_X1 NOR2_233( .ZN(g20947), .A1(g19734), .A2(g15335) );
  NOR2_X1 NOR2_234( .ZN(g20948), .A1(g19735), .A2(g15336) );
  NOR2_X1 NOR2_235( .ZN(g20949), .A1(g19741), .A2(g17673) );
  NOR2_X1 NOR2_236( .ZN(g20950), .A1(g19742), .A2(g17674) );
  NOR2_X1 NOR2_237( .ZN(g20951), .A1(g19743), .A2(g17675) );
  NOR2_X1 NOR2_238( .ZN(g20952), .A1(g19744), .A2(g15349) );
  NOR2_X1 NOR2_239( .ZN(g20953), .A1(g19752), .A2(g17695) );
  NOR2_X1 NOR2_240( .ZN(g20954), .A1(g19753), .A2(g17696) );
  NOR2_X1 NOR2_241( .ZN(g20955), .A1(g19754), .A2(g17697) );
  NOR2_X1 NOR2_242( .ZN(g20962), .A1(g19758), .A2(g17714) );
  NOR2_X1 NOR2_243( .ZN(g20963), .A1(g19759), .A2(g17715) );
  NOR2_X1 NOR2_244( .ZN(g20964), .A1(g19760), .A2(g17716) );
  NOR2_X1 NOR2_245( .ZN(g20965), .A1(g19761), .A2(g17717) );
  NOR2_X1 NOR2_246( .ZN(g20966), .A1(g19765), .A2(g17734) );
  NOR2_X1 NOR2_247( .ZN(g20967), .A1(g19766), .A2(g17735) );
  NOR2_X1 NOR2_248( .ZN(g20968), .A1(g19767), .A2(g17736) );
  NOR2_X1 NOR2_249( .ZN(g20969), .A1(g19768), .A2(g15402) );
  NOR2_X1 NOR2_250( .ZN(g20970), .A1(g19769), .A2(g15403) );
  NOR2_X1 NOR2_251( .ZN(g20972), .A1(g19774), .A2(g17752) );
  NOR2_X1 NOR2_252( .ZN(g20973), .A1(g19775), .A2(g17753) );
  NOR2_X1 NOR2_253( .ZN(g20974), .A1(g19776), .A2(g17754) );
  NOR2_X1 NOR2_254( .ZN(g20975), .A1(g19777), .A2(g15421) );
  NOR2_X1 NOR2_255( .ZN(g20976), .A1(g19778), .A2(g15422) );
  NOR2_X1 NOR2_256( .ZN(g20977), .A1(g19784), .A2(g17773) );
  NOR2_X1 NOR2_257( .ZN(g20978), .A1(g19785), .A2(g17774) );
  NOR2_X1 NOR2_258( .ZN(g20979), .A1(g19786), .A2(g17775) );
  NOR2_X1 NOR2_259( .ZN(g20980), .A1(g19787), .A2(g15435) );
  NOR2_X1 NOR2_260( .ZN(g20981), .A1(g19795), .A2(g17795) );
  NOR2_X1 NOR2_261( .ZN(g20982), .A1(g19796), .A2(g17796) );
  NOR2_X1 NOR2_262( .ZN(g20983), .A1(g19797), .A2(g17797) );
  NOR2_X1 NOR2_263( .ZN(g20989), .A1(g19802), .A2(g17812) );
  NOR2_X1 NOR2_264( .ZN(g20990), .A1(g19803), .A2(g17813) );
  NOR2_X1 NOR2_265( .ZN(g20991), .A1(g19804), .A2(g17814) );
  NOR2_X1 NOR2_266( .ZN(g20992), .A1(g19805), .A2(g15470) );
  NOR2_X1 NOR2_267( .ZN(g20993), .A1(g19807), .A2(g17835) );
  NOR2_X1 NOR2_268( .ZN(g20994), .A1(g19808), .A2(g17836) );
  NOR2_X1 NOR2_269( .ZN(g20995), .A1(g19809), .A2(g17837) );
  NOR2_X1 NOR2_270( .ZN(g20996), .A1(g19810), .A2(g15486) );
  NOR2_X1 NOR2_271( .ZN(g20997), .A1(g19811), .A2(g15487) );
  NOR2_X1 NOR2_272( .ZN(g20999), .A1(g19816), .A2(g17853) );
  NOR2_X1 NOR2_273( .ZN(g21000), .A1(g19817), .A2(g17854) );
  NOR2_X1 NOR2_274( .ZN(g21001), .A1(g19818), .A2(g17855) );
  NOR2_X1 NOR2_275( .ZN(g21002), .A1(g19819), .A2(g15505) );
  NOR2_X1 NOR2_276( .ZN(g21003), .A1(g19820), .A2(g15506) );
  NOR2_X1 NOR2_277( .ZN(g21004), .A1(g19826), .A2(g17874) );
  NOR2_X1 NOR2_278( .ZN(g21005), .A1(g19827), .A2(g17875) );
  NOR2_X1 NOR2_279( .ZN(g21006), .A1(g19828), .A2(g17876) );
  NOR2_X1 NOR2_280( .ZN(g21007), .A1(g19829), .A2(g15519) );
  NOR2_X1 NOR2_281( .ZN(g21008), .A1(g19836), .A2(g17877) );
  NOR2_X1 NOR2_282( .ZN(g21009), .A1(g19839), .A2(g17900) );
  NOR2_X1 NOR2_283( .ZN(g21010), .A1(g19840), .A2(g17901) );
  NOR2_X1 NOR2_284( .ZN(g21011), .A1(g19841), .A2(g17902) );
  NOR2_X1 NOR2_285( .ZN(g21015), .A1(g19846), .A2(g17924) );
  NOR2_X1 NOR2_286( .ZN(g21016), .A1(g19847), .A2(g17925) );
  NOR2_X1 NOR2_287( .ZN(g21017), .A1(g19848), .A2(g17926) );
  NOR2_X1 NOR2_288( .ZN(g21018), .A1(g19849), .A2(g15556) );
  NOR2_X1 NOR2_289( .ZN(g21019), .A1(g19851), .A2(g17947) );
  NOR2_X1 NOR2_290( .ZN(g21020), .A1(g19852), .A2(g17948) );
  NOR2_X1 NOR2_291( .ZN(g21021), .A1(g19853), .A2(g17949) );
  NOR2_X1 NOR2_292( .ZN(g21022), .A1(g19854), .A2(g15572) );
  NOR2_X1 NOR2_293( .ZN(g21023), .A1(g19855), .A2(g15573) );
  NOR2_X1 NOR2_294( .ZN(g21025), .A1(g19860), .A2(g17965) );
  NOR2_X1 NOR2_295( .ZN(g21026), .A1(g19861), .A2(g17966) );
  NOR2_X1 NOR2_296( .ZN(g21027), .A1(g19862), .A2(g17967) );
  NOR2_X1 NOR2_297( .ZN(g21028), .A1(g19863), .A2(g15591) );
  NOR2_X1 NOR2_298( .ZN(g21029), .A1(g19864), .A2(g15592) );
  NOR2_X1 NOR2_299( .ZN(g21031), .A1(g19869), .A2(g17989) );
  NOR2_X1 NOR2_300( .ZN(g21032), .A1(g19870), .A2(g17990) );
  NOR2_X1 NOR2_301( .ZN(g21033), .A1(g19872), .A2(g18011) );
  NOR2_X1 NOR2_302( .ZN(g21034), .A1(g19873), .A2(g18012) );
  NOR2_X1 NOR2_303( .ZN(g21035), .A1(g19874), .A2(g18013) );
  NOR2_X1 NOR2_304( .ZN(g21039), .A1(g19879), .A2(g18035) );
  NOR2_X1 NOR2_305( .ZN(g21040), .A1(g19880), .A2(g18036) );
  NOR2_X1 NOR2_306( .ZN(g21041), .A1(g19881), .A2(g18037) );
  NOR2_X1 NOR2_307( .ZN(g21042), .A1(g19882), .A2(g15634) );
  NOR2_X1 NOR2_308( .ZN(g21043), .A1(g19884), .A2(g18058) );
  NOR2_X1 NOR2_309( .ZN(g21044), .A1(g19885), .A2(g18059) );
  NOR2_X1 NOR2_310( .ZN(g21045), .A1(g19886), .A2(g18060) );
  NOR2_X1 NOR2_311( .ZN(g21046), .A1(g19887), .A2(g15650) );
  NOR2_X1 NOR2_312( .ZN(g21047), .A1(g19888), .A2(g15651) );
  NOR2_X1 NOR2_313( .ZN(g21048), .A1(g19889), .A2(g18062) );
  NOR2_X1 NOR2_314( .ZN(g21051), .A1(g19895), .A2(g18088) );
  NOR2_X1 NOR2_315( .ZN(g21052), .A1(g19900), .A2(g18106) );
  NOR2_X1 NOR2_316( .ZN(g21053), .A1(g19901), .A2(g18107) );
  NOR2_X1 NOR2_317( .ZN(g21054), .A1(g19903), .A2(g18128) );
  NOR2_X1 NOR2_318( .ZN(g21055), .A1(g19904), .A2(g18129) );
  NOR2_X1 NOR2_319( .ZN(g21056), .A1(g19905), .A2(g18130) );
  NOR2_X1 NOR2_320( .ZN(g21060), .A1(g19910), .A2(g18152) );
  NOR2_X1 NOR2_321( .ZN(g21061), .A1(g19911), .A2(g18153) );
  NOR2_X1 NOR2_322( .ZN(g21062), .A1(g19912), .A2(g18154) );
  NOR2_X1 NOR2_323( .ZN(g21063), .A1(g19913), .A2(g15710) );
  NOR2_X1 NOR2_324( .ZN(g21065), .A1(g19914), .A2(g18169) );
  NOR2_X1 NOR2_325( .ZN(g21070), .A1(g19920), .A2(g18204) );
  NOR2_X1 NOR2_326( .ZN(g21071), .A1(g19925), .A2(g18222) );
  NOR2_X1 NOR2_327( .ZN(g21072), .A1(g19926), .A2(g18223) );
  NOR2_X1 NOR2_328( .ZN(g21073), .A1(g19928), .A2(g18244) );
  NOR2_X1 NOR2_329( .ZN(g21074), .A1(g19929), .A2(g18245) );
  NOR2_X1 NOR2_330( .ZN(g21075), .A1(g19930), .A2(g18246) );
  NOR2_X1 NOR2_331( .ZN(g21080), .A1(g19935), .A2(g18311) );
  NOR2_X1 NOR2_332( .ZN(g21081), .A1(g19940), .A2(g18329) );
  NOR2_X1 NOR2_333( .ZN(g21082), .A1(g19941), .A2(g18330) );
  NOR2_X1 NOR2_334( .ZN(g21083), .A1(g19943), .A2(g18333) );
  NOR2_X1 NOR2_335( .ZN(g21084), .A1(g20011), .A2(g20048) );
  NOR2_X1 NOR2_336( .ZN(g21094), .A1(g19952), .A2(g18404) );
  NOR3_X1 NOR3_317( .ZN(g21095), .A1(g20012), .A2(g20049), .A3(g20084) );
  NOR3_X1 NOR3_318( .ZN(g21096), .A1(g20013), .A2(g20051), .A3(g20087) );
  NOR3_X1 NOR3_319( .ZN(g21104), .A1(g20050), .A2(g20085), .A3(g20106) );
  NOR3_X1 NOR3_320( .ZN(g21105), .A1(g20052), .A2(g20088), .A3(g20109) );
  NOR3_X1 NOR3_321( .ZN(g21106), .A1(g20053), .A2(g20090), .A3(g20112) );
  NOR3_X1 NOR3_322( .ZN(g21116), .A1(g20086), .A2(g20107), .A3(g20131) );
  NOR3_X1 NOR3_323( .ZN(g21117), .A1(g20089), .A2(g20110), .A3(g20133) );
  NOR3_X1 NOR3_324( .ZN(g21118), .A1(g20091), .A2(g20113), .A3(g20136) );
  NOR3_X1 NOR3_325( .ZN(g21119), .A1(g20092), .A2(g20115), .A3(g20139) );
  NOR3_X1 NOR3_326( .ZN(g21133), .A1(g20108), .A2(g20132), .A3(g20156) );
  NOR3_X1 NOR3_327( .ZN(g21134), .A1(g20111), .A2(g20134), .A3(g20157) );
  NOR3_X1 NOR3_328( .ZN(g21135), .A1(g20114), .A2(g20137), .A3(g20160) );
  NOR3_X1 NOR3_329( .ZN(g21147), .A1(g20135), .A2(g20158), .A3(g20188) );
  NOR3_X1 NOR3_330( .ZN(g21148), .A1(g20138), .A2(g20161), .A3(g20190) );
  NOR2_X1 NOR2_337( .ZN(g21149), .A1(g20015), .A2(g19981) );
  NOR2_X1 NOR2_338( .ZN(g21167), .A1(g20159), .A2(g20189) );
  NOR3_X1 NOR3_331( .ZN(g21168), .A1(g20162), .A2(g20191), .A3(g20220) );
  NOR2_X1 NOR2_339( .ZN(g21169), .A1(g20057), .A2(g20019) );
  NOR2_X1 NOR2_340( .ZN(g21183), .A1(g20192), .A2(g20221) );
  NOR2_X1 NOR2_341( .ZN(g21189), .A1(g20098), .A2(g20061) );
  NOR2_X1 NOR2_342( .ZN(g21204), .A1(g20123), .A2(g20102) );
  NOR2_X1 NOR2_343( .ZN(g21211), .A1(g19240), .A2(g19230) );
  NOR2_X1 NOR2_344( .ZN(g21219), .A1(g19253), .A2(g19243) );
  NOR3_X1 NOR3_332( .ZN(g21227), .A1(g18414), .A2(g18485), .A3(g20295) );
  NOR2_X1 NOR2_345( .ZN(g21228), .A1(g19388), .A2(g17118) );
  NOR2_X1 NOR2_346( .ZN(g21230), .A1(g19266), .A2(g19256) );
  NOR2_X1 NOR2_347( .ZN(g21233), .A1(g19418), .A2(g17145) );
  NOR2_X1 NOR2_348( .ZN(g21235), .A1(g19281), .A2(g19269) );
  NOR2_X1 NOR2_349( .ZN(g21238), .A1(g19954), .A2(g5890) );
  NOR2_X1 NOR2_350( .ZN(g21242), .A1(g19455), .A2(g17168) );
  NOR2_X1 NOR2_351( .ZN(g21246), .A1(g19984), .A2(g5929) );
  NOR2_X1 NOR2_352( .ZN(g21250), .A1(g19482), .A2(g17183) );
  NOR2_X1 NOR2_353( .ZN(g21255), .A1(g20022), .A2(g5963) );
  NOR2_X1 NOR2_354( .ZN(g21263), .A1(g20064), .A2(g5992) );
  NOR2_X1 NOR2_355( .ZN(g21316), .A1(g20460), .A2(g16111) );
  NOR2_X1 NOR2_356( .ZN(g21331), .A1(g20472), .A2(g16153) );
  NOR2_X1 NOR2_357( .ZN(g21346), .A1(g20480), .A2(g13247) );
  NOR2_X1 NOR2_358( .ZN(g21364), .A1(g20486), .A2(g13266) );
  NOR2_X1 NOR2_359( .ZN(g21385), .A1(g20492), .A2(g13289) );
  NOR2_X2 NOR2_360( .ZN(g21407), .A1(g20499), .A2(g13316) );
  NOR2_X2 NOR2_361( .ZN(g21432), .A1(g20502), .A2(g13335) );
  NOR2_X2 NOR2_362( .ZN(g21435), .A1(g20503), .A2(g16385) );
  NOR2_X1 NOR2_363( .ZN(g21467), .A1(g20506), .A2(g13355) );
  NOR2_X1 NOR2_364( .ZN(g21470), .A1(g20512), .A2(g16417) );
  NOR2_X1 NOR2_365( .ZN(g21502), .A1(g20525), .A2(g16445) );
  NOR2_X1 NOR2_366( .ZN(g21615), .A1(g16567), .A2(g19957) );
  NOR3_X1 NOR3_333( .ZN(g21618), .A1(g20016), .A2(g14079), .A3(g14165) );
  NOR2_X1 NOR2_367( .ZN(g21636), .A1(g20473), .A2(g6513) );
  NOR2_X1 NOR2_368( .ZN(g21643), .A1(g16591), .A2(g19987) );
  NOR3_X1 NOR3_334( .ZN(g21646), .A1(g20058), .A2(g14194), .A3(g14280) );
  NOR2_X1 NOR2_369( .ZN(g21665), .A1(g20507), .A2(g18352) );
  NOR2_X1 NOR2_370( .ZN(g21667), .A1(g20481), .A2(g6777) );
  NOR2_X1 NOR2_371( .ZN(g21674), .A1(g16611), .A2(g20025) );
  NOR3_X2 NOR3_335( .ZN(g21677), .A1(g20099), .A2(g14309), .A3(g14402) );
  NOR2_X1 NOR2_372( .ZN(g21694), .A1(g20526), .A2(g18447) );
  NOR2_X1 NOR2_373( .ZN(g21696), .A1(g20487), .A2(g7079) );
  NOR2_X1 NOR2_374( .ZN(g21703), .A1(g16629), .A2(g20067) );
  NOR3_X1 NOR3_336( .ZN(g21706), .A1(g20124), .A2(g14431), .A3(g14514) );
  NOR2_X1 NOR2_375( .ZN(g21711), .A1(g19830), .A2(g15780) );
  NOR2_X1 NOR2_376( .ZN(g21730), .A1(g20545), .A2(g18520) );
  NOR2_X1 NOR2_377( .ZN(g21732), .A1(g20493), .A2(g7329) );
  NOR3_X1 NOR3_337( .ZN(g21738), .A1(g19444), .A2(g17893), .A3(g14079) );
  NOR2_X1 NOR2_378( .ZN(g21739), .A1(g20507), .A2(g18430) );
  NOR2_X1 NOR2_379( .ZN(g21756), .A1(g19070), .A2(g18584) );
  NOR3_X1 NOR3_338( .ZN(g21762), .A1(g19471), .A2(g18004), .A3(g14194) );
  NOR2_X1 NOR2_380( .ZN(g21763), .A1(g20526), .A2(g18503) );
  NOR3_X1 NOR3_339( .ZN(g21778), .A1(g19494), .A2(g18121), .A3(g14309) );
  NOR2_X1 NOR2_381( .ZN(g21779), .A1(g20545), .A2(g18567) );
  NOR3_X1 NOR3_340( .ZN(g21793), .A1(g19515), .A2(g18237), .A3(g14431) );
  NOR2_X1 NOR2_382( .ZN(g21794), .A1(g19070), .A2(g18617) );
  NOR2_X1 NOR2_383( .ZN(g21796), .A1(g19830), .A2(g13004) );
  NOR2_X1 NOR2_384( .ZN(g21842), .A1(g13609), .A2(g19150) );
  NOR2_X1 NOR2_385( .ZN(g21843), .A1(g13619), .A2(g19155) );
  NOR2_X1 NOR2_386( .ZN(g21845), .A1(g13631), .A2(g19161) );
  NOR2_X1 NOR2_387( .ZN(g21847), .A1(g13642), .A2(g19166) );
  NOR2_X1 NOR2_388( .ZN(g21851), .A1(g19252), .A2(g8842) );
  NOR2_X1 NOR2_389( .ZN(g21878), .A1(g16964), .A2(g19228) );
  NOR2_X1 NOR2_390( .ZN(g21880), .A1(g13854), .A2(g19236) );
  NOR2_X1 NOR2_391( .ZN(g21882), .A1(g13862), .A2(g19248) );
  NOR2_X1 NOR2_392( .ZN(g21884), .A1(g19260), .A2(g19284) );
  NOR2_X1 NOR2_393( .ZN(g21887), .A1(g13519), .A2(g19289) );
  NOR2_X1 NOR2_394( .ZN(g21889), .A1(g19285), .A2(g19316) );
  NOR2_X1 NOR2_395( .ZN(g21890), .A1(g13530), .A2(g19307) );
  NOR2_X1 NOR2_396( .ZN(g21893), .A1(g13541), .A2(g19328) );
  NOR2_X1 NOR2_397( .ZN(g21894), .A1(g19317), .A2(g19356) );
  NOR2_X1 NOR2_398( .ZN(g21901), .A1(g13552), .A2(g19355) );
  NOR2_X1 NOR2_399( .ZN(g21968), .A1(g21234), .A2(g19476) );
  NOR2_X1 NOR2_400( .ZN(g21969), .A1(g20895), .A2(g10133) );
  NOR2_X1 NOR2_401( .ZN(g21970), .A1(g17182), .A2(g21226) );
  NOR2_X1 NOR2_402( .ZN(g21971), .A1(g21243), .A2(g19499) );
  NOR2_X1 NOR2_403( .ZN(g21972), .A1(g20914), .A2(g10238) );
  NOR2_X1 NOR2_404( .ZN(g21973), .A1(g21251), .A2(g19520) );
  NOR2_X1 NOR2_405( .ZN(g21974), .A1(g20938), .A2(g10340) );
  NOR2_X1 NOR2_406( .ZN(g21975), .A1(g21245), .A2(g21259) );
  NOR3_X1 NOR3_341( .ZN(g21980), .A1(g21252), .A2(g19531), .A3(g19540) );
  NOR2_X1 NOR2_407( .ZN(g21981), .A1(g21254), .A2(g21267) );
  NOR3_X1 NOR3_342( .ZN(g21987), .A1(g21260), .A2(g19541), .A3(g19544) );
  NOR2_X1 NOR2_408( .ZN(g21988), .A1(g21262), .A2(g21276) );
  NOR3_X1 NOR3_343( .ZN(g22000), .A1(g21268), .A2(g19545), .A3(g19547) );
  NOR2_X1 NOR2_409( .ZN(g22001), .A1(g21270), .A2(g21283) );
  NOR3_X1 NOR3_344( .ZN(g22013), .A1(g21277), .A2(g19548), .A3(g19551) );
  NOR2_X1 NOR2_410( .ZN(g22025), .A1(g21284), .A2(g19549) );
  NOR2_X1 NOR2_411( .ZN(g22026), .A1(g21083), .A2(g18407) );
  NOR2_X1 NOR2_412( .ZN(g22027), .A1(g21290), .A2(g19553) );
  NOR2_X1 NOR2_413( .ZN(g22028), .A1(g21291), .A2(g19554) );
  NOR2_X1 NOR2_414( .ZN(g22029), .A1(g21292), .A2(g19555) );
  NOR2_X1 NOR2_415( .ZN(g22030), .A1(g21298), .A2(g19557) );
  NOR2_X1 NOR2_416( .ZN(g22031), .A1(g21299), .A2(g19558) );
  NOR2_X1 NOR2_417( .ZN(g22032), .A1(g21300), .A2(g19559) );
  NOR2_X2 NOR2_418( .ZN(g22033), .A1(g21301), .A2(g19560) );
  NOR2_X1 NOR2_419( .ZN(g22034), .A1(g21302), .A2(g19561) );
  NOR2_X1 NOR2_420( .ZN(g22035), .A1(g21303), .A2(g19562) );
  NOR2_X1 NOR2_421( .ZN(g22037), .A1(g21304), .A2(g19564) );
  NOR2_X1 NOR2_422( .ZN(g22038), .A1(g21305), .A2(g19565) );
  NOR2_X1 NOR2_423( .ZN(g22039), .A1(g21306), .A2(g19566) );
  NOR2_X1 NOR2_424( .ZN(g22040), .A1(g21307), .A2(g19567) );
  NOR2_X1 NOR2_425( .ZN(g22041), .A1(g21308), .A2(g19568) );
  NOR2_X1 NOR2_426( .ZN(g22042), .A1(g21309), .A2(g19569) );
  NOR2_X1 NOR2_427( .ZN(g22043), .A1(g21310), .A2(g19570) );
  NOR2_X1 NOR2_428( .ZN(g22044), .A1(g21311), .A2(g19571) );
  NOR2_X1 NOR2_429( .ZN(g22045), .A1(g21312), .A2(g19572) );
  NOR2_X1 NOR2_430( .ZN(g22047), .A1(g21313), .A2(g19574) );
  NOR2_X1 NOR2_431( .ZN(g22048), .A1(g21314), .A2(g19575) );
  NOR2_X1 NOR2_432( .ZN(g22049), .A1(g21315), .A2(g19576) );
  NOR2_X1 NOR2_433( .ZN(g22054), .A1(g21319), .A2(g19586) );
  NOR2_X1 NOR2_434( .ZN(g22055), .A1(g21320), .A2(g19587) );
  NOR2_X1 NOR2_435( .ZN(g22056), .A1(g21321), .A2(g19588) );
  NOR2_X1 NOR2_436( .ZN(g22057), .A1(g21322), .A2(g19589) );
  NOR2_X1 NOR2_437( .ZN(g22058), .A1(g21323), .A2(g19590) );
  NOR2_X1 NOR2_438( .ZN(g22059), .A1(g21324), .A2(g19591) );
  NOR2_X1 NOR2_439( .ZN(g22060), .A1(g21325), .A2(g19592) );
  NOR2_X1 NOR2_440( .ZN(g22061), .A1(g21326), .A2(g19593) );
  NOR2_X1 NOR2_441( .ZN(g22063), .A1(g21328), .A2(g19597) );
  NOR2_X1 NOR2_442( .ZN(g22064), .A1(g21329), .A2(g19598) );
  NOR2_X1 NOR2_443( .ZN(g22065), .A1(g21330), .A2(g19599) );
  NOR2_X1 NOR2_444( .ZN(g22066), .A1(g21334), .A2(g19604) );
  NOR2_X1 NOR2_445( .ZN(g22067), .A1(g21335), .A2(g19605) );
  NOR2_X1 NOR2_446( .ZN(g22068), .A1(g21336), .A2(g19606) );
  NOR2_X1 NOR2_447( .ZN(g22073), .A1(g21337), .A2(g19616) );
  NOR2_X1 NOR2_448( .ZN(g22074), .A1(g21338), .A2(g19617) );
  NOR2_X1 NOR2_449( .ZN(g22075), .A1(g21339), .A2(g19618) );
  NOR2_X1 NOR2_450( .ZN(g22076), .A1(g21340), .A2(g19619) );
  NOR2_X1 NOR2_451( .ZN(g22077), .A1(g21341), .A2(g19620) );
  NOR2_X1 NOR2_452( .ZN(g22078), .A1(g21342), .A2(g19621) );
  NOR2_X1 NOR2_453( .ZN(g22079), .A1(g21343), .A2(g19623) );
  NOR2_X1 NOR2_454( .ZN(g22080), .A1(g21344), .A2(g19624) );
  NOR2_X1 NOR2_455( .ZN(g22081), .A1(g21345), .A2(g19625) );
  NOR2_X1 NOR2_456( .ZN(g22087), .A1(g21349), .A2(g19630) );
  NOR2_X1 NOR2_457( .ZN(g22088), .A1(g21350), .A2(g19631) );
  NOR2_X1 NOR2_458( .ZN(g22089), .A1(g21351), .A2(g19632) );
  NOR2_X1 NOR2_459( .ZN(g22090), .A1(g21352), .A2(g19637) );
  NOR2_X1 NOR2_460( .ZN(g22091), .A1(g21353), .A2(g19638) );
  NOR2_X1 NOR2_461( .ZN(g22092), .A1(g21354), .A2(g19639) );
  NOR2_X1 NOR2_462( .ZN(g22097), .A1(g21355), .A2(g19649) );
  NOR2_X1 NOR2_463( .ZN(g22098), .A1(g21356), .A2(g19650) );
  NOR2_X1 NOR2_464( .ZN(g22099), .A1(g21357), .A2(g19651) );
  NOR2_X1 NOR2_465( .ZN(g22100), .A1(g21360), .A2(g19653) );
  NOR2_X1 NOR2_466( .ZN(g22101), .A1(g21361), .A2(g19654) );
  NOR2_X1 NOR2_467( .ZN(g22102), .A1(g21362), .A2(g19655) );
  NOR2_X1 NOR2_468( .ZN(g22103), .A1(g21363), .A2(g19656) );
  NOR2_X1 NOR2_469( .ZN(g22104), .A1(g21367), .A2(g19663) );
  NOR2_X1 NOR2_470( .ZN(g22105), .A1(g21368), .A2(g19664) );
  NOR2_X1 NOR2_471( .ZN(g22106), .A1(g21369), .A2(g19665) );
  NOR2_X1 NOR2_472( .ZN(g22112), .A1(g21370), .A2(g19670) );
  NOR2_X1 NOR2_473( .ZN(g22113), .A1(g21371), .A2(g19671) );
  NOR2_X1 NOR2_474( .ZN(g22114), .A1(g21372), .A2(g19672) );
  NOR2_X2 NOR2_475( .ZN(g22115), .A1(g21373), .A2(g19677) );
  NOR2_X1 NOR2_476( .ZN(g22116), .A1(g21374), .A2(g19678) );
  NOR2_X1 NOR2_477( .ZN(g22117), .A1(g21375), .A2(g19679) );
  NOR2_X1 NOR2_478( .ZN(g22122), .A1(g21378), .A2(g19692) );
  NOR2_X1 NOR2_479( .ZN(g22123), .A1(g21379), .A2(g19693) );
  NOR2_X1 NOR2_480( .ZN(g22124), .A1(g21380), .A2(g19694) );
  NOR2_X1 NOR2_481( .ZN(g22125), .A1(g21381), .A2(g19695) );
  NOR2_X1 NOR2_482( .ZN(g22126), .A1(g21389), .A2(g19701) );
  NOR2_X1 NOR2_483( .ZN(g22127), .A1(g21390), .A2(g19702) );
  NOR2_X1 NOR2_484( .ZN(g22128), .A1(g21391), .A2(g19703) );
  NOR2_X1 NOR2_485( .ZN(g22129), .A1(g21392), .A2(g19704) );
  NOR2_X1 NOR2_486( .ZN(g22130), .A1(g21393), .A2(g19711) );
  NOR2_X1 NOR2_487( .ZN(g22131), .A1(g21394), .A2(g19712) );
  NOR2_X1 NOR2_488( .ZN(g22132), .A1(g21395), .A2(g19713) );
  NOR2_X1 NOR2_489( .ZN(g22138), .A1(g21396), .A2(g19718) );
  NOR2_X1 NOR2_490( .ZN(g22139), .A1(g21397), .A2(g19719) );
  NOR2_X1 NOR2_491( .ZN(g22140), .A1(g21398), .A2(g19720) );
  NOR2_X1 NOR2_492( .ZN(g22141), .A1(g21401), .A2(g19727) );
  NOR2_X1 NOR2_493( .ZN(g22142), .A1(g21402), .A2(g19728) );
  NOR2_X1 NOR2_494( .ZN(g22143), .A1(g21403), .A2(g19729) );
  NOR2_X1 NOR2_495( .ZN(g22144), .A1(g21410), .A2(g19730) );
  NOR2_X1 NOR2_496( .ZN(g22145), .A1(g21411), .A2(g19736) );
  NOR2_X1 NOR2_497( .ZN(g22146), .A1(g21412), .A2(g19737) );
  NOR2_X1 NOR2_498( .ZN(g22147), .A1(g21413), .A2(g19738) );
  NOR2_X1 NOR2_499( .ZN(g22148), .A1(g21414), .A2(g19739) );
  NOR2_X1 NOR2_500( .ZN(g22149), .A1(g21419), .A2(g19745) );
  NOR2_X1 NOR2_501( .ZN(g22150), .A1(g21420), .A2(g19746) );
  NOR2_X1 NOR2_502( .ZN(g22151), .A1(g21421), .A2(g19747) );
  NOR2_X1 NOR2_503( .ZN(g22152), .A1(g21422), .A2(g19748) );
  NOR2_X1 NOR2_504( .ZN(g22153), .A1(g21423), .A2(g19755) );
  NOR2_X1 NOR2_505( .ZN(g22154), .A1(g21424), .A2(g19756) );
  NOR2_X1 NOR2_506( .ZN(g22155), .A1(g21425), .A2(g19757) );
  NOR2_X1 NOR2_507( .ZN(g22161), .A1(g21428), .A2(g19764) );
  NOR2_X1 NOR2_508( .ZN(g22162), .A1(g21438), .A2(g19770) );
  NOR2_X1 NOR2_509( .ZN(g22163), .A1(g21439), .A2(g19771) );
  NOR2_X1 NOR2_510( .ZN(g22164), .A1(g21440), .A2(g19772) );
  NOR2_X1 NOR2_511( .ZN(g22165), .A1(g21444), .A2(g19773) );
  NOR2_X1 NOR2_512( .ZN(g22166), .A1(g21445), .A2(g19779) );
  NOR2_X1 NOR2_513( .ZN(g22167), .A1(g21446), .A2(g19780) );
  NOR2_X1 NOR2_514( .ZN(g22168), .A1(g21447), .A2(g19781) );
  NOR2_X1 NOR2_515( .ZN(g22169), .A1(g21448), .A2(g19782) );
  NOR2_X1 NOR2_516( .ZN(g22170), .A1(g21453), .A2(g19788) );
  NOR2_X1 NOR2_517( .ZN(g22171), .A1(g21454), .A2(g19789) );
  NOR2_X1 NOR2_518( .ZN(g22172), .A1(g21455), .A2(g19790) );
  NOR2_X1 NOR2_519( .ZN(g22173), .A1(g21456), .A2(g19791) );
  NOR2_X1 NOR2_520( .ZN(g22174), .A1(g19868), .A2(g21593) );
  NOR2_X1 NOR2_521( .ZN(g22177), .A1(g21476), .A2(g19806) );
  NOR2_X1 NOR2_522( .ZN(g22178), .A1(g21480), .A2(g19812) );
  NOR2_X1 NOR2_523( .ZN(g22179), .A1(g21481), .A2(g19813) );
  NOR2_X1 NOR2_524( .ZN(g22180), .A1(g21482), .A2(g19814) );
  NOR2_X1 NOR2_525( .ZN(g22181), .A1(g21486), .A2(g19815) );
  NOR2_X1 NOR2_526( .ZN(g22182), .A1(g21487), .A2(g19821) );
  NOR2_X1 NOR2_527( .ZN(g22183), .A1(g21488), .A2(g19822) );
  NOR2_X1 NOR2_528( .ZN(g22184), .A1(g21489), .A2(g19823) );
  NOR2_X1 NOR2_529( .ZN(g22185), .A1(g21490), .A2(g19824) );
  NOR2_X1 NOR2_530( .ZN(g22186), .A1(g21497), .A2(g19837) );
  NOR2_X1 NOR2_531( .ZN(g22189), .A1(g19899), .A2(g21622) );
  NOR2_X1 NOR2_532( .ZN(g22191), .A1(g21517), .A2(g19850) );
  NOR2_X1 NOR2_533( .ZN(g22192), .A1(g21521), .A2(g19856) );
  NOR2_X1 NOR2_534( .ZN(g22193), .A1(g21522), .A2(g19857) );
  NOR2_X1 NOR2_535( .ZN(g22194), .A1(g21523), .A2(g19858) );
  NOR2_X1 NOR2_536( .ZN(g22195), .A1(g21527), .A2(g19859) );
  NOR2_X1 NOR2_537( .ZN(g22198), .A1(g19924), .A2(g21650) );
  NOR2_X1 NOR2_538( .ZN(g22200), .A1(g21553), .A2(g19883) );
  NOR2_X1 NOR2_539( .ZN(g22204), .A1(g19939), .A2(g21681) );
  NOR2_X1 NOR2_540( .ZN(g22210), .A1(g21610), .A2(g19932) );
  NOR2_X1 NOR2_541( .ZN(g22216), .A1(g21635), .A2(g19944) );
  NOR2_X1 NOR2_542( .ZN(g22218), .A1(g21639), .A2(g19949) );
  NOR2_X1 NOR2_543( .ZN(g22227), .A1(g21658), .A2(g19953) );
  NOR2_X1 NOR2_544( .ZN(g22231), .A1(g21666), .A2(g19971) );
  NOR2_X1 NOR2_545( .ZN(g22234), .A1(g21670), .A2(g19976) );
  NOR2_X1 NOR2_546( .ZN(g22242), .A1(g21687), .A2(g19983) );
  NOR2_X1 NOR2_547( .ZN(g22247), .A1(g21695), .A2(g20001) );
  NOR2_X1 NOR2_548( .ZN(g22249), .A1(g21699), .A2(g20006) );
  NOR2_X1 NOR2_549( .ZN(g22263), .A1(g21723), .A2(g20021) );
  NOR2_X1 NOR2_550( .ZN(g22267), .A1(g21731), .A2(g20039) );
  NOR2_X1 NOR2_551( .ZN(g22269), .A1(g21735), .A2(g20044) );
  NOR2_X1 NOR2_552( .ZN(g22280), .A1(g21749), .A2(g20063) );
  NOR2_X1 NOR2_553( .ZN(g22284), .A1(g21757), .A2(g20081) );
  NOR2_X1 NOR2_554( .ZN(g22288), .A1(g20144), .A2(g21805) );
  NOR2_X1 NOR2_555( .ZN(g22299), .A1(g21773), .A2(g20104) );
  NOR2_X1 NOR2_556( .ZN(g22308), .A1(g20182), .A2(g21812) );
  NOR2_X1 NOR2_557( .ZN(g22336), .A1(g20216), .A2(g21818) );
  NOR2_X1 NOR2_558( .ZN(g22361), .A1(g20246), .A2(g21822) );
  NOR2_X1 NOR2_559( .ZN(g22454), .A1(g17012), .A2(g21891) );
  NOR2_X1 NOR2_560( .ZN(g22493), .A1(g17042), .A2(g21899) );
  NOR2_X1 NOR2_561( .ZN(g22536), .A1(g17076), .A2(g21911) );
  NOR2_X1 NOR2_562( .ZN(g22576), .A1(g17111), .A2(g21925) );
  NOR2_X1 NOR2_563( .ZN(g22578), .A1(g21892), .A2(g18982) );
  NOR2_X1 NOR2_564( .ZN(g22615), .A1(g21900), .A2(g18990) );
  NOR2_X1 NOR2_565( .ZN(g22651), .A1(g21912), .A2(g18997) );
  NOR2_X1 NOR2_566( .ZN(g22687), .A1(g21926), .A2(g19010) );
  NOR2_X1 NOR2_567( .ZN(g22755), .A1(g21271), .A2(g20842) );
  NOR2_X1 NOR2_568( .ZN(g22784), .A1(g16075), .A2(g20885) );
  NOR2_X1 NOR2_569( .ZN(g22789), .A1(g21278), .A2(g20850) );
  NOR3_X1 NOR3_345( .ZN(g22810), .A1(g16075), .A2(g20842), .A3(g21271) );
  NOR2_X1 NOR2_570( .ZN(g22826), .A1(g16113), .A2(g20904) );
  NOR2_X1 NOR2_571( .ZN(g22831), .A1(g21285), .A2(g20858) );
  NOR3_X1 NOR3_346( .ZN(g22851), .A1(g16113), .A2(g20850), .A3(g21278) );
  NOR2_X1 NOR2_572( .ZN(g22865), .A1(g16164), .A2(g20928) );
  NOR2_X1 NOR2_573( .ZN(g22870), .A1(g21293), .A2(g20866) );
  NOR3_X1 NOR3_347( .ZN(g22886), .A1(g16164), .A2(g20858), .A3(g21285) );
  NOR2_X1 NOR2_574( .ZN(g22900), .A1(g16223), .A2(g20956) );
  NOR3_X1 NOR3_348( .ZN(g22921), .A1(g16223), .A2(g20866), .A3(g21293) );
  NOR2_X1 NOR2_575( .ZN(g22935), .A1(g21903), .A2(g7466) );
  NOR2_X1 NOR2_576( .ZN(g22953), .A1(g20700), .A2(g7595) );
  NOR2_X1 NOR2_577( .ZN(g22985), .A1(g21618), .A2(g21049) );
  NOR2_X1 NOR2_578( .ZN(g22987), .A1(g21646), .A2(g21068) );
  NOR2_X1 NOR2_579( .ZN(g22990), .A1(g21677), .A2(g21078) );
  NOR2_X1 NOR2_580( .ZN(g22997), .A1(g21706), .A2(g21092) );
  NOR2_X1 NOR2_581( .ZN(g22999), .A1(g21085), .A2(g19241) );
  NOR2_X1 NOR2_582( .ZN(g23000), .A1(g16909), .A2(g21067) );
  NOR2_X1 NOR2_583( .ZN(g23009), .A1(g21738), .A2(g21107) );
  NOR2_X2 NOR2_584( .ZN(g23013), .A1(g21097), .A2(g19254) );
  NOR2_X2 NOR2_585( .ZN(g23014), .A1(g16939), .A2(g21077) );
  NOR2_X1 NOR2_586( .ZN(g23022), .A1(g16968), .A2(g21086) );
  NOR3_X1 NOR3_349( .ZN(g23023), .A1(g14256), .A2(g14175), .A3(g21123) );
  NOR2_X1 NOR2_587( .ZN(g23025), .A1(g21762), .A2(g21124) );
  NOR2_X1 NOR2_588( .ZN(g23029), .A1(g21111), .A2(g19267) );
  NOR2_X1 NOR2_589( .ZN(g23030), .A1(g16970), .A2(g21091) );
  NOR2_X1 NOR2_590( .ZN(g23039), .A1(g16989), .A2(g21098) );
  NOR3_X1 NOR3_350( .ZN(g23040), .A1(g14378), .A2(g14290), .A3(g21142) );
  NOR2_X1 NOR2_591( .ZN(g23042), .A1(g21778), .A2(g21143) );
  NOR2_X1 NOR2_592( .ZN(g23046), .A1(g21128), .A2(g19282) );
  NOR2_X1 NOR2_593( .ZN(g23047), .A1(g16991), .A2(g21103) );
  NOR2_X1 NOR2_594( .ZN(g23051), .A1(g21121), .A2(g21153) );
  NOR2_X1 NOR2_595( .ZN(g23058), .A1(g16999), .A2(g21112) );
  NOR3_X1 NOR3_351( .ZN(g23059), .A1(g14490), .A2(g14412), .A3(g21162) );
  NOR2_X1 NOR2_596( .ZN(g23061), .A1(g21793), .A2(g21163) );
  NOR3_X1 NOR3_352( .ZN(g23066), .A1(g21138), .A2(g19303), .A3(g19320) );
  NOR2_X1 NOR2_597( .ZN(g23067), .A1(g17015), .A2(g21122) );
  NOR2_X1 NOR2_598( .ZN(g23070), .A1(g21140), .A2(g21173) );
  NOR2_X1 NOR2_599( .ZN(g23076), .A1(g17023), .A2(g21129) );
  NOR3_X1 NOR3_353( .ZN(g23077), .A1(g14577), .A2(g14524), .A3(g21182) );
  NOR3_X1 NOR3_354( .ZN(g23080), .A1(g21158), .A2(g19324), .A3(g19347) );
  NOR2_X1 NOR2_600( .ZN(g23081), .A1(g17045), .A2(g21141) );
  NOR2_X1 NOR2_601( .ZN(g23083), .A1(g21160), .A2(g21193) );
  NOR2_X1 NOR2_602( .ZN(g23092), .A1(g17055), .A2(g21154) );
  NOR2_X1 NOR2_603( .ZN(g23093), .A1(g17056), .A2(g21155) );
  NOR3_X1 NOR3_355( .ZN(g23096), .A1(g21178), .A2(g19351), .A3(g19381) );
  NOR2_X1 NOR2_604( .ZN(g23097), .A1(g17079), .A2(g21161) );
  NOR2_X1 NOR2_605( .ZN(g23099), .A1(g21180), .A2(g21208) );
  NOR2_X1 NOR2_606( .ZN(g23110), .A1(g17090), .A2(g21174) );
  NOR2_X1 NOR2_607( .ZN(g23111), .A1(g17091), .A2(g21175) );
  NOR3_X1 NOR3_356( .ZN(g23113), .A1(g21198), .A2(g19385), .A3(g19413) );
  NOR2_X1 NOR2_608( .ZN(g23114), .A1(g17114), .A2(g21181) );
  NOR2_X1 NOR2_609( .ZN(g23117), .A1(g17117), .A2(g21188) );
  NOR2_X1 NOR2_610( .ZN(g23123), .A1(g17128), .A2(g21194) );
  NOR2_X1 NOR2_611( .ZN(g23124), .A1(g17129), .A2(g21195) );
  NOR2_X1 NOR2_612( .ZN(g23126), .A1(g17144), .A2(g21203) );
  NOR2_X1 NOR2_613( .ZN(g23132), .A1(g17155), .A2(g21209) );
  NOR2_X1 NOR2_614( .ZN(g23133), .A1(g17156), .A2(g21210) );
  NOR2_X1 NOR2_615( .ZN(g23135), .A1(g21229), .A2(g19449) );
  NOR2_X1 NOR2_616( .ZN(g23136), .A1(g20878), .A2(g10024) );
  NOR2_X1 NOR2_617( .ZN(g23137), .A1(g17167), .A2(g21218) );
  NOR2_X1 NOR2_618( .ZN(g23324), .A1(g22144), .A2(g10024) );
  NOR2_X1 NOR2_619( .ZN(g23329), .A1(g22165), .A2(g10133) );
  NOR2_X1 NOR2_620( .ZN(g23330), .A1(g22186), .A2(g22777) );
  NOR2_X1 NOR2_621( .ZN(g23339), .A1(g22181), .A2(g10238) );
  NOR2_X1 NOR2_622( .ZN(g23348), .A1(g22195), .A2(g10340) );
  NOR2_X1 NOR2_623( .ZN(g23357), .A1(g22210), .A2(g20127) );
  NOR2_X1 NOR2_624( .ZN(g23358), .A1(g22227), .A2(g18407) );
  NOR2_X1 NOR2_625( .ZN(g23359), .A1(g22216), .A2(g22907) );
  NOR2_X1 NOR2_626( .ZN(g23385), .A1(g17393), .A2(g22517) );
  NOR2_X1 NOR2_627( .ZN(g23386), .A1(g22483), .A2(g21388) );
  NOR2_X1 NOR2_628( .ZN(g23392), .A1(g17460), .A2(g22557) );
  NOR2_X1 NOR2_629( .ZN(g23393), .A1(g22526), .A2(g21418) );
  NOR2_X1 NOR2_630( .ZN(g23399), .A1(g17506), .A2(g22581) );
  NOR2_X1 NOR2_631( .ZN(g23400), .A1(g17540), .A2(g22597) );
  NOR2_X1 NOR2_632( .ZN(g23401), .A1(g22566), .A2(g21452) );
  NOR2_X1 NOR2_633( .ZN(g23406), .A1(g17597), .A2(g22618) );
  NOR2_X1 NOR2_634( .ZN(g23407), .A1(g17630), .A2(g22634) );
  NOR2_X1 NOR2_635( .ZN(g23408), .A1(g22606), .A2(g21494) );
  NOR2_X1 NOR2_636( .ZN(g23413), .A1(g17694), .A2(g22654) );
  NOR2_X1 NOR2_637( .ZN(g23418), .A1(g17794), .A2(g22690) );
  NOR2_X1 NOR2_638( .ZN(g23427), .A1(g22699), .A2(g21589) );
  NOR2_X1 NOR2_639( .ZN(g23433), .A1(g22726), .A2(g21611) );
  NOR2_X1 NOR2_640( .ZN(g23461), .A1(g22841), .A2(g21707) );
  NOR2_X1 NOR2_641( .ZN(g23477), .A1(g22906), .A2(g21758) );
  NOR2_X1 NOR2_642( .ZN(g23497), .A1(g22876), .A2(g5606) );
  NOR2_X1 NOR2_643( .ZN(g23513), .A1(g22911), .A2(g5631) );
  NOR2_X1 NOR2_644( .ZN(g23528), .A1(g22936), .A2(g5659) );
  NOR2_X1 NOR2_645( .ZN(g23539), .A1(g22942), .A2(g5697) );
  NOR2_X2 NOR2_646( .ZN(g23545), .A1(g22984), .A2(g20285) );
  NOR3_X1 NOR3_357( .ZN(g23823), .A1(g23009), .A2(g18490), .A3(g4456) );
  NOR3_X1 NOR3_358( .ZN(g23858), .A1(g23025), .A2(g18554), .A3(g4632) );
  NOR3_X1 NOR3_359( .ZN(g23892), .A1(g23042), .A2(g18604), .A3(g4809) );
  NOR3_X1 NOR3_360( .ZN(g23913), .A1(g23061), .A2(g18636), .A3(g4985) );
  NOR2_X1 NOR2_647( .ZN(g23922), .A1(g4456), .A2(g22985) );
  NOR3_X1 NOR3_361( .ZN(g23945), .A1(g4456), .A2(g13565), .A3(g23009) );
  NOR2_X1 NOR2_648( .ZN(g23950), .A1(g22992), .A2(g6707) );
  NOR2_X1 NOR2_649( .ZN(g23954), .A1(g4632), .A2(g22987) );
  NOR3_X1 NOR3_362( .ZN(g23974), .A1(g4632), .A2(g13573), .A3(g23025) );
  NOR2_X1 NOR2_650( .ZN(g23979), .A1(g23003), .A2(g7009) );
  NOR2_X1 NOR2_651( .ZN(g23983), .A1(g4809), .A2(g22990) );
  NOR3_X1 NOR3_363( .ZN(g24004), .A1(g4809), .A2(g13582), .A3(g23042) );
  NOR2_X1 NOR2_652( .ZN(g24009), .A1(g23017), .A2(g7259) );
  NOR2_X1 NOR2_653( .ZN(g24013), .A1(g4985), .A2(g22997) );
  NOR3_X1 NOR3_364( .ZN(g24038), .A1(g4985), .A2(g13602), .A3(g23061) );
  NOR2_X1 NOR2_654( .ZN(g24043), .A1(g23033), .A2(g7455) );
  NOR2_X1 NOR2_655( .ZN(g24059), .A1(g21990), .A2(g20809) );
  NOR2_X1 NOR2_656( .ZN(g24072), .A1(g22004), .A2(g20826) );
  NOR2_X1 NOR2_657( .ZN(g24083), .A1(g22015), .A2(g20836) );
  NOR2_X1 NOR2_658( .ZN(g24092), .A1(g22020), .A2(g20840) );
  NOR2_X1 NOR2_659( .ZN(g24174), .A1(g16894), .A2(g22206) );
  NOR2_X1 NOR2_660( .ZN(g24178), .A1(g16908), .A2(g22211) );
  NOR2_X1 NOR2_661( .ZN(g24179), .A1(g16923), .A2(g22214) );
  NOR2_X1 NOR2_662( .ZN(g24181), .A1(g16938), .A2(g22220) );
  NOR2_X1 NOR2_663( .ZN(g24182), .A1(g16953), .A2(g22223) );
  NOR2_X1 NOR2_664( .ZN(g24206), .A1(g16966), .A2(g22228) );
  NOR2_X1 NOR2_665( .ZN(g24207), .A1(g16967), .A2(g22229) );
  NOR2_X1 NOR2_666( .ZN(g24208), .A1(g16969), .A2(g22235) );
  NOR2_X1 NOR2_667( .ZN(g24209), .A1(g16984), .A2(g22238) );
  NOR2_X1 NOR2_668( .ZN(g24212), .A1(g16987), .A2(g22244) );
  NOR2_X1 NOR2_669( .ZN(g24213), .A1(g16988), .A2(g22245) );
  NOR2_X1 NOR2_670( .ZN(g24214), .A1(g16990), .A2(g22250) );
  NOR2_X1 NOR2_671( .ZN(g24215), .A1(g16993), .A2(g22254) );
  NOR2_X1 NOR2_672( .ZN(g24216), .A1(g16994), .A2(g22255) );
  NOR2_X1 NOR2_673( .ZN(g24218), .A1(g16997), .A2(g22264) );
  NOR2_X1 NOR2_674( .ZN(g24219), .A1(g16998), .A2(g22265) );
  NOR2_X1 NOR2_675( .ZN(g24222), .A1(g17017), .A2(g22272) );
  NOR2_X1 NOR2_676( .ZN(g24223), .A1(g17018), .A2(g22273) );
  NOR2_X1 NOR2_677( .ZN(g24225), .A1(g17021), .A2(g22281) );
  NOR2_X1 NOR2_678( .ZN(g24226), .A1(g17022), .A2(g22282) );
  NOR2_X1 NOR2_679( .ZN(g24227), .A1(g22270), .A2(g21137) );
  NOR2_X1 NOR2_680( .ZN(g24228), .A1(g17028), .A2(g22285) );
  NOR2_X1 NOR2_681( .ZN(g24230), .A1(g17047), .A2(g22291) );
  NOR2_X1 NOR2_682( .ZN(g24231), .A1(g17048), .A2(g22292) );
  NOR2_X1 NOR2_683( .ZN(g24232), .A1(g22637), .A2(g22665) );
  NOR2_X1 NOR2_684( .ZN(g24234), .A1(g22289), .A2(g21157) );
  NOR2_X1 NOR2_685( .ZN(g24235), .A1(g17062), .A2(g22305) );
  NOR2_X1 NOR2_686( .ZN(g24237), .A1(g17081), .A2(g22311) );
  NOR2_X1 NOR2_687( .ZN(g24238), .A1(g17082), .A2(g22312) );
  NOR2_X1 NOR2_688( .ZN(g24242), .A1(g22309), .A2(g21177) );
  NOR2_X1 NOR2_689( .ZN(g24243), .A1(g17097), .A2(g22333) );
  NOR2_X1 NOR2_690( .ZN(g24249), .A1(g22337), .A2(g21197) );
  NOR2_X1 NOR2_691( .ZN(g24250), .A1(g17135), .A2(g22358) );
  NOR2_X1 NOR2_692( .ZN(g24426), .A1(g23386), .A2(g10024) );
  NOR2_X1 NOR2_693( .ZN(g24428), .A1(g23544), .A2(g22398) );
  NOR2_X1 NOR2_694( .ZN(g24430), .A1(g23393), .A2(g10133) );
  NOR2_X1 NOR2_695( .ZN(g24434), .A1(g23401), .A2(g10238) );
  NOR2_X1 NOR2_696( .ZN(g24438), .A1(g23408), .A2(g10340) );
  NOR2_X1 NOR2_697( .ZN(g24445), .A1(g23427), .A2(g22777) );
  NOR2_X1 NOR2_698( .ZN(g24446), .A1(g23433), .A2(g22907) );
  NOR2_X1 NOR2_699( .ZN(g24473), .A1(g23461), .A2(g18407) );
  NOR2_X1 NOR2_700( .ZN(g24476), .A1(g23477), .A2(g20127) );
  NOR2_X1 NOR2_701( .ZN(g24479), .A1(g23593), .A2(g22516) );
  NOR2_X1 NOR2_702( .ZN(g24480), .A1(g23617), .A2(g23659) );
  NOR2_X1 NOR2_703( .ZN(g24481), .A1(g23618), .A2(g19696) );
  NOR2_X1 NOR2_704( .ZN(g24485), .A1(g23625), .A2(g22556) );
  NOR2_X1 NOR2_705( .ZN(g24486), .A1(g23643), .A2(g22577) );
  NOR2_X1 NOR2_706( .ZN(g24487), .A1(g23666), .A2(g23709) );
  NOR2_X1 NOR2_707( .ZN(g24488), .A1(g23667), .A2(g19740) );
  NOR2_X1 NOR2_708( .ZN(g24489), .A1(g23674), .A2(g22596) );
  NOR2_X1 NOR2_709( .ZN(g24490), .A1(g23686), .A2(g22607) );
  NOR2_X1 NOR2_710( .ZN(g24491), .A1(g15247), .A2(g23735) );
  NOR2_X1 NOR2_711( .ZN(g24492), .A1(g23689), .A2(g22610) );
  NOR2_X1 NOR2_712( .ZN(g24493), .A1(g23693), .A2(g22614) );
  NOR2_X1 NOR2_713( .ZN(g24494), .A1(g23716), .A2(g23763) );
  NOR2_X1 NOR2_714( .ZN(g24495), .A1(g23717), .A2(g19783) );
  NOR2_X1 NOR2_715( .ZN(g24496), .A1(g23724), .A2(g22633) );
  NOR2_X1 NOR2_716( .ZN(g24497), .A1(g23734), .A2(g22638) );
  NOR2_X1 NOR2_717( .ZN(g24498), .A1(g15324), .A2(g23777) );
  NOR2_X1 NOR2_718( .ZN(g24499), .A1(g15325), .A2(g23778) );
  NOR2_X1 NOR2_719( .ZN(g24500), .A1(g23740), .A2(g22643) );
  NOR2_X1 NOR2_720( .ZN(g24501), .A1(g15339), .A2(g23790) );
  NOR2_X1 NOR2_721( .ZN(g24502), .A1(g23743), .A2(g22646) );
  NOR2_X1 NOR2_722( .ZN(g24503), .A1(g23747), .A2(g22650) );
  NOR2_X1 NOR2_723( .ZN(g24504), .A1(g23770), .A2(g23818) );
  NOR2_X1 NOR2_724( .ZN(g24505), .A1(g23771), .A2(g19825) );
  NOR2_X1 NOR2_725( .ZN(g24506), .A1(g23776), .A2(g22667) );
  NOR2_X1 NOR2_726( .ZN(g24507), .A1(g15391), .A2(g23824) );
  NOR2_X1 NOR2_727( .ZN(g24508), .A1(g15392), .A2(g23825) );
  NOR2_X1 NOR2_728( .ZN(g24509), .A1(g23789), .A2(g22674) );
  NOR2_X1 NOR2_729( .ZN(g24510), .A1(g15410), .A2(g23830) );
  NOR2_X1 NOR2_730( .ZN(g24511), .A1(g15411), .A2(g23831) );
  NOR2_X1 NOR2_731( .ZN(g24512), .A1(g23795), .A2(g22679) );
  NOR2_X1 NOR2_732( .ZN(g24513), .A1(g15425), .A2(g23843) );
  NOR2_X1 NOR2_733( .ZN(g24514), .A1(g23798), .A2(g22682) );
  NOR2_X1 NOR2_734( .ZN(g24515), .A1(g23802), .A2(g22686) );
  NOR2_X1 NOR2_735( .ZN(g24516), .A1(g23820), .A2(g22700) );
  NOR2_X1 NOR2_736( .ZN(g24517), .A1(g23822), .A2(g22701) );
  NOR2_X1 NOR2_737( .ZN(g24519), .A1(g15459), .A2(g23855) );
  NOR2_X1 NOR2_738( .ZN(g24520), .A1(g23829), .A2(g22707) );
  NOR2_X1 NOR2_739( .ZN(g24521), .A1(g15475), .A2(g23859) );
  NOR2_X1 NOR2_740( .ZN(g24522), .A1(g15476), .A2(g23860) );
  NOR2_X2 NOR2_741( .ZN(g24523), .A1(g23842), .A2(g22714) );
  NOR2_X2 NOR2_742( .ZN(g24524), .A1(g15494), .A2(g23865) );
  NOR2_X2 NOR2_743( .ZN(g24525), .A1(g15495), .A2(g23866) );
  NOR2_X1 NOR2_744( .ZN(g24526), .A1(g23848), .A2(g22719) );
  NOR2_X1 NOR2_745( .ZN(g24527), .A1(g15509), .A2(g23878) );
  NOR2_X1 NOR2_746( .ZN(g24528), .A1(g23851), .A2(g22722) );
  NOR2_X1 NOR2_747( .ZN(g24530), .A1(g23857), .A2(g22732) );
  NOR2_X1 NOR2_748( .ZN(g24532), .A1(g15545), .A2(g23889) );
  NOR2_X1 NOR2_749( .ZN(g24533), .A1(g23864), .A2(g22738) );
  NOR2_X1 NOR2_750( .ZN(g24534), .A1(g15561), .A2(g23893) );
  NOR2_X1 NOR2_751( .ZN(g24535), .A1(g15562), .A2(g23894) );
  NOR2_X1 NOR2_752( .ZN(g24536), .A1(g23877), .A2(g22745) );
  NOR2_X1 NOR2_753( .ZN(g24537), .A1(g15580), .A2(g23899) );
  NOR2_X1 NOR2_754( .ZN(g24538), .A1(g15581), .A2(g23900) );
  NOR2_X1 NOR2_755( .ZN(g24543), .A1(g23891), .A2(g22764) );
  NOR2_X1 NOR2_756( .ZN(g24545), .A1(g15623), .A2(g23910) );
  NOR2_X1 NOR2_757( .ZN(g24546), .A1(g23898), .A2(g22770) );
  NOR2_X1 NOR2_758( .ZN(g24547), .A1(g15639), .A2(g23914) );
  NOR2_X1 NOR2_759( .ZN(g24548), .A1(g15640), .A2(g23915) );
  NOR2_X1 NOR2_760( .ZN(g24555), .A1(g23912), .A2(g22798) );
  NOR2_X1 NOR2_761( .ZN(g24557), .A1(g15699), .A2(g23942) );
  NOR2_X1 NOR2_762( .ZN(g24558), .A1(g23917), .A2(g22804) );
  NOR2_X1 NOR2_763( .ZN(g24566), .A1(g23944), .A2(g22842) );
  NOR2_X1 NOR2_764( .ZN(g24575), .A1(g23972), .A2(g22874) );
  NOR2_X1 NOR2_765( .ZN(g24606), .A1(g24183), .A2(g537) );
  NOR2_X1 NOR2_766( .ZN(g24613), .A1(g23592), .A2(g22515) );
  NOR2_X1 NOR2_767( .ZN(g24622), .A1(g23616), .A2(g22546) );
  NOR2_X1 NOR2_768( .ZN(g24623), .A1(g24183), .A2(g529) );
  NOR2_X1 NOR2_769( .ZN(g24624), .A1(g23624), .A2(g22555) );
  NOR2_X1 NOR2_770( .ZN(g24636), .A1(g24183), .A2(g530) );
  NOR2_X1 NOR2_771( .ZN(g24637), .A1(g23665), .A2(g22587) );
  NOR2_X1 NOR2_772( .ZN(g24638), .A1(g23673), .A2(g22595) );
  NOR2_X1 NOR2_773( .ZN(g24652), .A1(g24183), .A2(g531) );
  NOR2_X1 NOR2_774( .ZN(g24656), .A1(g23715), .A2(g22624) );
  NOR2_X1 NOR2_775( .ZN(g24657), .A1(g23723), .A2(g22632) );
  NOR2_X1 NOR2_776( .ZN(g24663), .A1(g24183), .A2(g532) );
  NOR2_X1 NOR2_777( .ZN(g24675), .A1(g23769), .A2(g22660) );
  NOR2_X1 NOR2_778( .ZN(g24681), .A1(g24183), .A2(g533) );
  NOR2_X1 NOR2_779( .ZN(g24682), .A1(g23688), .A2(g24183) );
  NOR2_X1 NOR2_780( .ZN(g24694), .A1(g24183), .A2(g534) );
  NOR2_X1 NOR2_781( .ZN(g24708), .A1(g23854), .A2(g22727) );
  NOR2_X1 NOR2_782( .ZN(g24711), .A1(g24183), .A2(g536) );
  NOR2_X1 NOR2_783( .ZN(g24717), .A1(g23886), .A2(g22754) );
  NOR2_X1 NOR2_784( .ZN(g24720), .A1(g23888), .A2(g22759) );
  NOR2_X1 NOR2_785( .ZN(g24728), .A1(g23907), .A2(g22788) );
  NOR2_X1 NOR2_786( .ZN(g24731), .A1(g23909), .A2(g22793) );
  NOR2_X1 NOR2_787( .ZN(g24736), .A1(g23939), .A2(g22830) );
  NOR2_X1 NOR2_788( .ZN(g24739), .A1(g23941), .A2(g22835) );
  NOR2_X1 NOR2_789( .ZN(g24742), .A1(g23971), .A2(g22869) );
  NOR2_X1 NOR2_790( .ZN(g24756), .A1(g16089), .A2(g24211) );
  NOR2_X1 NOR2_791( .ZN(g24770), .A1(g16119), .A2(g24217) );
  NOR2_X1 NOR2_792( .ZN(g24782), .A1(g16160), .A2(g24221) );
  NOR2_X1 NOR2_793( .ZN(g24783), .A1(g16161), .A2(g24224) );
  NOR2_X1 NOR2_794( .ZN(g24800), .A1(g16211), .A2(g24229) );
  NOR2_X1 NOR2_795( .ZN(g24819), .A1(g16262), .A2(g24236) );
  NOR2_X1 NOR2_796( .ZN(g24836), .A1(g16309), .A2(g24241) );
  NOR2_X1 NOR2_797( .ZN(g24845), .A1(g16350), .A2(g24246) );
  NOR2_X1 NOR2_798( .ZN(g24847), .A1(g16356), .A2(g24247) );
  NOR2_X1 NOR2_799( .ZN(g24859), .A1(g16390), .A2(g24253) );
  NOR2_X1 NOR2_800( .ZN(g24871), .A1(g16422), .A2(g24256) );
  NOR2_X1 NOR2_801( .ZN(g25027), .A1(g24227), .A2(g17001) );
  NOR2_X1 NOR2_802( .ZN(g25042), .A1(g24234), .A2(g17031) );
  NOR2_X1 NOR2_803( .ZN(g25056), .A1(g24242), .A2(g17065) );
  NOR2_X1 NOR2_804( .ZN(g25067), .A1(g24249), .A2(g17100) );
  NOR2_X1 NOR2_805( .ZN(g25075), .A1(g13880), .A2(g23483) );
  NOR2_X1 NOR2_806( .ZN(g25076), .A1(g23409), .A2(g22187) );
  NOR2_X1 NOR2_807( .ZN(g25077), .A1(g23414), .A2(g22196) );
  NOR2_X1 NOR2_808( .ZN(g25078), .A1(g23419), .A2(g22201) );
  NOR2_X1 NOR2_809( .ZN(g25081), .A1(g23423), .A2(g22202) );
  NOR2_X1 NOR2_810( .ZN(g25082), .A1(g23428), .A2(g22207) );
  NOR2_X1 NOR2_811( .ZN(g25085), .A1(g23432), .A2(g22208) );
  NOR2_X1 NOR2_812( .ZN(g25091), .A1(g23434), .A2(g22215) );
  NOR2_X1 NOR2_813( .ZN(g25099), .A1(g23440), .A2(g22224) );
  NOR2_X1 NOR2_814( .ZN(g25125), .A1(g23510), .A2(g22340) );
  NOR2_X1 NOR2_815( .ZN(g25127), .A1(g23525), .A2(g22363) );
  NOR2_X1 NOR2_816( .ZN(g25129), .A1(g23536), .A2(g22383) );
  NOR2_X1 NOR2_817( .ZN(g25185), .A1(g24492), .A2(g10024) );
  NOR2_X1 NOR2_818( .ZN(g25189), .A1(g24502), .A2(g10133) );
  NOR2_X1 NOR2_819( .ZN(g25191), .A1(g24516), .A2(g22777) );
  NOR2_X1 NOR2_820( .ZN(g25194), .A1(g24514), .A2(g10238) );
  NOR2_X1 NOR2_821( .ZN(g25197), .A1(g24528), .A2(g10340) );
  NOR2_X1 NOR2_822( .ZN(g25199), .A1(g24558), .A2(g20127) );
  NOR2_X1 NOR2_823( .ZN(g25201), .A1(g24575), .A2(g18407) );
  NOR2_X1 NOR2_824( .ZN(g25202), .A1(g24566), .A2(g22907) );
  NOR2_X1 NOR2_825( .ZN(g25204), .A1(g24745), .A2(g23547) );
  NOR2_X1 NOR2_826( .ZN(g25206), .A1(g24746), .A2(g23550) );
  NOR2_X1 NOR2_827( .ZN(g25207), .A1(g24747), .A2(g23551) );
  NOR2_X1 NOR2_828( .ZN(g25208), .A1(g24748), .A2(g23552) );
  NOR2_X1 NOR2_829( .ZN(g25209), .A1(g24749), .A2(g23554) );
  NOR2_X1 NOR2_830( .ZN(g25211), .A1(g24750), .A2(g23558) );
  NOR2_X1 NOR2_831( .ZN(g25212), .A1(g24751), .A2(g23559) );
  NOR2_X1 NOR2_832( .ZN(g25213), .A1(g24752), .A2(g23560) );
  NOR2_X1 NOR2_833( .ZN(g25214), .A1(g24754), .A2(g23563) );
  NOR2_X1 NOR2_834( .ZN(g25215), .A1(g24755), .A2(g23564) );
  NOR2_X1 NOR2_835( .ZN(g25216), .A1(g24757), .A2(g23565) );
  NOR2_X1 NOR2_836( .ZN(g25217), .A1(g24758), .A2(g23567) );
  NOR2_X1 NOR2_837( .ZN(g25218), .A1(g24760), .A2(g23571) );
  NOR2_X1 NOR2_838( .ZN(g25219), .A1(g24761), .A2(g23572) );
  NOR2_X1 NOR2_839( .ZN(g25220), .A1(g24762), .A2(g23573) );
  NOR2_X1 NOR2_840( .ZN(g25221), .A1(g24767), .A2(g23577) );
  NOR2_X1 NOR2_841( .ZN(g25222), .A1(g24768), .A2(g23578) );
  NOR2_X1 NOR2_842( .ZN(g25223), .A1(g24769), .A2(g23579) );
  NOR2_X1 NOR2_843( .ZN(g25224), .A1(g24772), .A2(g23582) );
  NOR2_X1 NOR2_844( .ZN(g25225), .A1(g24773), .A2(g23583) );
  NOR2_X1 NOR2_845( .ZN(g25226), .A1(g24774), .A2(g23584) );
  NOR2_X1 NOR2_846( .ZN(g25227), .A1(g24775), .A2(g23586) );
  NOR2_X1 NOR2_847( .ZN(g25228), .A1(g24776), .A2(g23590) );
  NOR2_X1 NOR2_848( .ZN(g25229), .A1(g24777), .A2(g23591) );
  NOR2_X1 NOR2_849( .ZN(g25230), .A1(g24779), .A2(g23598) );
  NOR2_X1 NOR2_850( .ZN(g25231), .A1(g24780), .A2(g23599) );
  NOR2_X1 NOR2_851( .ZN(g25232), .A1(g24781), .A2(g23600) );
  NOR2_X1 NOR2_852( .ZN(g25233), .A1(g24788), .A2(g23604) );
  NOR2_X1 NOR2_853( .ZN(g25234), .A1(g24789), .A2(g23605) );
  NOR2_X1 NOR2_854( .ZN(g25235), .A1(g24790), .A2(g23606) );
  NOR2_X1 NOR2_855( .ZN(g25236), .A1(g24792), .A2(g23609) );
  NOR2_X1 NOR2_856( .ZN(g25237), .A1(g24793), .A2(g23610) );
  NOR2_X1 NOR2_857( .ZN(g25238), .A1(g24794), .A2(g23611) );
  NOR2_X1 NOR2_858( .ZN(g25239), .A1(g24796), .A2(g23615) );
  NOR2_X1 NOR2_859( .ZN(g25240), .A1(g24798), .A2(g23622) );
  NOR2_X1 NOR2_860( .ZN(g25241), .A1(g24799), .A2(g23623) );
  NOR2_X1 NOR2_861( .ZN(g25242), .A1(g24802), .A2(g23630) );
  NOR2_X1 NOR2_862( .ZN(g25243), .A1(g24803), .A2(g23631) );
  NOR2_X1 NOR2_863( .ZN(g25244), .A1(g24804), .A2(g23632) );
  NOR2_X1 NOR2_864( .ZN(g25245), .A1(g24809), .A2(g23636) );
  NOR2_X1 NOR2_865( .ZN(g25246), .A1(g24810), .A2(g23637) );
  NOR2_X1 NOR2_866( .ZN(g25247), .A1(g24811), .A2(g23638) );
  NOR2_X1 NOR2_867( .ZN(g25248), .A1(g24818), .A2(g23664) );
  NOR2_X1 NOR2_868( .ZN(g25249), .A1(g24821), .A2(g23671) );
  NOR2_X1 NOR2_869( .ZN(g25250), .A1(g24822), .A2(g23672) );
  NOR2_X1 NOR2_870( .ZN(g25251), .A1(g24824), .A2(g23679) );
  NOR2_X1 NOR2_871( .ZN(g25252), .A1(g24825), .A2(g23680) );
  NOR2_X1 NOR2_872( .ZN(g25253), .A1(g24826), .A2(g23681) );
  NOR2_X1 NOR2_873( .ZN(g25254), .A1(g24831), .A2(g23687) );
  NOR2_X1 NOR2_874( .ZN(g25255), .A1(g24838), .A2(g23714) );
  NOR2_X1 NOR2_875( .ZN(g25256), .A1(g24840), .A2(g23721) );
  NOR2_X1 NOR2_876( .ZN(g25257), .A1(g24841), .A2(g23722) );
  NOR2_X1 NOR2_877( .ZN(g25258), .A1(g24846), .A2(g23741) );
  NOR2_X1 NOR2_878( .ZN(g25259), .A1(g24853), .A2(g23768) );
  NOR2_X1 NOR2_879( .ZN(g25260), .A1(g24858), .A2(g17737) );
  NOR2_X1 NOR2_880( .ZN(g25261), .A1(g24861), .A2(g23796) );
  NOR2_X1 NOR2_881( .ZN(g25262), .A1(g24869), .A2(g17824) );
  NOR2_X1 NOR2_882( .ZN(g25263), .A1(g24874), .A2(g17838) );
  NOR2_X1 NOR2_883( .ZN(g25264), .A1(g24876), .A2(g23849) );
  NOR2_X1 NOR2_884( .ZN(g25265), .A1(g24878), .A2(g23852) );
  NOR2_X1 NOR2_885( .ZN(g25266), .A1(g24881), .A2(g17912) );
  NOR2_X1 NOR2_886( .ZN(g25267), .A1(g24884), .A2(g17936) );
  NOR2_X1 NOR2_887( .ZN(g25268), .A1(g24888), .A2(g17950) );
  NOR2_X1 NOR2_888( .ZN(g25270), .A1(g24898), .A2(g18023) );
  NOR2_X1 NOR2_889( .ZN(g25271), .A1(g24901), .A2(g18047) );
  NOR2_X1 NOR2_890( .ZN(g25272), .A1(g24905), .A2(g18061) );
  NOR2_X1 NOR2_891( .ZN(g25273), .A1(g24907), .A2(g23904) );
  NOR2_X1 NOR2_892( .ZN(g25279), .A1(g24921), .A2(g18140) );
  NOR2_X1 NOR2_893( .ZN(g25280), .A1(g24924), .A2(g18164) );
  NOR2_X1 NOR2_894( .ZN(g25288), .A1(g24938), .A2(g18256) );
  NOR2_X1 NOR2_895( .ZN(g25311), .A1(g24964), .A2(g24029) );
  NOR2_X1 NOR2_896( .ZN(g25343), .A1(g24975), .A2(g5623) );
  NOR2_X1 NOR2_897( .ZN(g25357), .A1(g24986), .A2(g5651) );
  NOR2_X1 NOR2_898( .ZN(g25372), .A1(g24997), .A2(g5689) );
  NOR2_X1 NOR2_899( .ZN(g25389), .A1(g25005), .A2(g5741) );
  NOR2_X1 NOR2_900( .ZN(g25418), .A1(g24482), .A2(g22319) );
  NOR2_X1 NOR2_901( .ZN(g25426), .A1(g24183), .A2(g24616) );
  NOR2_X1 NOR2_902( .ZN(g25429), .A1(g24482), .A2(g22319) );
  NOR2_X1 NOR2_903( .ZN(g25450), .A1(g16018), .A2(g25086) );
  NOR2_X1 NOR2_904( .ZN(g25451), .A1(g16048), .A2(g25102) );
  NOR2_X1 NOR2_905( .ZN(g25452), .A1(g16101), .A2(g25117) );
  NOR2_X1 NOR2_906( .ZN(g25523), .A1(g20842), .A2(g24429) );
  NOR2_X1 NOR2_907( .ZN(g25539), .A1(g25088), .A2(g6157) );
  NOR2_X1 NOR2_908( .ZN(g25569), .A1(g24708), .A2(g24490) );
  NOR2_X1 NOR2_909( .ZN(g25589), .A1(g20850), .A2(g24433) );
  NOR2_X1 NOR2_910( .ZN(g25605), .A1(g25096), .A2(g6184) );
  NOR2_X1 NOR2_911( .ZN(g25631), .A1(g24717), .A2(g24497) );
  NOR2_X1 NOR2_912( .ZN(g25648), .A1(g24720), .A2(g24500) );
  NOR2_X1 NOR2_913( .ZN(g25668), .A1(g20858), .A2(g24437) );
  NOR2_X1 NOR2_914( .ZN(g25684), .A1(g25106), .A2(g6216) );
  NOR2_X2 NOR2_915( .ZN(g25699), .A1(g24613), .A2(g24506) );
  NOR2_X2 NOR2_916( .ZN(g25708), .A1(g24728), .A2(g24509) );
  NOR2_X2 NOR2_917( .ZN(g25725), .A1(g24731), .A2(g24512) );
  NOR2_X1 NOR2_918( .ZN(g25745), .A1(g20866), .A2(g24440) );
  NOR2_X1 NOR2_919( .ZN(g25761), .A1(g25112), .A2(g6305) );
  NOR2_X1 NOR2_920( .ZN(g25764), .A1(g25076), .A2(g21615) );
  NOR2_X1 NOR2_921( .ZN(g25772), .A1(g24624), .A2(g24520) );
  NOR2_X1 NOR2_922( .ZN(g25781), .A1(g24736), .A2(g24523) );
  NOR2_X1 NOR2_923( .ZN(g25798), .A1(g24739), .A2(g24526) );
  NOR2_X1 NOR2_924( .ZN(g25818), .A1(g25077), .A2(g21643) );
  NOR2_X1 NOR2_925( .ZN(g25826), .A1(g24638), .A2(g24533) );
  NOR2_X1 NOR2_926( .ZN(g25835), .A1(g24742), .A2(g24536) );
  NOR3_X1 NOR3_365( .ZN(g25852), .A1(g4456), .A2(g14831), .A3(g25078) );
  NOR2_X1 NOR2_927( .ZN(g25853), .A1(g25081), .A2(g21674) );
  NOR2_X1 NOR2_928( .ZN(g25861), .A1(g24657), .A2(g24546) );
  NOR3_X1 NOR4_16_A( .ZN(extra16), .A1(g4456), .A2(g25078), .A3(g18429) );
  NOR2_X1 NOR4_16( .ZN(g25870), .A1(extra16), .A2(g16075) );
  NOR3_X1 NOR3_366( .ZN(g25873), .A1(g4632), .A2(g14904), .A3(g25082) );
  NOR2_X1 NOR2_929( .ZN(g25874), .A1(g25085), .A2(g21703) );
  NOR3_X1 NOR4_17_A( .ZN(extra17), .A1(g4632), .A2(g25082), .A3(g18502) );
  NOR2_X1 NOR4_17( .ZN(g25882), .A1(extra17), .A2(g16113) );
  NOR3_X1 NOR3_367( .ZN(g25885), .A1(g4809), .A2(g14985), .A3(g25091) );
  NOR3_X1 NOR4_18_A( .ZN(extra18), .A1(g4809), .A2(g25091), .A3(g18566) );
  NOR2_X1 NOR4_18( .ZN(g25887), .A1(extra18), .A2(g16164) );
  NOR3_X1 NOR3_368( .ZN(g25890), .A1(g4985), .A2(g15074), .A3(g25099) );
  NOR3_X1 NOR4_19_A( .ZN(extra19), .A1(g4985), .A2(g25099), .A3(g18616) );
  NOR2_X1 NOR4_19( .ZN(g25892), .A1(extra19), .A2(g16223) );
  NOR2_X1 NOR2_930( .ZN(g25932), .A1(g25125), .A2(g17001) );
  NOR2_X1 NOR2_931( .ZN(g25935), .A1(g25127), .A2(g17031) );
  NOR2_X1 NOR2_932( .ZN(g25938), .A1(g25129), .A2(g17065) );
  NOR2_X1 NOR2_933( .ZN(g25940), .A1(g24428), .A2(g17100) );
  NOR2_X1 NOR2_934( .ZN(g25941), .A1(g24529), .A2(g24540) );
  NOR2_X1 NOR2_935( .ZN(g25943), .A1(g24541), .A2(g24550) );
  NOR2_X1 NOR2_936( .ZN(g25944), .A1(g24542), .A2(g24552) );
  NOR2_X1 NOR2_937( .ZN(g25946), .A1(g24553), .A2(g24561) );
  NOR2_X1 NOR2_938( .ZN(g25947), .A1(g24554), .A2(g24563) );
  NOR2_X1 NOR2_939( .ZN(g25948), .A1(g24564), .A2(g24571) );
  NOR2_X1 NOR2_940( .ZN(g25949), .A1(g24565), .A2(g24573) );
  NOR2_X1 NOR2_941( .ZN(g25950), .A1(g24574), .A2(g24580) );
  NOR2_X1 NOR2_942( .ZN(g25962), .A1(g24591), .A2(g23496) );
  NOR2_X1 NOR2_943( .ZN(g25967), .A1(g24596), .A2(g23512) );
  NOR2_X1 NOR2_944( .ZN(g25974), .A1(g24604), .A2(g23527) );
  NOR2_X1 NOR2_945( .ZN(g25979), .A1(g24611), .A2(g23538) );
  NOR2_X1 NOR2_946( .ZN(g26025), .A1(g25392), .A2(g17193) );
  NOR2_X1 NOR2_947( .ZN(g26031), .A1(g25273), .A2(g22777) );
  NOR2_X1 NOR2_948( .ZN(g26037), .A1(g25311), .A2(g18407) );
  NOR2_X1 NOR2_949( .ZN(g26041), .A1(g25475), .A2(g24855) );
  NOR2_X1 NOR2_950( .ZN(g26042), .A1(g25505), .A2(g24867) );
  NOR2_X1 NOR2_951( .ZN(g26043), .A1(g25506), .A2(g24870) );
  NOR2_X1 NOR2_952( .ZN(g26044), .A1(g25552), .A2(g24882) );
  NOR2_X1 NOR2_953( .ZN(g26045), .A1(g25553), .A2(g24885) );
  NOR2_X1 NOR2_954( .ZN(g26046), .A1(g25618), .A2(g24899) );
  NOR2_X1 NOR2_955( .ZN(g26047), .A1(g25619), .A2(g24902) );
  NOR2_X1 NOR2_956( .ZN(g26048), .A1(g25628), .A2(g24906) );
  NOR2_X1 NOR2_957( .ZN(g26049), .A1(g25629), .A2(g24908) );
  NOR2_X1 NOR2_958( .ZN(g26050), .A1(g25697), .A2(g24922) );
  NOR2_X1 NOR2_959( .ZN(g26055), .A1(g25881), .A2(g24974) );
  NOR2_X1 NOR2_960( .ZN(g26081), .A1(g25470), .A2(g25482) );
  NOR2_X1 NOR2_961( .ZN(g26083), .A1(g25426), .A2(g22319) );
  NOR2_X1 NOR2_962( .ZN(g26084), .A1(g25487), .A2(g25513) );
  NOR3_X1 NOR3_369( .ZN(g26087), .A1(g6068), .A2(g24183), .A3(g25319) );
  NOR2_X1 NOR2_963( .ZN(g26090), .A1(g25518), .A2(g25560) );
  NOR3_X1 NOR3_370( .ZN(g26096), .A1(g6068), .A2(g24183), .A3(g25394) );
  NOR3_X1 NOR3_371( .ZN(g26099), .A1(g6068), .A2(g24183), .A3(g25313) );
  NOR2_X1 NOR2_964( .ZN(g26103), .A1(g25565), .A2(g25626) );
  NOR3_X1 NOR3_372( .ZN(g26107), .A1(g6068), .A2(g24183), .A3(g25383) );
  NOR3_X1 NOR3_373( .ZN(g26110), .A1(g6068), .A2(g24183), .A3(g25305) );
  NOR2_X1 NOR2_965( .ZN(g26113), .A1(g25426), .A2(g22319) );
  NOR3_X1 NOR3_374( .ZN(g26126), .A1(g6068), .A2(g24183), .A3(g25368) );
  NOR3_X1 NOR3_375( .ZN(g26137), .A1(g6068), .A2(g24183), .A3(g25355) );
  NOR2_X1 NOR2_966( .ZN(g26140), .A1(g24183), .A2(g25430) );
  NOR3_X1 NOR3_376( .ZN(g26145), .A1(g6068), .A2(g24183), .A3(g25347) );
  NOR3_X1 NOR3_377( .ZN(g26151), .A1(g6068), .A2(g24183), .A3(g25335) );
  NOR3_X1 NOR3_378( .ZN(g26154), .A1(g6068), .A2(g24183), .A3(g25329) );
  NOR2_X1 NOR2_967( .ZN(g26160), .A1(g25951), .A2(g16162) );
  NOR2_X1 NOR2_968( .ZN(g26168), .A1(g25953), .A2(g16212) );
  NOR2_X1 NOR2_969( .ZN(g26183), .A1(g25957), .A2(g13270) );
  NOR2_X1 NOR2_970( .ZN(g26199), .A1(g25961), .A2(g13291) );
  NOR2_X1 NOR2_971( .ZN(g26217), .A1(g25963), .A2(g13320) );
  NOR2_X1 NOR2_972( .ZN(g26240), .A1(g25968), .A2(g13340) );
  NOR2_X1 NOR2_973( .ZN(g26265), .A1(g25972), .A2(g13360) );
  NOR2_X1 NOR2_974( .ZN(g26272), .A1(g25973), .A2(g16423) );
  NOR2_X1 NOR2_975( .ZN(g26283), .A1(g25954), .A2(g24486) );
  NOR2_X1 NOR2_976( .ZN(g26295), .A1(g25977), .A2(g13385) );
  NOR2_X1 NOR2_977( .ZN(g26304), .A1(g25978), .A2(g16451) );
  NOR2_X1 NOR2_978( .ZN(g26327), .A1(g25958), .A2(g24493) );
  NOR2_X1 NOR2_979( .ZN(g26336), .A1(g25981), .A2(g13481) );
  NOR2_X1 NOR2_980( .ZN(g26374), .A1(g25964), .A2(g24503) );
  NOR2_X1 NOR2_981( .ZN(g26417), .A1(g25969), .A2(g24515) );
  NOR2_X1 NOR2_982( .ZN(g26529), .A1(g25962), .A2(g17001) );
  NOR2_X1 NOR2_983( .ZN(g26530), .A1(g25967), .A2(g17031) );
  NOR2_X1 NOR2_984( .ZN(g26531), .A1(g25974), .A2(g17065) );
  NOR2_X1 NOR2_985( .ZN(g26532), .A1(g25979), .A2(g17100) );
  NOR2_X1 NOR2_986( .ZN(g26534), .A1(g25321), .A2(g8869) );
  NOR2_X1 NOR2_987( .ZN(g26541), .A1(g13755), .A2(g25269) );
  NOR2_X1 NOR2_988( .ZN(g26545), .A1(g13790), .A2(g25277) );
  NOR2_X1 NOR2_989( .ZN(g26547), .A1(g13796), .A2(g25278) );
  NOR2_X1 NOR2_990( .ZN(g26553), .A1(g13816), .A2(g25282) );
  NOR2_X1 NOR2_991( .ZN(g26557), .A1(g13818), .A2(g25286) );
  NOR2_X1 NOR2_992( .ZN(g26559), .A1(g13824), .A2(g25287) );
  NOR2_X1 NOR2_993( .ZN(g26560), .A1(g25281), .A2(g24559) );
  NOR2_X1 NOR2_994( .ZN(g26569), .A1(g13837), .A2(g25290) );
  NOR2_X1 NOR2_995( .ZN(g26573), .A1(g13839), .A2(g25294) );
  NOR2_X1 NOR2_996( .ZN(g26575), .A1(g13845), .A2(g25295) );
  NOR2_X1 NOR2_997( .ZN(g26583), .A1(g25289), .A2(g24569) );
  NOR2_X1 NOR2_998( .ZN(g26592), .A1(g13851), .A2(g25300) );
  NOR2_X1 NOR2_999( .ZN(g26596), .A1(g13853), .A2(g25304) );
  NOR2_X1 NOR2_1000( .ZN(g26607), .A1(g25299), .A2(g24578) );
  NOR2_X1 NOR2_1001( .ZN(g26616), .A1(g13860), .A2(g25310) );
  NOR2_X1 NOR2_1002( .ZN(g26630), .A1(g25309), .A2(g24585) );
  NOR2_X1 NOR2_1003( .ZN(g26655), .A1(g25328), .A2(g17084) );
  NOR2_X1 NOR2_1004( .ZN(g26659), .A1(g25334), .A2(g17116) );
  NOR2_X1 NOR2_1005( .ZN(g26660), .A1(g25208), .A2(g10024) );
  NOR2_X1 NOR2_1006( .ZN(g26661), .A1(g25337), .A2(g17122) );
  NOR2_X1 NOR2_1007( .ZN(g26664), .A1(g25346), .A2(g17138) );
  NOR2_X1 NOR2_1008( .ZN(g26665), .A1(g25348), .A2(g17143) );
  NOR2_X1 NOR2_1009( .ZN(g26666), .A1(g25216), .A2(g10133) );
  NOR2_X1 NOR2_1010( .ZN(g26667), .A1(g25351), .A2(g17149) );
  NOR2_X1 NOR2_1011( .ZN(g26669), .A1(g25360), .A2(g17161) );
  NOR2_X1 NOR2_1012( .ZN(g26670), .A1(g25362), .A2(g17166) );
  NOR2_X1 NOR2_1013( .ZN(g26671), .A1(g25226), .A2(g10238) );
  NOR2_X1 NOR2_1014( .ZN(g26672), .A1(g25365), .A2(g17172) );
  NOR2_X1 NOR2_1015( .ZN(g26675), .A1(g25375), .A2(g17176) );
  NOR2_X1 NOR2_1016( .ZN(g26676), .A1(g25377), .A2(g17181) );
  NOR2_X1 NOR2_1017( .ZN(g26677), .A1(g25238), .A2(g10340) );
  NOR2_X1 NOR2_1018( .ZN(g26776), .A1(g26042), .A2(g10024) );
  NOR2_X1 NOR2_1019( .ZN(g26781), .A1(g26044), .A2(g10133) );
  NOR2_X1 NOR2_1020( .ZN(g26786), .A1(g26049), .A2(g22777) );
  NOR2_X1 NOR2_1021( .ZN(g26789), .A1(g26046), .A2(g10238) );
  NOR2_X1 NOR2_1022( .ZN(g26795), .A1(g26050), .A2(g10340) );
  NOR2_X1 NOR2_1023( .ZN(g26798), .A1(g26055), .A2(g18407) );
  NOR2_X1 NOR2_1024( .ZN(g26799), .A1(g26158), .A2(g25453) );
  NOR2_X1 NOR2_1025( .ZN(g26800), .A1(g26163), .A2(g25457) );
  NOR2_X1 NOR2_1026( .ZN(g26801), .A1(g26171), .A2(g25461) );
  NOR2_X1 NOR2_1027( .ZN(g26802), .A1(g26188), .A2(g25466) );
  NOR2_X1 NOR2_1028( .ZN(g26803), .A1(g15105), .A2(g26213) );
  NOR2_X1 NOR2_1029( .ZN(g26804), .A1(g15172), .A2(g26235) );
  NOR2_X1 NOR2_1030( .ZN(g26805), .A1(g15173), .A2(g26236) );
  NOR2_X1 NOR2_1031( .ZN(g26806), .A1(g15197), .A2(g26244) );
  NOR2_X1 NOR2_1032( .ZN(g26807), .A1(g15245), .A2(g26261) );
  NOR2_X1 NOR2_1033( .ZN(g26808), .A1(g15246), .A2(g26262) );
  NOR2_X1 NOR2_1034( .ZN(g26809), .A1(g15258), .A2(g26270) );
  NOR2_X1 NOR2_1035( .ZN(g26810), .A1(g15259), .A2(g26271) );
  NOR2_X1 NOR2_1036( .ZN(g26811), .A1(g15283), .A2(g26279) );
  NOR2_X1 NOR2_1037( .ZN(g26812), .A1(g15321), .A2(g26291) );
  NOR2_X1 NOR2_1038( .ZN(g26813), .A1(g15337), .A2(g26302) );
  NOR2_X1 NOR2_1039( .ZN(g26814), .A1(g15338), .A2(g26303) );
  NOR2_X1 NOR2_1040( .ZN(g26815), .A1(g15350), .A2(g26311) );
  NOR2_X1 NOR2_1041( .ZN(g26816), .A1(g15351), .A2(g26312) );
  NOR2_X1 NOR2_1042( .ZN(g26817), .A1(g15375), .A2(g26317) );
  NOR2_X1 NOR2_1043( .ZN(g26818), .A1(g15407), .A2(g26335) );
  NOR2_X1 NOR2_1044( .ZN(g26820), .A1(g15423), .A2(g26346) );
  NOR2_X1 NOR2_1045( .ZN(g26821), .A1(g15424), .A2(g26347) );
  NOR2_X1 NOR2_1046( .ZN(g26822), .A1(g15436), .A2(g26352) );
  NOR2_X1 NOR2_1047( .ZN(g26823), .A1(g15437), .A2(g26353) );
  NOR2_X1 NOR2_1048( .ZN(g26824), .A1(g15491), .A2(g26382) );
  NOR2_X1 NOR2_1049( .ZN(g26825), .A1(g15507), .A2(g26390) );
  NOR2_X1 NOR2_1050( .ZN(g26826), .A1(g15508), .A2(g26391) );
  NOR2_X1 NOR2_1051( .ZN(g26827), .A1(g15577), .A2(g26425) );
  NOR2_X1 NOR2_1052( .ZN(g26869), .A1(g26458), .A2(g5642) );
  NOR2_X1 NOR2_1053( .ZN(g26873), .A1(g25483), .A2(g26260) );
  NOR2_X1 NOR2_1054( .ZN(g26877), .A1(g26140), .A2(g22319) );
  NOR2_X1 NOR2_1055( .ZN(g26878), .A1(g26482), .A2(g5680) );
  NOR2_X1 NOR2_1056( .ZN(g26882), .A1(g25514), .A2(g26301) );
  NOR2_X1 NOR2_1057( .ZN(g26885), .A1(g26140), .A2(g22319) );
  NOR2_X1 NOR2_1058( .ZN(g26887), .A1(g26498), .A2(g5732) );
  NOR2_X1 NOR2_1059( .ZN(g26891), .A1(g25561), .A2(g26345) );
  NOR2_X1 NOR2_1060( .ZN(g26897), .A1(g26513), .A2(g5790) );
  NOR2_X1 NOR2_1061( .ZN(g26901), .A1(g25627), .A2(g26389) );
  NOR2_X1 NOR2_1062( .ZN(g26905), .A1(g26096), .A2(g22319) );
  NOR2_X1 NOR2_1063( .ZN(g26914), .A1(g26107), .A2(g22319) );
  NOR2_X1 NOR2_1064( .ZN(g26988), .A1(g24893), .A2(g26023) );
  NOR2_X1 NOR2_1065( .ZN(g26989), .A1(g26663), .A2(g21913) );
  NOR2_X1 NOR2_1066( .ZN(g27011), .A1(g24916), .A2(g26026) );
  NOR2_X1 NOR2_1067( .ZN(g27012), .A1(g26668), .A2(g21931) );
  NOR2_X1 NOR2_1068( .ZN(g27037), .A1(g24933), .A2(g26028) );
  NOR2_X2 NOR2_1069( .ZN(g27038), .A1(g26674), .A2(g20640) );
  NOR2_X2 NOR2_1070( .ZN(g27051), .A1(g4456), .A2(g26081) );
  NOR2_X1 NOR2_1071( .ZN(g27065), .A1(g24945), .A2(g26029) );
  NOR2_X1 NOR2_1072( .ZN(g27066), .A1(g26024), .A2(g20665) );
  NOR2_X1 NOR2_1073( .ZN(g27078), .A1(g4632), .A2(g26084) );
  NOR2_X1 NOR2_1074( .ZN(g27094), .A1(g4809), .A2(g26090) );
  NOR2_X1 NOR2_1075( .ZN(g27106), .A1(g4985), .A2(g26103) );
  NOR2_X1 NOR2_1076( .ZN(g27120), .A1(g26560), .A2(g17001) );
  NOR2_X1 NOR2_1077( .ZN(g27123), .A1(g26583), .A2(g17031) );
  NOR2_X1 NOR2_1078( .ZN(g27129), .A1(g26607), .A2(g17065) );
  NOR2_X1 NOR2_1079( .ZN(g27131), .A1(g26630), .A2(g17100) );
  NOR2_X1 NOR2_1080( .ZN(g27144), .A1(g23451), .A2(g26052) );
  NOR2_X1 NOR2_1081( .ZN(g27147), .A1(g23458), .A2(g26054) );
  NOR2_X1 NOR2_1082( .ZN(g27149), .A1(g23462), .A2(g26060) );
  NOR2_X1 NOR2_1083( .ZN(g27152), .A1(g23467), .A2(g26062) );
  NOR2_X1 NOR2_1084( .ZN(g27157), .A1(g23471), .A2(g26067) );
  NOR2_X1 NOR2_1085( .ZN(g27160), .A1(g23476), .A2(g26069) );
  NOR2_X1 NOR2_1086( .ZN(g27165), .A1(g23484), .A2(g26074) );
  NOR2_X1 NOR2_1087( .ZN(g27174), .A1(g23494), .A2(g26080) );
  NOR2_X1 NOR2_1088( .ZN(g27175), .A1(g26075), .A2(g25342) );
  NOR2_X1 NOR2_1089( .ZN(g27179), .A1(g26082), .A2(g25356) );
  NOR2_X1 NOR2_1090( .ZN(g27184), .A1(g26085), .A2(g25371) );
  NOR2_X1 NOR2_1091( .ZN(g27188), .A1(g26091), .A2(g25388) );
  NOR2_X1 NOR2_1092( .ZN(g27243), .A1(g26802), .A2(g10340) );
  NOR2_X1 NOR2_1093( .ZN(g27250), .A1(g26955), .A2(g26166) );
  NOR2_X1 NOR2_1094( .ZN(g27251), .A1(g26958), .A2(g26186) );
  NOR2_X1 NOR2_1095( .ZN(g27252), .A1(g26963), .A2(g26207) );
  NOR2_X1 NOR2_1096( .ZN(g27253), .A1(g26965), .A2(g26212) );
  NOR2_X1 NOR2_1097( .ZN(g27254), .A1(g26968), .A2(g26231) );
  NOR2_X1 NOR2_1098( .ZN(g27255), .A1(g26969), .A2(g26233) );
  NOR2_X1 NOR2_1099( .ZN(g27256), .A1(g26970), .A2(g26234) );
  NOR2_X1 NOR2_1100( .ZN(g27257), .A1(g26971), .A2(g26243) );
  NOR2_X1 NOR2_1101( .ZN(g27258), .A1(g26977), .A2(g26257) );
  NOR2_X1 NOR2_1102( .ZN(g27259), .A1(g26978), .A2(g26258) );
  NOR2_X1 NOR2_1103( .ZN(g27260), .A1(g26979), .A2(g26259) );
  NOR2_X1 NOR2_1104( .ZN(g27261), .A1(g26980), .A2(g26263) );
  NOR2_X1 NOR2_1105( .ZN(g27262), .A1(g26981), .A2(g26268) );
  NOR2_X1 NOR2_1106( .ZN(g27263), .A1(g26982), .A2(g26269) );
  NOR2_X1 NOR2_1107( .ZN(g27264), .A1(g26984), .A2(g26278) );
  NOR2_X1 NOR2_1108( .ZN(g27265), .A1(g26993), .A2(g26288) );
  NOR2_X1 NOR2_1109( .ZN(g27266), .A1(g26994), .A2(g26289) );
  NOR2_X1 NOR2_1110( .ZN(g27267), .A1(g26995), .A2(g26290) );
  NOR2_X1 NOR2_1111( .ZN(g27268), .A1(g26996), .A2(g26292) );
  NOR2_X1 NOR2_1112( .ZN(g27269), .A1(g26997), .A2(g26293) );
  NOR2_X1 NOR2_1113( .ZN(g27270), .A1(g26998), .A2(g26298) );
  NOR2_X1 NOR2_1114( .ZN(g27271), .A1(g26999), .A2(g26299) );
  NOR2_X1 NOR2_1115( .ZN(g27272), .A1(g27000), .A2(g26300) );
  NOR2_X1 NOR2_1116( .ZN(g27273), .A1(g27001), .A2(g26307) );
  NOR2_X1 NOR2_1117( .ZN(g27274), .A1(g27002), .A2(g26309) );
  NOR2_X1 NOR2_1118( .ZN(g27275), .A1(g27003), .A2(g26310) );
  NOR2_X1 NOR2_1119( .ZN(g27276), .A1(g27004), .A2(g26316) );
  NOR2_X1 NOR2_1120( .ZN(g27277), .A1(g27005), .A2(g26318) );
  NOR2_X1 NOR2_1121( .ZN(g27278), .A1(g27006), .A2(g26319) );
  NOR2_X1 NOR2_1122( .ZN(g27279), .A1(g27007), .A2(g26324) );
  NOR2_X1 NOR2_1123( .ZN(g27280), .A1(g27008), .A2(g26325) );
  NOR2_X1 NOR2_1124( .ZN(g27281), .A1(g27009), .A2(g26326) );
  NOR2_X1 NOR2_1125( .ZN(g27282), .A1(g27016), .A2(g26332) );
  NOR2_X1 NOR2_1126( .ZN(g27283), .A1(g27017), .A2(g26333) );
  NOR2_X1 NOR2_1127( .ZN(g27284), .A1(g27018), .A2(g26334) );
  NOR2_X1 NOR2_1128( .ZN(g27285), .A1(g27019), .A2(g26339) );
  NOR2_X1 NOR2_1129( .ZN(g27286), .A1(g27020), .A2(g26340) );
  NOR2_X1 NOR2_1130( .ZN(g27287), .A1(g27021), .A2(g26342) );
  NOR2_X1 NOR2_1131( .ZN(g27288), .A1(g27022), .A2(g26343) );
  NOR2_X1 NOR2_1132( .ZN(g27289), .A1(g27023), .A2(g26344) );
  NOR2_X1 NOR2_1133( .ZN(g27290), .A1(g27024), .A2(g26348) );
  NOR2_X1 NOR2_1134( .ZN(g27291), .A1(g27025), .A2(g26350) );
  NOR2_X1 NOR2_1135( .ZN(g27292), .A1(g27026), .A2(g26351) );
  NOR2_X1 NOR2_1136( .ZN(g27293), .A1(g27027), .A2(g26357) );
  NOR2_X1 NOR2_1137( .ZN(g27294), .A1(g27028), .A2(g26361) );
  NOR2_X1 NOR2_1138( .ZN(g27295), .A1(g27029), .A2(g26362) );
  NOR2_X1 NOR2_1139( .ZN(g27296), .A1(g27030), .A2(g26363) );
  NOR2_X1 NOR2_1140( .ZN(g27297), .A1(g27031), .A2(g26365) );
  NOR2_X1 NOR2_1141( .ZN(g27298), .A1(g27032), .A2(g26366) );
  NOR2_X1 NOR2_1142( .ZN(g27299), .A1(g27033), .A2(g26371) );
  NOR2_X1 NOR2_1143( .ZN(g27300), .A1(g27034), .A2(g26372) );
  NOR2_X1 NOR2_1144( .ZN(g27301), .A1(g27035), .A2(g26373) );
  NOR2_X1 NOR2_1145( .ZN(g27302), .A1(g27042), .A2(g26379) );
  NOR2_X1 NOR2_1146( .ZN(g27303), .A1(g27043), .A2(g26380) );
  NOR2_X1 NOR2_1147( .ZN(g27304), .A1(g27044), .A2(g26381) );
  NOR2_X1 NOR2_1148( .ZN(g27305), .A1(g27045), .A2(g26383) );
  NOR2_X1 NOR2_1149( .ZN(g27306), .A1(g27046), .A2(g26384) );
  NOR2_X1 NOR2_1150( .ZN(g27307), .A1(g27047), .A2(g26386) );
  NOR2_X1 NOR2_1151( .ZN(g27308), .A1(g27048), .A2(g26387) );
  NOR2_X1 NOR2_1152( .ZN(g27309), .A1(g27049), .A2(g26388) );
  NOR2_X1 NOR2_1153( .ZN(g27310), .A1(g27050), .A2(g26392) );
  NOR2_X1 NOR2_1154( .ZN(g27311), .A1(g27053), .A2(g26396) );
  NOR2_X1 NOR2_1155( .ZN(g27312), .A1(g27054), .A2(g26397) );
  NOR2_X1 NOR2_1156( .ZN(g27313), .A1(g27055), .A2(g26400) );
  NOR2_X1 NOR2_1157( .ZN(g27314), .A1(g27056), .A2(g26404) );
  NOR2_X1 NOR2_1158( .ZN(g27315), .A1(g27057), .A2(g26405) );
  NOR2_X1 NOR2_1159( .ZN(g27316), .A1(g27058), .A2(g26406) );
  NOR2_X1 NOR2_1160( .ZN(g27317), .A1(g27059), .A2(g26408) );
  NOR2_X1 NOR2_1161( .ZN(g27318), .A1(g27060), .A2(g26409) );
  NOR2_X1 NOR2_1162( .ZN(g27319), .A1(g27061), .A2(g26414) );
  NOR2_X1 NOR2_1163( .ZN(g27320), .A1(g27062), .A2(g26415) );
  NOR2_X1 NOR2_1164( .ZN(g27321), .A1(g27063), .A2(g26416) );
  NOR2_X1 NOR2_1165( .ZN(g27322), .A1(g27070), .A2(g26422) );
  NOR2_X1 NOR2_1166( .ZN(g27323), .A1(g27071), .A2(g26423) );
  NOR2_X1 NOR2_1167( .ZN(g27324), .A1(g27072), .A2(g26424) );
  NOR2_X1 NOR2_1168( .ZN(g27325), .A1(g27073), .A2(g26426) );
  NOR2_X1 NOR2_1169( .ZN(g27326), .A1(g27074), .A2(g26427) );
  NOR2_X1 NOR2_1170( .ZN(g27327), .A1(g27077), .A2(g26432) );
  NOR2_X1 NOR2_1171( .ZN(g27328), .A1(g27080), .A2(g26437) );
  NOR2_X1 NOR2_1172( .ZN(g27329), .A1(g27081), .A2(g26438) );
  NOR2_X1 NOR2_1173( .ZN(g27330), .A1(g27082), .A2(g26441) );
  NOR2_X1 NOR2_1174( .ZN(g27331), .A1(g27083), .A2(g26445) );
  NOR2_X1 NOR2_1175( .ZN(g27332), .A1(g27084), .A2(g26446) );
  NOR2_X1 NOR2_1176( .ZN(g27333), .A1(g27085), .A2(g26447) );
  NOR2_X1 NOR2_1177( .ZN(g27334), .A1(g27086), .A2(g26449) );
  NOR2_X1 NOR2_1178( .ZN(g27335), .A1(g27087), .A2(g26450) );
  NOR2_X1 NOR2_1179( .ZN(g27336), .A1(g27088), .A2(g26455) );
  NOR2_X1 NOR2_1180( .ZN(g27337), .A1(g27089), .A2(g26456) );
  NOR2_X1 NOR2_1181( .ZN(g27338), .A1(g27090), .A2(g26457) );
  NOR2_X1 NOR2_1182( .ZN(g27339), .A1(g27093), .A2(g26464) );
  NOR2_X1 NOR2_1183( .ZN(g27340), .A1(g27096), .A2(g26469) );
  NOR2_X1 NOR2_1184( .ZN(g27341), .A1(g27097), .A2(g26470) );
  NOR2_X1 NOR2_1185( .ZN(g27342), .A1(g27098), .A2(g26473) );
  NOR2_X1 NOR2_1186( .ZN(g27343), .A1(g27099), .A2(g26477) );
  NOR2_X1 NOR2_1187( .ZN(g27344), .A1(g27100), .A2(g26478) );
  NOR2_X1 NOR2_1188( .ZN(g27345), .A1(g27101), .A2(g26479) );
  NOR2_X1 NOR2_1189( .ZN(g27346), .A1(g27105), .A2(g26488) );
  NOR2_X1 NOR2_1190( .ZN(g27347), .A1(g27108), .A2(g26493) );
  NOR2_X1 NOR2_1191( .ZN(g27348), .A1(g27109), .A2(g26494) );
  NOR2_X1 NOR2_1192( .ZN(g27354), .A1(g27112), .A2(g26504) );
  NOR2_X1 NOR2_1193( .ZN(g27414), .A1(g26770), .A2(g25187) );
  NOR3_X1 NOR3_379( .ZN(g27415), .A1(g23104), .A2(g27181), .A3(g25128) );
  NOR2_X1 NOR2_1194( .ZN(g27435), .A1(g26777), .A2(g25193) );
  NOR3_X1 NOR3_380( .ZN(g27436), .A1(g23118), .A2(g27187), .A3(g24427) );
  NOR2_X1 NOR2_1195( .ZN(g27450), .A1(g26902), .A2(g24613) );
  NOR2_X1 NOR2_1196( .ZN(g27454), .A1(g26783), .A2(g25196) );
  NOR3_X1 NOR3_381( .ZN(g27455), .A1(g23127), .A2(g26758), .A3(g24431) );
  NOR2_X1 NOR2_1197( .ZN(g27462), .A1(g26892), .A2(g24622) );
  NOR2_X1 NOR2_1198( .ZN(g27464), .A1(g27178), .A2(g25975) );
  NOR2_X1 NOR2_1199( .ZN(g27466), .A1(g26915), .A2(g24624) );
  NOR2_X1 NOR2_1200( .ZN(g27470), .A1(g26790), .A2(g25198) );
  NOR3_X1 NOR3_382( .ZN(g27471), .A1(g23138), .A2(g26764), .A3(g24435) );
  NOR2_X1 NOR2_1201( .ZN(g27478), .A1(g26754), .A2(g24432) );
  NOR2_X1 NOR2_1202( .ZN(g27481), .A1(g27182), .A2(g25980) );
  NOR2_X1 NOR2_1203( .ZN(g27482), .A1(g26906), .A2(g24637) );
  NOR2_X1 NOR2_1204( .ZN(g27485), .A1(g26928), .A2(g24638) );
  NOR3_X1 NOR3_383( .ZN(g27492), .A1(g24958), .A2(g24633), .A3(g26771) );
  NOR2_X1 NOR2_1205( .ZN(g27496), .A1(g27185), .A2(g25178) );
  NOR2_X1 NOR2_1206( .ZN(g27501), .A1(g26763), .A2(g24436) );
  NOR2_X1 NOR2_1207( .ZN(g27504), .A1(g26918), .A2(g24656) );
  NOR2_X1 NOR2_1208( .ZN(g27507), .A1(g26941), .A2(g24657) );
  NOR3_X1 NOR3_384( .ZN(g27513), .A1(g24969), .A2(g24653), .A3(g26778) );
  NOR2_X1 NOR2_1209( .ZN(g27521), .A1(g26766), .A2(g24439) );
  NOR2_X1 NOR2_1210( .ZN(g27524), .A1(g26931), .A2(g24675) );
  NOR2_X1 NOR2_1211( .ZN(g27527), .A1(g26759), .A2(g19087) );
  NOR2_X1 NOR2_1212( .ZN(g27529), .A1(g4456), .A2(g26873) );
  NOR2_X1 NOR2_1213( .ZN(g27531), .A1(g26760), .A2(g25181) );
  NOR2_X1 NOR2_1214( .ZN(g27532), .A1(g26761), .A2(g25182) );
  NOR3_X1 NOR3_385( .ZN(g27538), .A1(g24982), .A2(g24672), .A3(g26784) );
  NOR2_X1 NOR2_1215( .ZN(g27546), .A1(g26769), .A2(g24441) );
  NOR2_X1 NOR2_1216( .ZN(g27549), .A1(g26765), .A2(g19093) );
  NOR2_X1 NOR2_1217( .ZN(g27551), .A1(g4632), .A2(g26882) );
  NOR3_X1 NOR3_386( .ZN(g27558), .A1(g24993), .A2(g24691), .A3(g26791) );
  NOR2_X1 NOR2_1218( .ZN(g27563), .A1(g26922), .A2(g24708) );
  NOR2_X1 NOR2_1219( .ZN(g27564), .A1(g26767), .A2(g25184) );
  NOR2_X1 NOR2_1220( .ZN(g27565), .A1(g26768), .A2(g19100) );
  NOR2_X1 NOR2_1221( .ZN(g27567), .A1(g4809), .A2(g26891) );
  NOR2_X1 NOR2_1222( .ZN(g27572), .A1(g26911), .A2(g24717) );
  NOR2_X1 NOR2_1223( .ZN(g27573), .A1(g26773), .A2(g25188) );
  NOR2_X1 NOR2_1224( .ZN(g27574), .A1(g26935), .A2(g24720) );
  NOR2_X1 NOR2_1225( .ZN(g27575), .A1(g26774), .A2(g19107) );
  NOR2_X1 NOR2_1226( .ZN(g27577), .A1(g4985), .A2(g26901) );
  NOR2_X1 NOR2_1227( .ZN(g27579), .A1(g26775), .A2(g25192) );
  NOR2_X1 NOR2_1228( .ZN(g27581), .A1(g26925), .A2(g24728) );
  NOR2_X1 NOR2_1229( .ZN(g27582), .A1(g26944), .A2(g24731) );
  NOR2_X1 NOR2_1230( .ZN(g27584), .A1(g26938), .A2(g24736) );
  NOR2_X1 NOR2_1231( .ZN(g27585), .A1(g26950), .A2(g24739) );
  NOR2_X1 NOR2_1232( .ZN(g27588), .A1(g26947), .A2(g24742) );
  NOR2_X1 NOR2_1233( .ZN(g27594), .A1(g27175), .A2(g17001) );
  NOR2_X1 NOR2_1234( .ZN(g27603), .A1(g27179), .A2(g17031) );
  NOR2_X1 NOR2_1235( .ZN(g27612), .A1(g27184), .A2(g17065) );
  NOR2_X1 NOR2_1236( .ZN(g27621), .A1(g27188), .A2(g17100) );
  NOR2_X1 NOR2_1237( .ZN(g27629), .A1(g26829), .A2(g26051) );
  NOR2_X1 NOR2_1238( .ZN(g27631), .A1(g26833), .A2(g26053) );
  NOR2_X1 NOR2_1239( .ZN(g27655), .A1(g26842), .A2(g26061) );
  NOR2_X1 NOR2_1240( .ZN(g27658), .A1(g26851), .A2(g26068) );
  NOR2_X1 NOR2_1241( .ZN(g27672), .A1(g26799), .A2(g10024) );
  NOR2_X1 NOR2_1242( .ZN(g27678), .A1(g26800), .A2(g10133) );
  NOR2_X1 NOR2_1243( .ZN(g27682), .A1(g26801), .A2(g10238) );
  NOR2_X1 NOR2_1244( .ZN(g27718), .A1(g27251), .A2(g10133) );
  NOR2_X1 NOR2_1245( .ZN(g27722), .A1(g27252), .A2(g10238) );
  NOR2_X1 NOR2_1246( .ZN(g27724), .A1(g27254), .A2(g10340) );
  NOR2_X1 NOR2_1247( .ZN(g27735), .A1(g27394), .A2(g26961) );
  NOR2_X1 NOR2_1248( .ZN(g27736), .A1(g27396), .A2(g26962) );
  NOR2_X1 NOR2_1249( .ZN(g27741), .A1(g27407), .A2(g26966) );
  NOR2_X1 NOR2_1250( .ZN(g27742), .A1(g27409), .A2(g26967) );
  NOR2_X1 NOR2_1251( .ZN(g27746), .A1(g27425), .A2(g26972) );
  NOR2_X1 NOR2_1252( .ZN(g27747), .A1(g27427), .A2(g26973) );
  NOR2_X1 NOR2_1253( .ZN(g27754), .A1(g27446), .A2(g26985) );
  NOR2_X1 NOR2_1254( .ZN(g27755), .A1(g27448), .A2(g26986) );
  NOR2_X1 NOR2_1255( .ZN(g27759), .A1(g27495), .A2(g27052) );
  NOR2_X1 NOR2_1256( .ZN(g27760), .A1(g27509), .A2(g27076) );
  NOR2_X1 NOR2_1257( .ZN(g27761), .A1(g27516), .A2(g27079) );
  NOR2_X1 NOR2_1258( .ZN(g27762), .A1(g27530), .A2(g27091) );
  NOR2_X1 NOR2_1259( .ZN(g27763), .A1(g27534), .A2(g27092) );
  NOR2_X1 NOR2_1260( .ZN(g27764), .A1(g27541), .A2(g27095) );
  NOR2_X1 NOR2_1261( .ZN(g27765), .A1(g27552), .A2(g27103) );
  NOR2_X1 NOR2_1262( .ZN(g27766), .A1(g27554), .A2(g27104) );
  NOR2_X1 NOR2_1263( .ZN(g27767), .A1(g27561), .A2(g27107) );
  NOR2_X1 NOR2_1264( .ZN(g27768), .A1(g27568), .A2(g27110) );
  NOR2_X1 NOR2_1265( .ZN(g27769), .A1(g27570), .A2(g27111) );
  NOR2_X1 NOR2_1266( .ZN(g27771), .A1(g27578), .A2(g27115) );
  NOR2_X1 NOR2_1267( .ZN(g27798), .A1(g27632), .A2(g1223) );
  NOR3_X1 NOR3_387( .ZN(g27802), .A1(g6087), .A2(g27632), .A3(g25330) );
  NOR2_X1 NOR2_1268( .ZN(g27810), .A1(g27632), .A2(g1215) );
  NOR3_X1 NOR3_388( .ZN(g27811), .A1(g6087), .A2(g27632), .A3(g25404) );
  NOR3_X1 NOR3_389( .ZN(g27814), .A1(g6087), .A2(g27632), .A3(g25322) );
  NOR2_X1 NOR2_1269( .ZN(g27823), .A1(g27632), .A2(g1216) );
  NOR3_X1 NOR3_390( .ZN(g27824), .A1(g6087), .A2(g27632), .A3(g25399) );
  NOR3_X1 NOR3_391( .ZN(g27827), .A1(g6087), .A2(g27632), .A3(g25314) );
  NOR2_X1 NOR2_1270( .ZN(g27834), .A1(g27478), .A2(g14630) );
  NOR2_X1 NOR2_1271( .ZN(g27842), .A1(g27632), .A2(g1217) );
  NOR2_X1 NOR2_1272( .ZN(g27850), .A1(g27501), .A2(g14650) );
  NOR2_X1 NOR2_1273( .ZN(g27854), .A1(g27632), .A2(g1218) );
  NOR3_X1 NOR3_392( .ZN(g27855), .A1(g6087), .A2(g27632), .A3(g25385) );
  NOR2_X1 NOR2_1274( .ZN(g27864), .A1(g27632), .A2(g1219) );
  NOR3_X1 NOR3_393( .ZN(g27865), .A1(g6087), .A2(g27632), .A3(g25370) );
  NOR2_X1 NOR2_1275( .ZN(g27868), .A1(g23742), .A2(g27632) );
  NOR2_X1 NOR2_1276( .ZN(g27869), .A1(g27632), .A2(g25437) );
  NOR2_X1 NOR2_1277( .ZN(g27875), .A1(g27521), .A2(g14677) );
  NOR2_X1 NOR2_1278( .ZN(g27882), .A1(g27632), .A2(g1220) );
  NOR3_X1 NOR3_394( .ZN(g27883), .A1(g6087), .A2(g27632), .A3(g25361) );
  NOR2_X1 NOR2_1279( .ZN(g27886), .A1(g27632), .A2(g24627) );
  NOR2_X1 NOR2_1280( .ZN(g27892), .A1(g27546), .A2(g14711) );
  NOR2_X1 NOR2_1281( .ZN(g27896), .A1(g27632), .A2(g1222) );
  NOR3_X1 NOR3_395( .ZN(g27897), .A1(g6087), .A2(g27632), .A3(g25349) );
  NOR3_X1 NOR3_396( .ZN(g27900), .A1(g6087), .A2(g27632), .A3(g25338) );
  NOR2_X1 NOR2_1282( .ZN(g27906), .A1(g16127), .A2(g27656) );
  NOR2_X1 NOR2_1283( .ZN(g27911), .A1(g16170), .A2(g27657) );
  NOR2_X1 NOR2_1284( .ZN(g27916), .A1(g16219), .A2(g27659) );
  NOR2_X1 NOR2_1285( .ZN(g27917), .A1(g16220), .A2(g27660) );
  NOR2_X1 NOR2_1286( .ZN(g27925), .A1(g16276), .A2(g27661) );
  NOR2_X1 NOR2_1287( .ZN(g27937), .A1(g16321), .A2(g27666) );
  NOR2_X1 NOR2_1288( .ZN(g27950), .A1(g16367), .A2(g27673) );
  NOR2_X1 NOR2_1289( .ZN(g27962), .A1(g16394), .A2(g27679) );
  NOR2_X1 NOR2_1290( .ZN(g27964), .A1(g16400), .A2(g27680) );
  NOR2_X1 NOR2_1291( .ZN(g27980), .A1(g16428), .A2(g27681) );
  NOR2_X1 NOR2_1292( .ZN(g27997), .A1(g16456), .A2(g27242) );
  NOR2_X1 NOR2_1293( .ZN(g28002), .A1(g26032), .A2(g27246) );
  NOR2_X1 NOR2_1294( .ZN(g28029), .A1(g26033), .A2(g27247) );
  NOR2_X1 NOR2_1295( .ZN(g28059), .A1(g26034), .A2(g27248) );
  NOR2_X1 NOR2_1296( .ZN(g28088), .A1(g26036), .A2(g27249) );
  NOR2_X1 NOR2_1297( .ZN(g28145), .A1(g27629), .A2(g17001) );
  NOR2_X1 NOR2_1298( .ZN(g28146), .A1(g27631), .A2(g17031) );
  NOR2_X1 NOR2_1299( .ZN(g28147), .A1(g27655), .A2(g17065) );
  NOR2_X1 NOR2_1300( .ZN(g28148), .A1(g27658), .A2(g17100) );
  NOR2_X1 NOR2_1301( .ZN(g28157), .A1(g13902), .A2(g27370) );
  NOR2_X1 NOR2_1302( .ZN(g28185), .A1(g27356), .A2(g26845) );
  NOR2_X1 NOR2_1303( .ZN(g28189), .A1(g27359), .A2(g26853) );
  NOR2_X1 NOR2_1304( .ZN(g28191), .A1(g27365), .A2(g26860) );
  NOR2_X1 NOR2_1305( .ZN(g28192), .A1(g27372), .A2(g26866) );
  NOR2_X1 NOR2_1306( .ZN(g28199), .A1(g27250), .A2(g10024) );
  NOR2_X1 NOR2_1307( .ZN(g28321), .A1(g27742), .A2(g10133) );
  NOR2_X1 NOR2_1308( .ZN(g28325), .A1(g27747), .A2(g10238) );
  NOR2_X1 NOR2_1309( .ZN(g28328), .A1(g27755), .A2(g10340) );
  NOR2_X1 NOR2_1310( .ZN(g28342), .A1(g15460), .A2(g28008) );
  NOR2_X1 NOR2_1311( .ZN(g28344), .A1(g15526), .A2(g28027) );
  NOR2_X1 NOR2_1312( .ZN(g28345), .A1(g15527), .A2(g28028) );
  NOR2_X1 NOR2_1313( .ZN(g28346), .A1(g15546), .A2(g28035) );
  NOR2_X1 NOR2_1314( .ZN(g28348), .A1(g15594), .A2(g28050) );
  NOR2_X1 NOR2_1315( .ZN(g28349), .A1(g15595), .A2(g28051) );
  NOR2_X1 NOR2_1316( .ZN(g28350), .A1(g15604), .A2(g28057) );
  NOR2_X1 NOR2_1317( .ZN(g28351), .A1(g15605), .A2(g28058) );
  NOR2_X1 NOR2_1318( .ZN(g28352), .A1(g15624), .A2(g28065) );
  NOR2_X1 NOR2_1319( .ZN(g28353), .A1(g15666), .A2(g28073) );
  NOR2_X1 NOR2_1320( .ZN(g28354), .A1(g15670), .A2(g28079) );
  NOR2_X1 NOR2_1321( .ZN(g28355), .A1(g15671), .A2(g28080) );
  NOR2_X1 NOR2_1322( .ZN(g28356), .A1(g15680), .A2(g28086) );
  NOR2_X1 NOR2_1323( .ZN(g28357), .A1(g15681), .A2(g28087) );
  NOR2_X1 NOR2_1324( .ZN(g28358), .A1(g15700), .A2(g28094) );
  NOR2_X1 NOR2_1325( .ZN(g28360), .A1(g15725), .A2(g28098) );
  NOR2_X1 NOR2_1326( .ZN(g28361), .A1(g15729), .A2(g28104) );
  NOR2_X1 NOR2_1327( .ZN(g28362), .A1(g15730), .A2(g28105) );
  NOR2_X1 NOR2_1328( .ZN(g28363), .A1(g15739), .A2(g28111) );
  NOR2_X1 NOR2_1329( .ZN(g28364), .A1(g15740), .A2(g28112) );
  NOR2_X1 NOR2_1330( .ZN(g28366), .A1(g15765), .A2(g28116) );
  NOR2_X1 NOR2_1331( .ZN(g28367), .A1(g15769), .A2(g28122) );
  NOR2_X1 NOR2_1332( .ZN(g28368), .A1(g15770), .A2(g28123) );
  NOR2_X1 NOR2_1333( .ZN(g28371), .A1(g15793), .A2(g28127) );
  NOR2_X1 NOR2_1334( .ZN(g28392), .A1(g27886), .A2(g22344) );
  NOR2_X1 NOR2_1335( .ZN(g28394), .A1(g27869), .A2(g22344) );
  NOR2_X1 NOR2_1336( .ZN(g28397), .A1(g27869), .A2(g22344) );
  NOR2_X1 NOR2_1337( .ZN(g28400), .A1(g27886), .A2(g22344) );
  NOR2_X1 NOR2_1338( .ZN(g28403), .A1(g27811), .A2(g22344) );
  NOR2_X1 NOR2_1339( .ZN(g28406), .A1(g27824), .A2(g22344) );
  NOR2_X1 NOR2_1340( .ZN(g28409), .A1(g24676), .A2(g27801) );
  NOR2_X1 NOR2_1341( .ZN(g28410), .A1(g27748), .A2(g22344) );
  NOR2_X1 NOR2_1342( .ZN(g28413), .A1(g24695), .A2(g27809) );
  NOR2_X1 NOR2_1343( .ZN(g28414), .A1(g27748), .A2(g22344) );
  NOR2_X1 NOR2_1344( .ZN(g28417), .A1(g24712), .A2(g27830) );
  NOR2_X1 NOR2_1345( .ZN(g28418), .A1(g24723), .A2(g27846) );
  NOR2_X1 NOR2_1346( .ZN(g28420), .A1(g16031), .A2(g28171) );
  NOR2_X1 NOR2_1347( .ZN(g28421), .A1(g16068), .A2(g28176) );
  NOR2_X1 NOR2_1348( .ZN(g28425), .A1(g16133), .A2(g28188) );
  NOR2_X1 NOR2_1349( .ZN(g28449), .A1(g27727), .A2(g26780) );
  NOR2_X2 NOR2_1350( .ZN(g28461), .A1(g27729), .A2(g26787) );
  NOR2_X2 NOR2_1351( .ZN(g28470), .A1(g27671), .A2(g28193) );
  NOR2_X1 NOR2_1352( .ZN(g28473), .A1(g27730), .A2(g26794) );
  NOR2_X1 NOR2_1353( .ZN(g28482), .A1(g27731), .A2(g26797) );
  NOR2_X1 NOR2_1354( .ZN(g28488), .A1(g26755), .A2(g27719) );
  NOR2_X1 NOR2_1355( .ZN(g28489), .A1(g26756), .A2(g27720) );
  NOR2_X1 NOR2_1356( .ZN(g28490), .A1(g27240), .A2(g27721) );
  NOR2_X1 NOR2_1357( .ZN(g28495), .A1(g27244), .A2(g27723) );
  NOR2_X1 NOR2_1358( .ZN(g28499), .A1(g26027), .A2(g27725) );
  NOR2_X1 NOR2_1359( .ZN(g28523), .A1(g26035), .A2(g27732) );
  NOR2_X1 NOR2_1360( .ZN(g28525), .A1(g27245), .A2(g27726) );
  NOR2_X1 NOR2_1361( .ZN(g28528), .A1(g26030), .A2(g27728) );
  NOR2_X1 NOR2_1362( .ZN(g28551), .A1(g26038), .A2(g27733) );
  NOR2_X1 NOR2_1363( .ZN(g28578), .A1(g26039), .A2(g27734) );
  NOR2_X1 NOR2_1364( .ZN(g28606), .A1(g26040), .A2(g27737) );
  NOR2_X1 NOR2_1365( .ZN(g28634), .A1(g28185), .A2(g17001) );
  NOR2_X1 NOR2_1366( .ZN(g28635), .A1(g28189), .A2(g17031) );
  NOR2_X1 NOR2_1367( .ZN(g28636), .A1(g28191), .A2(g17065) );
  NOR2_X1 NOR2_1368( .ZN(g28637), .A1(g28192), .A2(g17100) );
  NOR2_X1 NOR2_1369( .ZN(g28654), .A1(g27770), .A2(g27355) );
  NOR2_X1 NOR2_1370( .ZN(g28656), .A1(g27772), .A2(g27358) );
  NOR2_X1 NOR2_1371( .ZN(g28658), .A1(g27773), .A2(g27364) );
  NOR2_X1 NOR2_1372( .ZN(g28661), .A1(g27775), .A2(g27371) );
  NOR2_X1 NOR2_1373( .ZN(g28668), .A1(g27736), .A2(g10024) );
  NOR2_X1 NOR2_1374( .ZN(g28728), .A1(g28422), .A2(g27904) );
  NOR2_X1 NOR2_1375( .ZN(g28731), .A1(g28423), .A2(g27908) );
  NOR2_X1 NOR2_1376( .ZN(g28732), .A1(g14894), .A2(g28426) );
  NOR2_X1 NOR2_1377( .ZN(g28733), .A1(g28424), .A2(g27909) );
  NOR2_X1 NOR2_1378( .ZN(g28735), .A1(g14957), .A2(g28430) );
  NOR2_X1 NOR2_1379( .ZN(g28736), .A1(g28427), .A2(g27913) );
  NOR2_X1 NOR2_1380( .ZN(g28737), .A1(g28428), .A2(g27914) );
  NOR2_X1 NOR2_1381( .ZN(g28738), .A1(g14975), .A2(g28433) );
  NOR2_X1 NOR2_1382( .ZN(g28739), .A1(g28429), .A2(g27915) );
  NOR2_X1 NOR2_1383( .ZN(g28744), .A1(g15030), .A2(g28439) );
  NOR2_X1 NOR2_1384( .ZN(g28745), .A1(g28431), .A2(g27922) );
  NOR2_X1 NOR2_1385( .ZN(g28746), .A1(g15046), .A2(g28441) );
  NOR2_X1 NOR2_1386( .ZN(g28747), .A1(g28434), .A2(g27923) );
  NOR2_X1 NOR2_1387( .ZN(g28748), .A1(g28435), .A2(g27924) );
  NOR2_X1 NOR2_1388( .ZN(g28749), .A1(g15064), .A2(g28444) );
  NOR2_X1 NOR2_1389( .ZN(g28750), .A1(g28436), .A2(g27926) );
  NOR2_X1 NOR2_1390( .ZN(g28754), .A1(g28440), .A2(g27931) );
  NOR2_X1 NOR2_1391( .ZN(g28758), .A1(g15126), .A2(g28451) );
  NOR2_X1 NOR2_1392( .ZN(g28759), .A1(g28442), .A2(g27935) );
  NOR2_X1 NOR2_1393( .ZN(g28760), .A1(g15142), .A2(g28453) );
  NOR2_X1 NOR2_1394( .ZN(g28761), .A1(g28445), .A2(g27936) );
  NOR2_X1 NOR2_1395( .ZN(g28762), .A1(g28446), .A2(g27938) );
  NOR2_X1 NOR2_1396( .ZN(g28763), .A1(g15160), .A2(g28456) );
  NOR2_X1 NOR2_1397( .ZN(g28767), .A1(g28452), .A2(g27945) );
  NOR2_X1 NOR2_1398( .ZN(g28771), .A1(g15218), .A2(g28463) );
  NOR2_X1 NOR2_1399( .ZN(g28772), .A1(g28454), .A2(g27949) );
  NOR2_X1 NOR2_1400( .ZN(g28773), .A1(g15234), .A2(g28465) );
  NOR2_X1 NOR2_1401( .ZN(g28774), .A1(g28457), .A2(g27951) );
  NOR2_X1 NOR2_1402( .ZN(g28778), .A1(g28464), .A2(g27963) );
  NOR2_X1 NOR2_1403( .ZN(g28782), .A1(g15304), .A2(g28475) );
  NOR2_X1 NOR2_1404( .ZN(g28783), .A1(g28466), .A2(g27968) );
  NOR2_X1 NOR2_1405( .ZN(g28784), .A1(g28468), .A2(g27970) );
  NOR2_X1 NOR2_1406( .ZN(g28788), .A1(g28476), .A2(g27984) );
  NOR2_X1 NOR2_1407( .ZN(g28789), .A1(g28477), .A2(g27985) );
  NOR2_X1 NOR2_1408( .ZN(g28790), .A1(g28478), .A2(g27991) );
  NOR2_X2 NOR2_1409( .ZN(g28794), .A1(g28484), .A2(g28009) );
  NOR2_X2 NOR2_1410( .ZN(g28795), .A1(g28485), .A2(g28015) );
  NOR2_X1 NOR2_1411( .ZN(g28802), .A1(g28492), .A2(g28036) );
  NOR2_X1 NOR2_1412( .ZN(g28803), .A1(g28493), .A2(g28042) );
  NOR2_X1 NOR2_1413( .ZN(g28813), .A1(g28497), .A2(g28066) );
  NOR2_X1 NOR2_1414( .ZN(g28874), .A1(g28657), .A2(g16221) );
  NOR2_X1 NOR2_1415( .ZN(g28886), .A1(g28659), .A2(g16277) );
  NOR2_X1 NOR2_1416( .ZN(g28903), .A1(g28660), .A2(g13295) );
  NOR2_X1 NOR2_1417( .ZN(g28920), .A1(g28662), .A2(g13322) );
  NOR2_X1 NOR2_1418( .ZN(g28941), .A1(g28663), .A2(g13343) );
  NOR3_X1 NOR3_397( .ZN(g28954), .A1(g26673), .A2(g27241), .A3(g28323) );
  NOR2_X1 NOR2_1419( .ZN(g28963), .A1(g28664), .A2(g13365) );
  NOR2_X1 NOR2_1420( .ZN(g28982), .A1(g28665), .A2(g28670) );
  NOR2_X1 NOR2_1421( .ZN(g28987), .A1(g28666), .A2(g13390) );
  NOR2_X1 NOR2_1422( .ZN(g28990), .A1(g28667), .A2(g16457) );
  NOR2_X1 NOR2_1423( .ZN(g29009), .A1(g28669), .A2(g28320) );
  NOR2_X1 NOR2_1424( .ZN(g29013), .A1(g28671), .A2(g11607) );
  NOR2_X1 NOR2_1425( .ZN(g29016), .A1(g28672), .A2(g13487) );
  NOR2_X1 NOR2_1426( .ZN(g29031), .A1(g28319), .A2(g28324) );
  NOR2_X1 NOR2_1427( .ZN(g29039), .A1(g28322), .A2(g13500) );
  NOR2_X1 NOR2_1428( .ZN(g29063), .A1(g28326), .A2(g28329) );
  NOR2_X1 NOR2_1429( .ZN(g29064), .A1(g28327), .A2(g28330) );
  NOR2_X1 NOR2_1430( .ZN(g29083), .A1(g28331), .A2(g28333) );
  NOR2_X1 NOR2_1431( .ZN(g29090), .A1(g28332), .A2(g28334) );
  NOR2_X1 NOR2_1432( .ZN(g29097), .A1(g28335), .A2(g28336) );
  NOR2_X1 NOR2_1433( .ZN(g29109), .A1(g28654), .A2(g17001) );
  NOR2_X1 NOR2_1434( .ZN(g29110), .A1(g28656), .A2(g17031) );
  NOR2_X1 NOR2_1435( .ZN(g29111), .A1(g28658), .A2(g17065) );
  NOR2_X1 NOR2_1436( .ZN(g29112), .A1(g28661), .A2(g17100) );
  NOR2_X1 NOR2_1437( .ZN(g29113), .A1(g28381), .A2(g8907) );
  NOR2_X1 NOR2_1438( .ZN(g29126), .A1(g28373), .A2(g27774) );
  NOR2_X1 NOR2_1439( .ZN(g29127), .A1(g28376), .A2(g27779) );
  NOR2_X1 NOR2_1440( .ZN(g29128), .A1(g28380), .A2(g27783) );
  NOR2_X1 NOR2_1441( .ZN(g29129), .A1(g28385), .A2(g27790) );
  NOR2_X1 NOR2_1442( .ZN(g29167), .A1(g28841), .A2(g28396) );
  NOR2_X1 NOR2_1443( .ZN(g29169), .A1(g28843), .A2(g28398) );
  NOR2_X1 NOR2_1444( .ZN(g29170), .A1(g28844), .A2(g28399) );
  NOR2_X1 NOR2_1445( .ZN(g29172), .A1(g28846), .A2(g28401) );
  NOR2_X1 NOR2_1446( .ZN(g29173), .A1(g28847), .A2(g28402) );
  NOR2_X1 NOR2_1447( .ZN(g29178), .A1(g28848), .A2(g28404) );
  NOR2_X1 NOR2_1448( .ZN(g29179), .A1(g28849), .A2(g28405) );
  NOR2_X1 NOR2_1449( .ZN(g29181), .A1(g28850), .A2(g28407) );
  NOR2_X1 NOR2_1450( .ZN(g29182), .A1(g28851), .A2(g28408) );
  NOR2_X1 NOR2_1451( .ZN(g29184), .A1(g28852), .A2(g28411) );
  NOR2_X1 NOR2_1452( .ZN(g29185), .A1(g28853), .A2(g28412) );
  NOR2_X1 NOR2_1453( .ZN(g29187), .A1(g28854), .A2(g28416) );
  NOR2_X1 NOR2_1454( .ZN(g29194), .A1(g14958), .A2(g28881) );
  NOR2_X1 NOR2_1455( .ZN(g29195), .A1(g28880), .A2(g28438) );
  NOR2_X1 NOR2_1456( .ZN(g29197), .A1(g15031), .A2(g28893) );
  NOR2_X1 NOR2_1457( .ZN(g29198), .A1(g15047), .A2(g28898) );
  NOR2_X1 NOR2_1458( .ZN(g29199), .A1(g28892), .A2(g28448) );
  NOR2_X1 NOR2_1459( .ZN(g29201), .A1(g15104), .A2(g28910) );
  NOR2_X1 NOR2_1460( .ZN(g29202), .A1(g28897), .A2(g28450) );
  NOR2_X2 NOR2_1461( .ZN(g29204), .A1(g15127), .A2(g28915) );
  NOR2_X1 NOR2_1462( .ZN(g29205), .A1(g15143), .A2(g28923) );
  NOR2_X1 NOR2_1463( .ZN(g29206), .A1(g28909), .A2(g28459) );
  NOR2_X1 NOR2_1464( .ZN(g29207), .A1(g28914), .A2(g28460) );
  NOR2_X1 NOR2_1465( .ZN(g29209), .A1(g15196), .A2(g28936) );
  NOR2_X1 NOR2_1466( .ZN(g29210), .A1(g28919), .A2(g28462) );
  NOR2_X1 NOR2_1467( .ZN(g29212), .A1(g15219), .A2(g28944) );
  NOR2_X1 NOR2_1468( .ZN(g29213), .A1(g15235), .A2(g28949) );
  NOR2_X1 NOR2_1469( .ZN(g29214), .A1(g28931), .A2(g28469) );
  NOR2_X1 NOR2_1470( .ZN(g29215), .A1(g28935), .A2(g28471) );
  NOR2_X1 NOR2_1471( .ZN(g29216), .A1(g28940), .A2(g28472) );
  NOR2_X1 NOR2_1472( .ZN(g29218), .A1(g15282), .A2(g28966) );
  NOR2_X1 NOR2_1473( .ZN(g29219), .A1(g28948), .A2(g28474) );
  NOR2_X1 NOR2_1474( .ZN(g29221), .A1(g15305), .A2(g28971) );
  NOR2_X1 NOR2_1475( .ZN(g29222), .A1(g28958), .A2(g28479) );
  NOR2_X1 NOR2_1476( .ZN(g29223), .A1(g28962), .A2(g28480) );
  NOR2_X1 NOR2_1477( .ZN(g29224), .A1(g28970), .A2(g28481) );
  NOR2_X1 NOR2_1478( .ZN(g29226), .A1(g15374), .A2(g28997) );
  NOR2_X1 NOR2_1479( .ZN(g29227), .A1(g28986), .A2(g28486) );
  NOR2_X1 NOR2_1480( .ZN(g29228), .A1(g28996), .A2(g28487) );
  NOR2_X1 NOR2_1481( .ZN(g29231), .A1(g29022), .A2(g28494) );
  NOR2_X1 NOR2_1482( .ZN(g29303), .A1(g28716), .A2(g19112) );
  NOR2_X1 NOR2_1483( .ZN(g29313), .A1(g28717), .A2(g19117) );
  NOR2_X1 NOR2_1484( .ZN(g29324), .A1(g28718), .A2(g19124) );
  NOR2_X1 NOR2_1485( .ZN(g29333), .A1(g28719), .A2(g19131) );
  NOR2_X1 NOR2_1486( .ZN(g29340), .A1(g28337), .A2(g28722) );
  NOR2_X1 NOR2_1487( .ZN(g29343), .A1(g28338), .A2(g28724) );
  NOR2_X1 NOR2_1488( .ZN(g29345), .A1(g28339), .A2(g28726) );
  NOR2_X1 NOR2_1489( .ZN(g29347), .A1(g28340), .A2(g28729) );
  NOR2_X1 NOR2_1490( .ZN(g29353), .A1(g29126), .A2(g17001) );
  NOR2_X1 NOR2_1491( .ZN(g29354), .A1(g29127), .A2(g17031) );
  NOR2_X1 NOR2_1492( .ZN(g29355), .A1(g29128), .A2(g17065) );
  NOR2_X1 NOR2_1493( .ZN(g29357), .A1(g29129), .A2(g17100) );
  NOR2_X1 NOR2_1494( .ZN(g29399), .A1(g28834), .A2(g28378) );
  NOR2_X1 NOR2_1495( .ZN(g29403), .A1(g28836), .A2(g28383) );
  NOR2_X1 NOR2_1496( .ZN(g29406), .A1(g28838), .A2(g28387) );
  NOR2_X1 NOR2_1497( .ZN(g29409), .A1(g28840), .A2(g28389) );
  NOR2_X1 NOR2_1498( .ZN(g29552), .A1(g29130), .A2(g29411) );
  NOR2_X1 NOR2_1499( .ZN(g29569), .A1(g28708), .A2(g29174) );
  NOR2_X1 NOR2_1500( .ZN(g29570), .A1(g28709), .A2(g29175) );
  NOR2_X1 NOR2_1501( .ZN(g29571), .A1(g28710), .A2(g29176) );
  NOR2_X1 NOR2_1502( .ZN(g29574), .A1(g28712), .A2(g29180) );
  NOR2_X1 NOR2_1503( .ZN(g29576), .A1(g28713), .A2(g29183) );
  NOR2_X1 NOR2_1504( .ZN(g29577), .A1(g28714), .A2(g29186) );
  NOR2_X1 NOR2_1505( .ZN(g29578), .A1(g28715), .A2(g29188) );
  NOR2_X1 NOR2_1506( .ZN(g29579), .A1(g29399), .A2(g17001) );
  NOR2_X1 NOR2_1507( .ZN(g29580), .A1(g29403), .A2(g17031) );
  NOR2_X1 NOR2_1508( .ZN(g29581), .A1(g29406), .A2(g17065) );
  NOR2_X1 NOR2_1509( .ZN(g29582), .A1(g29409), .A2(g17100) );
  NOR2_X1 NOR2_1510( .ZN(g29606), .A1(g13878), .A2(g29248) );
  NOR2_X1 NOR2_1511( .ZN(g29608), .A1(g13892), .A2(g29251) );
  NOR2_X1 NOR2_1512( .ZN(g29609), .A1(g13900), .A2(g29252) );
  NOR2_X1 NOR2_1513( .ZN(g29611), .A1(g13913), .A2(g29255) );
  NOR2_X1 NOR2_1514( .ZN(g29612), .A1(g13933), .A2(g29256) );
  NOR2_X1 NOR2_1515( .ZN(g29613), .A1(g13941), .A2(g29257) );
  NOR2_X1 NOR2_1516( .ZN(g29616), .A1(g13969), .A2(g29259) );
  NOR2_X1 NOR2_1517( .ZN(g29617), .A1(g13989), .A2(g29260) );
  NOR2_X1 NOR2_1518( .ZN(g29618), .A1(g13997), .A2(g29261) );
  NOR2_X1 NOR2_1519( .ZN(g29620), .A1(g14039), .A2(g29262) );
  NOR2_X1 NOR2_1520( .ZN(g29621), .A1(g14059), .A2(g29263) );
  NOR2_X2 NOR2_1521( .ZN(g29623), .A1(g14130), .A2(g29264) );
  NOR2_X1 NOR2_1522( .ZN(g29663), .A1(g29518), .A2(g29284) );
  NOR2_X1 NOR2_1523( .ZN(g29665), .A1(g29521), .A2(g29289) );
  NOR2_X1 NOR2_1524( .ZN(g29667), .A1(g29524), .A2(g29294) );
  NOR2_X1 NOR2_1525( .ZN(g29669), .A1(g29528), .A2(g29300) );
  NOR2_X1 NOR2_1526( .ZN(g29670), .A1(g29529), .A2(g29302) );
  NOR2_X1 NOR2_1527( .ZN(g29671), .A1(g29534), .A2(g29310) );
  NOR2_X1 NOR2_1528( .ZN(g29672), .A1(g29536), .A2(g29312) );
  NOR2_X1 NOR2_1529( .ZN(g29676), .A1(g29540), .A2(g29320) );
  NOR2_X1 NOR2_1530( .ZN(g29677), .A1(g29543), .A2(g29321) );
  NOR2_X1 NOR2_1531( .ZN(g29678), .A1(g29545), .A2(g29323) );
  NOR2_X1 NOR2_1532( .ZN(g29679), .A1(g29549), .A2(g29329) );
  NOR2_X1 NOR2_1533( .ZN(g29680), .A1(g29553), .A2(g29330) );
  NOR2_X1 NOR2_1534( .ZN(g29681), .A1(g29555), .A2(g29332) );
  NOR2_X1 NOR2_1535( .ZN(g29682), .A1(g29557), .A2(g29336) );
  NOR2_X1 NOR2_1536( .ZN(g29683), .A1(g29559), .A2(g29337) );
  NOR2_X1 NOR2_1537( .ZN(g29684), .A1(g29562), .A2(g29338) );
  NOR2_X1 NOR2_1538( .ZN(g29685), .A1(g29564), .A2(g29341) );
  NOR2_X1 NOR2_1539( .ZN(g29686), .A1(g29566), .A2(g29342) );
  NOR2_X1 NOR2_1540( .ZN(g29687), .A1(g29572), .A2(g29344) );
  NOR2_X1 NOR2_1541( .ZN(g29688), .A1(g29575), .A2(g29346) );
  NOR2_X1 NOR2_1542( .ZN(g29703), .A1(g29583), .A2(g1917) );
  NOR3_X1 NOR3_398( .ZN(g29705), .A1(g6104), .A2(g29583), .A3(g25339) );
  NOR2_X1 NOR2_1543( .ZN(g29709), .A1(g29583), .A2(g1909) );
  NOR3_X1 NOR3_399( .ZN(g29710), .A1(g6104), .A2(g29583), .A3(g25412) );
  NOR3_X1 NOR3_400( .ZN(g29713), .A1(g6104), .A2(g29583), .A3(g25332) );
  NOR2_X1 NOR2_1544( .ZN(g29717), .A1(g29583), .A2(g1910) );
  NOR3_X1 NOR3_401( .ZN(g29718), .A1(g6104), .A2(g29583), .A3(g25409) );
  NOR3_X1 NOR3_402( .ZN(g29721), .A1(g6104), .A2(g29583), .A3(g25323) );
  NOR2_X1 NOR2_1545( .ZN(g29725), .A1(g29583), .A2(g1911) );
  NOR2_X1 NOR2_1546( .ZN(g29727), .A1(g29583), .A2(g1912) );
  NOR3_X1 NOR3_403( .ZN(g29728), .A1(g6104), .A2(g29583), .A3(g25401) );
  NOR2_X1 NOR2_1547( .ZN(g29731), .A1(g29583), .A2(g1913) );
  NOR3_X1 NOR3_404( .ZN(g29732), .A1(g6104), .A2(g29583), .A3(g25387) );
  NOR2_X1 NOR2_1548( .ZN(g29735), .A1(g23797), .A2(g29583) );
  NOR2_X1 NOR2_1549( .ZN(g29736), .A1(g29583), .A2(g25444) );
  NOR2_X1 NOR2_1550( .ZN(g29740), .A1(g29583), .A2(g1914) );
  NOR3_X1 NOR3_405( .ZN(g29741), .A1(g6104), .A2(g29583), .A3(g25376) );
  NOR2_X1 NOR2_1551( .ZN(g29744), .A1(g29583), .A2(g24641) );
  NOR2_X1 NOR2_1552( .ZN(g29747), .A1(g29583), .A2(g1916) );
  NOR3_X1 NOR3_406( .ZN(g29748), .A1(g6104), .A2(g29583), .A3(g25363) );
  NOR3_X1 NOR3_407( .ZN(g29751), .A1(g6104), .A2(g29583), .A3(g25352) );
  NOR2_X1 NOR2_1553( .ZN(g29754), .A1(g16178), .A2(g29607) );
  NOR2_X1 NOR2_1554( .ZN(g29755), .A1(g16229), .A2(g29610) );
  NOR2_X1 NOR2_1555( .ZN(g29756), .A1(g16284), .A2(g29614) );
  NOR2_X1 NOR2_1556( .ZN(g29757), .A1(g16285), .A2(g29615) );
  NOR2_X1 NOR2_1557( .ZN(g29758), .A1(g16335), .A2(g29619) );
  NOR2_X1 NOR2_1558( .ZN(g29759), .A1(g16379), .A2(g29622) );
  NOR2_X1 NOR2_1559( .ZN(g29760), .A1(g16411), .A2(g29624) );
  NOR3_X1 NOR3_408( .ZN(g29761), .A1(g28707), .A2(g28711), .A3(g29466) );
  NOR2_X1 NOR2_1560( .ZN(g29762), .A1(g16432), .A2(g29625) );
  NOR2_X1 NOR2_1561( .ZN(g29763), .A1(g16438), .A2(g29626) );
  NOR2_X1 NOR2_1562( .ZN(g29764), .A1(g16462), .A2(g29464) );
  NOR2_X1 NOR2_1563( .ZN(g29765), .A1(g13492), .A2(g29465) );
  NOR2_X1 NOR2_1564( .ZN(g29766), .A1(g29467), .A2(g19142) );
  NOR2_X1 NOR2_1565( .ZN(g29767), .A1(g29468), .A2(g19143) );
  NOR2_X1 NOR2_1566( .ZN(g29768), .A1(g29469), .A2(g19146) );
  NOR2_X1 NOR2_1567( .ZN(g29769), .A1(g29470), .A2(g19148) );
  NOR2_X1 NOR2_1568( .ZN(g29770), .A1(g29471), .A2(g29196) );
  NOR2_X1 NOR2_1569( .ZN(g29771), .A1(g29472), .A2(g29200) );
  NOR2_X1 NOR2_1570( .ZN(g29772), .A1(g29473), .A2(g29203) );
  NOR2_X1 NOR2_1571( .ZN(g29773), .A1(g29474), .A2(g29208) );
  NOR2_X1 NOR2_1572( .ZN(g29774), .A1(g29475), .A2(g29211) );
  NOR2_X2 NOR2_1573( .ZN(g29775), .A1(g29476), .A2(g29217) );
  NOR2_X1 NOR2_1574( .ZN(g29776), .A1(g29477), .A2(g29220) );
  NOR2_X1 NOR2_1575( .ZN(g29777), .A1(g29478), .A2(g29225) );
  NOR2_X1 NOR2_1576( .ZN(g29778), .A1(g29479), .A2(g29229) );
  NOR2_X1 NOR2_1577( .ZN(g29779), .A1(g13943), .A2(g29502) );
  NOR2_X1 NOR2_1578( .ZN(g29780), .A1(g29480), .A2(g29232) );
  NOR2_X1 NOR2_1579( .ZN(g29781), .A1(g29481), .A2(g29233) );
  NOR2_X1 NOR2_1580( .ZN(g29782), .A1(g29482), .A2(g29234) );
  NOR2_X1 NOR2_1581( .ZN(g29783), .A1(g29483), .A2(g29235) );
  NOR2_X1 NOR2_1582( .ZN(g29784), .A1(g29484), .A2(g29236) );
  NOR2_X1 NOR2_1583( .ZN(g29785), .A1(g29485), .A2(g29238) );
  NOR2_X1 NOR2_1584( .ZN(g29786), .A1(g29486), .A2(g29239) );
  NOR2_X1 NOR2_1585( .ZN(g29787), .A1(g29487), .A2(g29240) );
  NOR2_X1 NOR2_1586( .ZN(g29788), .A1(g29488), .A2(g29241) );
  NOR2_X1 NOR2_1587( .ZN(g29789), .A1(g29489), .A2(g29242) );
  NOR2_X1 NOR2_1588( .ZN(g29791), .A1(g29490), .A2(g29243) );
  NOR2_X1 NOR2_1589( .ZN(g29912), .A1(g24676), .A2(g29716) );
  NOR2_X1 NOR2_1590( .ZN(g29914), .A1(g24695), .A2(g29724) );
  NOR2_X1 NOR2_1591( .ZN(g29916), .A1(g24712), .A2(g29726) );
  NOR2_X1 NOR2_1592( .ZN(g29918), .A1(g29744), .A2(g22367) );
  NOR2_X1 NOR2_1593( .ZN(g29919), .A1(g29736), .A2(g22367) );
  NOR2_X1 NOR2_1594( .ZN(g29920), .A1(g24723), .A2(g29739) );
  NOR2_X1 NOR2_1595( .ZN(g29921), .A1(g29736), .A2(g22367) );
  NOR2_X1 NOR2_1596( .ZN(g29922), .A1(g29744), .A2(g22367) );
  NOR2_X1 NOR2_1597( .ZN(g29924), .A1(g29710), .A2(g22367) );
  NOR2_X1 NOR2_1598( .ZN(g29926), .A1(g29718), .A2(g22367) );
  NOR2_X1 NOR2_1599( .ZN(g29928), .A1(g29673), .A2(g22367) );
  NOR2_X1 NOR2_1600( .ZN(g29929), .A1(g29673), .A2(g22367) );
  NOR2_X1 NOR2_1601( .ZN(g29936), .A1(g16049), .A2(g29790) );
  NOR2_X1 NOR2_1602( .ZN(g29939), .A1(g16102), .A2(g29792) );
  NOR2_X1 NOR2_1603( .ZN(g29941), .A1(g16182), .A2(g29793) );
  NOR2_X1 NOR2_1604( .ZN(g30010), .A1(g29520), .A2(g29942) );
  NOR2_X1 NOR2_1605( .ZN(g30011), .A1(g29522), .A2(g29944) );
  NOR2_X1 NOR2_1606( .ZN(g30012), .A1(g29523), .A2(g29945) );
  NOR2_X1 NOR2_1607( .ZN(g30013), .A1(g29525), .A2(g29946) );
  NOR2_X1 NOR2_1608( .ZN(g30014), .A1(g29526), .A2(g29947) );
  NOR2_X1 NOR2_1609( .ZN(g30015), .A1(g29527), .A2(g29948) );
  NOR2_X1 NOR2_1610( .ZN(g30016), .A1(g29531), .A2(g29949) );
  NOR2_X1 NOR2_1611( .ZN(g30017), .A1(g29532), .A2(g29950) );
  NOR2_X1 NOR2_1612( .ZN(g30018), .A1(g29533), .A2(g29951) );
  NOR2_X1 NOR2_1613( .ZN(g30019), .A1(g29538), .A2(g29952) );
  NOR2_X1 NOR2_1614( .ZN(g30020), .A1(g29539), .A2(g29953) );
  NOR2_X1 NOR2_1615( .ZN(g30021), .A1(g29541), .A2(g29954) );
  NOR2_X1 NOR2_1616( .ZN(g30022), .A1(g29547), .A2(g29955) );
  NOR2_X1 NOR2_1617( .ZN(g30023), .A1(g29548), .A2(g29956) );
  NOR2_X1 NOR2_1618( .ZN(g30024), .A1(g29550), .A2(g29957) );
  NOR2_X1 NOR2_1619( .ZN(g30025), .A1(g29558), .A2(g29958) );
  NOR2_X1 NOR2_1620( .ZN(g30026), .A1(g29560), .A2(g29959) );
  NOR2_X1 NOR2_1621( .ZN(g30027), .A1(g29565), .A2(g29960) );
  NOR2_X1 NOR2_1622( .ZN(g30028), .A1(g29567), .A2(g29961) );
  NOR2_X1 NOR2_1623( .ZN(g30029), .A1(g29573), .A2(g29962) );
  NOR2_X1 NOR2_1624( .ZN(g30030), .A1(g24676), .A2(g29923) );
  NOR2_X1 NOR2_1625( .ZN(g30031), .A1(g24695), .A2(g29925) );
  NOR2_X1 NOR2_1626( .ZN(g30032), .A1(g24712), .A2(g29927) );
  NOR2_X1 NOR2_1627( .ZN(g30033), .A1(g24723), .A2(g29931) );
  NOR2_X1 NOR2_1628( .ZN(g30053), .A1(g29963), .A2(g16286) );
  NOR2_X1 NOR2_1629( .ZN(g30054), .A1(g29964), .A2(g16336) );
  NOR2_X1 NOR2_1630( .ZN(g30055), .A1(g29965), .A2(g13326) );
  NOR2_X1 NOR2_1631( .ZN(g30056), .A1(g29966), .A2(g13345) );
  NOR2_X1 NOR2_1632( .ZN(g30057), .A1(g29967), .A2(g13368) );
  NOR2_X1 NOR2_1633( .ZN(g30058), .A1(g29968), .A2(g13395) );
  NOR2_X1 NOR2_1634( .ZN(g30059), .A1(g29969), .A2(g29811) );
  NOR2_X1 NOR2_1635( .ZN(g30060), .A1(g29970), .A2(g11612) );
  NOR2_X1 NOR2_1636( .ZN(g30061), .A1(g29971), .A2(g13493) );
  NOR2_X1 NOR2_1637( .ZN(g30062), .A1(g29810), .A2(g29815) );
  NOR2_X1 NOR2_1638( .ZN(g30063), .A1(g29812), .A2(g11637) );
  NOR2_X1 NOR2_1639( .ZN(g30064), .A1(g29813), .A2(g13506) );
  NOR2_X1 NOR2_1640( .ZN(g30065), .A1(g29814), .A2(g29817) );
  NOR2_X1 NOR2_1641( .ZN(g30066), .A1(g29816), .A2(g13517) );
  NOR2_X1 NOR2_1642( .ZN(g30067), .A1(g29818), .A2(g29820) );
  NOR2_X1 NOR2_1643( .ZN(g30068), .A1(g29819), .A2(g29821) );
  NOR2_X1 NOR2_1644( .ZN(g30069), .A1(g29822), .A2(g29828) );
  NOR2_X1 NOR2_1645( .ZN(g30070), .A1(g29827), .A2(g29833) );
  NOR2_X1 NOR2_1646( .ZN(g30071), .A1(g29834), .A2(g29839) );
  NOR2_X1 NOR2_1647( .ZN(g30072), .A1(g29910), .A2(g8947) );
  NOR2_X1 NOR2_1648( .ZN(g30245), .A1(g16074), .A2(g30077) );
  NOR2_X1 NOR2_1649( .ZN(g30246), .A1(g16107), .A2(g30079) );
  NOR2_X1 NOR2_1650( .ZN(g30247), .A1(g16112), .A2(g30080) );
  NOR2_X1 NOR2_1651( .ZN(g30248), .A1(g16139), .A2(g30081) );
  NOR2_X1 NOR2_1652( .ZN(g30249), .A1(g16158), .A2(g30082) );
  NOR2_X1 NOR2_1653( .ZN(g30250), .A1(g16163), .A2(g30083) );
  NOR2_X1 NOR2_1654( .ZN(g30251), .A1(g16198), .A2(g30085) );
  NOR2_X1 NOR2_1655( .ZN(g30252), .A1(g16217), .A2(g30086) );
  NOR2_X1 NOR2_1656( .ZN(g30253), .A1(g16222), .A2(g30087) );
  NOR2_X1 NOR2_1657( .ZN(g30254), .A1(g16242), .A2(g30088) );
  NOR2_X1 NOR2_1658( .ZN(g30255), .A1(g16263), .A2(g30089) );
  NOR2_X1 NOR2_1659( .ZN(g30256), .A1(g16282), .A2(g30090) );
  NOR2_X1 NOR2_1660( .ZN(g30257), .A1(g16290), .A2(g30091) );
  NOR2_X1 NOR2_1661( .ZN(g30258), .A1(g16291), .A2(g30092) );
  NOR2_X1 NOR2_1662( .ZN(g30259), .A1(g16301), .A2(g30093) );
  NOR2_X1 NOR2_1663( .ZN(g30260), .A1(g16322), .A2(g30094) );
  NOR2_X1 NOR2_1664( .ZN(g30261), .A1(g16342), .A2(g30095) );
  NOR2_X1 NOR2_1665( .ZN(g30262), .A1(g16343), .A2(g30096) );
  NOR2_X1 NOR2_1666( .ZN(g30263), .A1(g16344), .A2(g30097) );
  NOR2_X1 NOR2_1667( .ZN(g30264), .A1(g16348), .A2(g30098) );
  NOR2_X1 NOR2_1668( .ZN(g30265), .A1(g16349), .A2(g30099) );
  NOR2_X1 NOR2_1669( .ZN(g30266), .A1(g16359), .A2(g30100) );
  NOR2_X1 NOR2_1670( .ZN(g30267), .A1(g16380), .A2(g30101) );
  NOR2_X1 NOR2_1671( .ZN(g30268), .A1(g16382), .A2(g30102) );
  NOR2_X1 NOR2_1672( .ZN(g30269), .A1(g16386), .A2(g30103) );
  NOR2_X1 NOR2_1673( .ZN(g30270), .A1(g16387), .A2(g30104) );
  NOR2_X1 NOR2_1674( .ZN(g30271), .A1(g16388), .A2(g30105) );
  NOR2_X1 NOR2_1675( .ZN(g30272), .A1(g16392), .A2(g30106) );
  NOR2_X1 NOR2_1676( .ZN(g30273), .A1(g16393), .A2(g30107) );
  NOR2_X1 NOR2_1677( .ZN(g30274), .A1(g16403), .A2(g30108) );
  NOR2_X1 NOR2_1678( .ZN(g30275), .A1(g16413), .A2(g30109) );
  NOR2_X1 NOR2_1679( .ZN(g30276), .A1(g16415), .A2(g30110) );
  NOR2_X1 NOR2_1680( .ZN(g30277), .A1(g16418), .A2(g30111) );
  NOR2_X1 NOR2_1681( .ZN(g30278), .A1(g16420), .A2(g30112) );
  NOR2_X1 NOR2_1682( .ZN(g30279), .A1(g16424), .A2(g30113) );
  NOR2_X1 NOR2_1683( .ZN(g30280), .A1(g16425), .A2(g30114) );
  NOR2_X1 NOR2_1684( .ZN(g30281), .A1(g16426), .A2(g30115) );
  NOR2_X1 NOR2_1685( .ZN(g30282), .A1(g16430), .A2(g30117) );
  NOR2_X1 NOR2_1686( .ZN(g30283), .A1(g16431), .A2(g30118) );
  NOR2_X1 NOR2_1687( .ZN(g30284), .A1(g16444), .A2(g29980) );
  NOR2_X1 NOR2_1688( .ZN(g30285), .A1(g16447), .A2(g29981) );
  NOR2_X1 NOR2_1689( .ZN(g30286), .A1(g16449), .A2(g29982) );
  NOR2_X1 NOR2_1690( .ZN(g30287), .A1(g16452), .A2(g29983) );
  NOR2_X1 NOR2_1691( .ZN(g30288), .A1(g16454), .A2(g29984) );
  NOR2_X1 NOR2_1692( .ZN(g30289), .A1(g16458), .A2(g29985) );
  NOR2_X1 NOR2_1693( .ZN(g30290), .A1(g16459), .A2(g29986) );
  NOR2_X1 NOR2_1694( .ZN(g30291), .A1(g16460), .A2(g29987) );
  NOR2_X1 NOR2_1695( .ZN(g30292), .A1(g13477), .A2(g29988) );
  NOR2_X1 NOR2_1696( .ZN(g30293), .A1(g13480), .A2(g29989) );
  NOR2_X1 NOR2_1697( .ZN(g30294), .A1(g13483), .A2(g29990) );
  NOR2_X1 NOR2_1698( .ZN(g30295), .A1(g13485), .A2(g29991) );
  NOR2_X1 NOR2_1699( .ZN(g30296), .A1(g13488), .A2(g29993) );
  NOR2_X1 NOR2_1700( .ZN(g30297), .A1(g13490), .A2(g29994) );
  NOR2_X1 NOR2_1701( .ZN(g30298), .A1(g13496), .A2(g29995) );
  NOR2_X1 NOR2_1702( .ZN(g30299), .A1(g13499), .A2(g29996) );
  NOR2_X1 NOR2_1703( .ZN(g30300), .A1(g13502), .A2(g30001) );
  NOR2_X1 NOR2_1704( .ZN(g30301), .A1(g13504), .A2(g30002) );
  NOR2_X1 NOR2_1705( .ZN(g30302), .A1(g13513), .A2(g30003) );
  NOR2_X1 NOR2_1706( .ZN(g30303), .A1(g13516), .A2(g30005) );
  NOR2_X1 NOR2_1707( .ZN(g30304), .A1(g13527), .A2(g30007) );
  NOR2_X1 NOR2_1708( .ZN(g30338), .A1(g14297), .A2(g30225) );
  NOR2_X1 NOR2_1709( .ZN(g30341), .A1(g14328), .A2(g30226) );
  NOR2_X1 NOR2_1710( .ZN(g30356), .A1(g14419), .A2(g30227) );
  NOR2_X1 NOR2_1711( .ZN(g30399), .A1(g30116), .A2(g30123) );
  NOR2_X1 NOR2_1712( .ZN(g30400), .A1(g29997), .A2(g30127) );
  NOR2_X1 NOR2_1713( .ZN(g30401), .A1(g29998), .A2(g30128) );
  NOR2_X1 NOR2_1714( .ZN(g30402), .A1(g29999), .A2(g30129) );
  NOR2_X1 NOR2_1715( .ZN(g30403), .A1(g30004), .A2(g30131) );
  NOR2_X1 NOR2_1716( .ZN(g30404), .A1(g30006), .A2(g30132) );
  NOR2_X1 NOR2_1717( .ZN(g30405), .A1(g30008), .A2(g30133) );
  NOR2_X1 NOR2_1718( .ZN(g30406), .A1(g30009), .A2(g30138) );
  NOR2_X1 NOR2_1719( .ZN(g30455), .A1(g13953), .A2(g30216) );
  NOR2_X1 NOR2_1720( .ZN(g30468), .A1(g14007), .A2(g30217) );
  NOR2_X1 NOR2_1721( .ZN(g30470), .A1(g14023), .A2(g30218) );
  NOR2_X1 NOR2_1722( .ZN(g30482), .A1(g14067), .A2(g30219) );
  NOR2_X1 NOR2_1723( .ZN(g30485), .A1(g14098), .A2(g30220) );
  NOR2_X1 NOR2_1724( .ZN(g30487), .A1(g14114), .A2(g30221) );
  NOR2_X1 NOR2_1725( .ZN(g30500), .A1(g14182), .A2(g30222) );
  NOR2_X1 NOR2_1726( .ZN(g30503), .A1(g14213), .A2(g30223) );
  NOR2_X1 NOR2_1727( .ZN(g30505), .A1(g14229), .A2(g30224) );
  NOR2_X2 NOR2_1728( .ZN(g30566), .A1(g14327), .A2(g30398) );
  NOR2_X2 NOR2_1729( .ZN(g30584), .A1(g30412), .A2(g2611) );
  NOR3_X1 NOR3_409( .ZN(g30588), .A1(g6119), .A2(g30412), .A3(g25353) );
  NOR2_X2 NOR2_1730( .ZN(g30593), .A1(g30412), .A2(g2603) );
  NOR3_X1 NOR3_410( .ZN(g30594), .A1(g6119), .A2(g30412), .A3(g25419) );
  NOR3_X1 NOR3_411( .ZN(g30597), .A1(g6119), .A2(g30412), .A3(g25341) );
  NOR2_X2 NOR2_1731( .ZN(g30601), .A1(g30412), .A2(g2604) );
  NOR3_X2 NOR3_412( .ZN(g30602), .A1(g6119), .A2(g30412), .A3(g25417) );
  NOR3_X2 NOR3_413( .ZN(g30605), .A1(g6119), .A2(g30412), .A3(g25333) );
  NOR2_X2 NOR2_1732( .ZN(g30608), .A1(g30412), .A2(g2605) );
  NOR2_X1 NOR2_1733( .ZN(g30609), .A1(g30412), .A2(g2606) );
  NOR3_X1 NOR3_414( .ZN(g30610), .A1(g6119), .A2(g30412), .A3(g25411) );
  NOR2_X1 NOR2_1734( .ZN(g30613), .A1(g30412), .A2(g2607) );
  NOR3_X1 NOR3_415( .ZN(g30614), .A1(g6119), .A2(g30412), .A3(g25403) );
  NOR2_X1 NOR2_1735( .ZN(g30617), .A1(g23850), .A2(g30412) );
  NOR2_X1 NOR2_1736( .ZN(g30618), .A1(g30412), .A2(g25449) );
  NOR2_X1 NOR2_1737( .ZN(g30621), .A1(g30412), .A2(g2608) );
  NOR3_X1 NOR3_416( .ZN(g30622), .A1(g6119), .A2(g30412), .A3(g25393) );
  NOR2_X1 NOR2_1738( .ZN(g30625), .A1(g30412), .A2(g24660) );
  NOR2_X1 NOR2_1739( .ZN(g30628), .A1(g30412), .A2(g2610) );
  NOR3_X1 NOR3_417( .ZN(g30629), .A1(g6119), .A2(g30412), .A3(g25378) );
  NOR3_X1 NOR3_418( .ZN(g30632), .A1(g6119), .A2(g30412), .A3(g25366) );
  NOR2_X1 NOR2_1740( .ZN(g30635), .A1(g16108), .A2(g30407) );
  NOR2_X1 NOR2_1741( .ZN(g30636), .A1(g16140), .A2(g30409) );
  NOR2_X1 NOR2_1742( .ZN(g30637), .A1(g16141), .A2(g30410) );
  NOR2_X1 NOR2_1743( .ZN(g30638), .A1(g16159), .A2(g30411) );
  NOR2_X1 NOR2_1744( .ZN(g30639), .A1(g16186), .A2(g30436) );
  NOR2_X1 NOR2_1745( .ZN(g30640), .A1(g16187), .A2(g30437) );
  NOR2_X1 NOR2_1746( .ZN(g30641), .A1(g16188), .A2(g30438) );
  NOR2_X1 NOR2_1747( .ZN(g30642), .A1(g16199), .A2(g30440) );
  NOR2_X1 NOR2_1748( .ZN(g30643), .A1(g16200), .A2(g30441) );
  NOR2_X1 NOR2_1749( .ZN(g30644), .A1(g16218), .A2(g30442) );
  NOR2_X1 NOR2_1750( .ZN(g30645), .A1(g16240), .A2(g30444) );
  NOR2_X1 NOR2_1751( .ZN(g30646), .A1(g16241), .A2(g30445) );
  NOR2_X1 NOR2_1752( .ZN(g30647), .A1(g16251), .A2(g30447) );
  NOR2_X1 NOR2_1753( .ZN(g30648), .A1(g16252), .A2(g30448) );
  NOR2_X1 NOR2_1754( .ZN(g30649), .A1(g16253), .A2(g30449) );
  NOR2_X1 NOR2_1755( .ZN(g30650), .A1(g16264), .A2(g30451) );
  NOR2_X1 NOR2_1756( .ZN(g30651), .A1(g16265), .A2(g30452) );
  NOR2_X1 NOR2_1757( .ZN(g30652), .A1(g16283), .A2(g30453) );
  NOR2_X1 NOR2_1758( .ZN(g30653), .A1(g16289), .A2(g30454) );
  NOR2_X1 NOR2_1759( .ZN(g30654), .A1(g16299), .A2(g30457) );
  NOR2_X1 NOR2_1760( .ZN(g30655), .A1(g16300), .A2(g30458) );
  NOR2_X1 NOR2_1761( .ZN(g30656), .A1(g16310), .A2(g30460) );
  NOR2_X1 NOR2_1762( .ZN(g30657), .A1(g16311), .A2(g30461) );
  NOR2_X1 NOR2_1763( .ZN(g30658), .A1(g16312), .A2(g30462) );
  NOR2_X1 NOR2_1764( .ZN(g30659), .A1(g16323), .A2(g30464) );
  NOR2_X1 NOR2_1765( .ZN(g30660), .A1(g16324), .A2(g30465) );
  NOR2_X1 NOR2_1766( .ZN(g30661), .A1(g16345), .A2(g30467) );
  NOR2_X1 NOR2_1767( .ZN(g30662), .A1(g16347), .A2(g30469) );
  NOR2_X1 NOR2_1768( .ZN(g30663), .A1(g16357), .A2(g30472) );
  NOR2_X1 NOR2_1769( .ZN(g30664), .A1(g16358), .A2(g30473) );
  NOR2_X1 NOR2_1770( .ZN(g30665), .A1(g16368), .A2(g30475) );
  NOR2_X1 NOR2_1771( .ZN(g30666), .A1(g16369), .A2(g30476) );
  NOR2_X1 NOR2_1772( .ZN(g30667), .A1(g16370), .A2(g30477) );
  NOR2_X1 NOR2_1773( .ZN(g30668), .A1(g16381), .A2(g30478) );
  NOR2_X1 NOR2_1774( .ZN(g30669), .A1(g16383), .A2(g30481) );
  NOR2_X1 NOR2_1775( .ZN(g30670), .A1(g16389), .A2(g30484) );
  NOR2_X1 NOR2_1776( .ZN(g30671), .A1(g16391), .A2(g30486) );
  NOR2_X1 NOR2_1777( .ZN(g30672), .A1(g16401), .A2(g30489) );
  NOR2_X1 NOR2_1778( .ZN(g30673), .A1(g16402), .A2(g30490) );
  NOR2_X1 NOR2_1779( .ZN(g30674), .A1(g16414), .A2(g30492) );
  NOR2_X1 NOR2_1780( .ZN(g30675), .A1(g16416), .A2(g30495) );
  NOR2_X1 NOR2_1781( .ZN(g30676), .A1(g16419), .A2(g30496) );
  NOR2_X1 NOR2_1782( .ZN(g30677), .A1(g16421), .A2(g30499) );
  NOR2_X1 NOR2_1783( .ZN(g30678), .A1(g16427), .A2(g30502) );
  NOR2_X1 NOR2_1784( .ZN(g30679), .A1(g16429), .A2(g30504) );
  NOR2_X1 NOR2_1785( .ZN(g30680), .A1(g16443), .A2(g30327) );
  NOR2_X1 NOR2_1786( .ZN(g30681), .A1(g16448), .A2(g30330) );
  NOR2_X1 NOR2_1787( .ZN(g30682), .A1(g16450), .A2(g30333) );
  NOR2_X1 NOR2_1788( .ZN(g30683), .A1(g16453), .A2(g30334) );
  NOR2_X1 NOR2_1789( .ZN(g30684), .A1(g16455), .A2(g30337) );
  NOR3_X1 NOR3_419( .ZN(g30685), .A1(g29992), .A2(g30000), .A3(g30372) );
  NOR2_X1 NOR2_1790( .ZN(g30686), .A1(g16461), .A2(g30340) );
  NOR2_X1 NOR2_1791( .ZN(g30687), .A1(g13479), .A2(g30345) );
  NOR2_X1 NOR2_1792( .ZN(g30688), .A1(g13484), .A2(g30348) );
  NOR2_X1 NOR2_1793( .ZN(g30689), .A1(g13486), .A2(g30351) );
  NOR2_X1 NOR2_1794( .ZN(g30690), .A1(g13489), .A2(g30352) );
  NOR2_X1 NOR2_1795( .ZN(g30691), .A1(g13491), .A2(g30355) );
  NOR2_X1 NOR2_1796( .ZN(g30692), .A1(g13498), .A2(g30361) );
  NOR2_X1 NOR2_1797( .ZN(g30693), .A1(g13503), .A2(g30364) );
  NOR2_X1 NOR2_1798( .ZN(g30694), .A1(g13505), .A2(g30367) );
  NOR2_X1 NOR2_1799( .ZN(g30695), .A1(g13515), .A2(g30374) );
  NOR2_X1 NOR2_1800( .ZN(g30699), .A1(g13914), .A2(g30387) );
  NOR2_X1 NOR2_1801( .ZN(g30700), .A1(g13952), .A2(g30388) );
  NOR2_X1 NOR2_1802( .ZN(g30701), .A1(g13970), .A2(g30389) );
  NOR2_X1 NOR2_1803( .ZN(g30702), .A1(g14006), .A2(g30390) );
  NOR2_X1 NOR2_1804( .ZN(g30703), .A1(g14022), .A2(g30391) );
  NOR2_X1 NOR2_1805( .ZN(g30704), .A1(g14040), .A2(g30392) );
  NOR2_X1 NOR2_1806( .ZN(g30705), .A1(g14097), .A2(g30393) );
  NOR2_X1 NOR2_1807( .ZN(g30706), .A1(g14113), .A2(g30394) );
  NOR2_X1 NOR2_1808( .ZN(g30707), .A1(g14131), .A2(g30395) );
  NOR2_X1 NOR2_1809( .ZN(g30708), .A1(g14212), .A2(g30396) );
  NOR2_X1 NOR2_1810( .ZN(g30709), .A1(g14228), .A2(g30397) );
  NOR2_X1 NOR2_1811( .ZN(g30780), .A1(g30625), .A2(g22387) );
  NOR2_X1 NOR2_1812( .ZN(g30783), .A1(g30618), .A2(g22387) );
  NOR2_X1 NOR2_1813( .ZN(g30785), .A1(g30618), .A2(g22387) );
  NOR2_X1 NOR2_1814( .ZN(g30786), .A1(g30625), .A2(g22387) );
  NOR2_X1 NOR2_1815( .ZN(g30787), .A1(g30594), .A2(g22387) );
  NOR2_X1 NOR2_1816( .ZN(g30788), .A1(g30602), .A2(g22387) );
  NOR2_X1 NOR2_1817( .ZN(g30789), .A1(g30575), .A2(g22387) );
  NOR2_X1 NOR2_1818( .ZN(g30790), .A1(g30575), .A2(g22387) );
  NOR2_X1 NOR2_1819( .ZN(g30796), .A1(g16069), .A2(g30696) );
  NOR2_X1 NOR2_1820( .ZN(g30798), .A1(g16134), .A2(g30697) );
  NOR2_X1 NOR2_1821( .ZN(g30801), .A1(g16237), .A2(g30698) );
  NOR2_X1 NOR2_1822( .ZN(g30929), .A1(g30728), .A2(g30736) );
  NOR2_X1 NOR2_1823( .ZN(g30930), .A1(g30735), .A2(g30744) );
  NOR2_X1 NOR2_1824( .ZN(g30931), .A1(g30743), .A2(g30750) );
  NOR2_X2 NOR2_1825( .ZN(g30932), .A1(g30754), .A2(g30757) );
  NOR2_X2 NOR2_1826( .ZN(g30933), .A1(g30755), .A2(g30758) );
  NOR2_X2 NOR2_1827( .ZN(g30934), .A1(g30759), .A2(g30761) );
  NOR2_X1 NOR2_1828( .ZN(g30935), .A1(g30760), .A2(g30762) );
  NOR2_X1 NOR2_1829( .ZN(g30936), .A1(g30763), .A2(g30764) );
  NOR2_X1 NOR2_1830( .ZN(g30954), .A1(g30916), .A2(g30944) );
  NOR2_X1 NOR2_1831( .ZN(g30955), .A1(g30918), .A2(g30945) );
  NOR2_X1 NOR2_1832( .ZN(g30956), .A1(g30919), .A2(g30946) );
  NOR2_X1 NOR2_1833( .ZN(g30957), .A1(g30920), .A2(g30947) );
  NOR2_X1 NOR2_1834( .ZN(g30958), .A1(g30922), .A2(g30948) );
  NOR2_X1 NOR2_1835( .ZN(g30959), .A1(g30923), .A2(g30949) );
  NOR2_X1 NOR2_1836( .ZN(g30960), .A1(g30924), .A2(g30950) );
  NOR2_X1 NOR2_1837( .ZN(g30961), .A1(g30925), .A2(g30951) );
  NOR3_X2 NOR3_420( .ZN(g30970), .A1(g30917), .A2(g30921), .A3(g30953) );

endmodule
