// Verilog
// c3540
// Ninputs 50
// Noutputs 22
// NtotalGates 1669
// BUFF1 223
// NOT1 490
// OR2 35
// AND2 410
// NAND2 274
// NAND3 17
// AND3 76
// NOR2 25
// AND4 10
// NAND4 7
// OR3 56
// NOR3 27
// AND5 2
// NOR8 16
// OR4 1

module c3540(N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,
  N137,N143,N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,
  N270,N274,N283,N294,N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,N1713,N1947,N3195,N3833,
  N3987,N4028,N4145,N4589,N4667,N4815,N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,N5360,N5361);
input N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
  N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
  N303,N311,N317,N322,N326,N329,N330,N343,N349,N350;
output N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
  N5360,N5361;

  wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,N715,N724,N727,N736,N740,N749,
    N753,N763,N768,N769,N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,N825,N829,
    N832,N835,N836,N839,N842,N845,N848,N851,N854,N858,N861,N864,N867,N870,N874,N877,
    N880,N883,N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,N916,N917,N920,N923,
    N926,N929,N932,N935,N938,N941,N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,
    N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,
    N1261,N1262,N1263,N1264,N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,N1315,N1322,
    N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,
    N1351,N1352,N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
    N1409,N1426,N1427,N1452,N1459,N1460,N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,
    N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,N1508,N1509,N1510,N1511,N1512,N1520,
    N1562,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
    N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,
    N1670,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,N1694,N1714,N1715,N1718,
    N1721,N1722,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,
    N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,
    N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,N1824,N1833,
    N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,
    N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,N1878,N1879,N1880,N1883,
    N1884,N1885,N1888,N1889,N1890,N1893,N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,
    N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,
    N1960,N1961,N1966,N1981,N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,N2024,N2025,
    N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,
    N2068,N2073,N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,
    N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
    N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,N2178,N2179,N2180,N2181,N2183,N2184,
    N2185,N2188,N2191,N2194,N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,N2231,N2232,
    N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,
    N2287,N2294,N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,N2331,N2334,N2341,N2342,
    N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,
    N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,N2435,N2436,N2437,N2438,N2439,N2440,
    N2443,N2444,N2445,N2448,N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,N2477,N2478,
    N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,
    N2587,N2596,N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,
    N2643,N2644,N2645,N2646,N2647,N2648,N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,
    N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,N2729,N2730,N2731,N2732,N2733,N2734,
    N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,N2750,N2751,
    N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,
    N2970,N2973,N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,
    N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,
    N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,
    N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,
    N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,
    N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
    N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,
    N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,
    N3108,N3109,N3110,N3111,N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,N3138,N3141,
    N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,
    N3184,N3187,N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,
    N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,
    N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,
    N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,
    N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
    N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,
    N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,
    N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,
    N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,N3390,N3391,
    N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,
    N3410,N3413,N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,N3438,N3439,N3442,N3445,
    N3446,N3447,N3451,N3455,N3458,N3461,N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,
    N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,N3514,N3517,N3520,N3523,N3534,N3535,
    N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,
    N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,
    N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3648,N3651,N3652,N3653,
    N3654,N3657,N3658,N3661,N3662,N3663,N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,
    N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,N3696,N3697,N3700,N3703,N3704,N3705,
    N3706,N3707,N3708,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3731,N3734,
    N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,
    N3789,N3800,N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,N3835,N3838,N3845,N3850,
    N3855,N3858,N3861,N3865,N3868,N3884,N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,
    N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,N3936,N3937,N3940,N3947,N3948,N3950,
    N3953,N3956,N3959,N3962,N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,N4029,N4030,
    N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,
    N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,N4073,N4074,N4075,N4076,
    N4077,N4078,N4079,N4080,N4085,N4086,N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,
    N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,N4122,N4123,N4126,N4127,N4128,N4139,
    N4142,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,N4186,N4189,
    N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,
    N4241,N4242,N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,N4284,N4287,N4291,N4295,
    N4296,N4299,N4303,N4304,N4305,N4310,N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,
    N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,N4359,N4362,N4365,N4368,N4371,N4376,
    N4377,N4387,N4390,N4393,N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,N4447,N4448,
    N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,
    N4496,N4497,N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,N4527,N4528,N4529,N4530,
    N4531,N4534,N4537,N4540,N4545,N4549,N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,
    N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,N4602,N4603,N4608,N4613,N4616,N4619,
    N4623,N4628,N4629,N4630,N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,N4659,N4664,
    N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,
    N4704,N4705,N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,N4730,N4733,N4740,N4743,
    N4747,N4748,N4749,N4750,N4753,N4754,N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,
    N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,N4822,N4823,N4826,N4829,N4830,N4831,
    N4838,N4844,N4847,N4850,N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,N4889,N4895,
    N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,
    N4925,N4926,N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,N4952,N4953,N4954,N4957,
    N4964,N4965,N4968,N4969,N4970,N4973,N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,
    N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,N5039,N5042,N5046,N5050,N5055,N5058,
    N5061,N5066,N5070,N5080,N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,N5117,N5122,
    N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,
    N5183,N5184,N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,N5212,N5215,N5217,N5219,
    N5220,N5221,N5222,N5223,N5224,N5225,N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,
    N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,N5278,N5279,N5283,N5284,N5285,N5286,
    N5289,N5292,N5295,N5298,N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,N5335,N5340,
    N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,N5358,N5359,extra0,
    extra1,extra2,extra3,extra4,extra5,extra6,extra7,extra8,extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,
    extra17,extra18,extra19,extra20,extra21,extra22,extra23,extra24,extra25,extra26,extra27,extra28,extra29,extra30,extra31,extra32,
    extra33,extra34,extra35,extra36,extra37,extra38,extra39,extra40,extra41,extra42,extra43,extra44,extra45,extra46,extra47,extra48,
    extra49;

  BUF_X1 BUFF1_1( .Z(N655), .A(N50) );
  INV_X4 NOT1_2( .ZN(N665), .A(N50) );
  BUF_X1 BUFF1_3( .Z(N670), .A(N58) );
  INV_X4 NOT1_4( .ZN(N679), .A(N58) );
  BUF_X1 BUFF1_5( .Z(N683), .A(N68) );
  INV_X4 NOT1_6( .ZN(N686), .A(N68) );
  BUF_X1 BUFF1_7( .Z(N690), .A(N68) );
  BUF_X1 BUFF1_8( .Z(N699), .A(N77) );
  INV_X4 NOT1_9( .ZN(N702), .A(N77) );
  BUF_X1 BUFF1_10( .Z(N706), .A(N77) );
  BUF_X1 BUFF1_11( .Z(N715), .A(N87) );
  INV_X4 NOT1_12( .ZN(N724), .A(N87) );
  BUF_X1 BUFF1_13( .Z(N727), .A(N97) );
  INV_X1 NOT1_14( .ZN(N736), .A(N97) );
  BUF_X1 BUFF1_15( .Z(N740), .A(N107) );
  INV_X1 NOT1_16( .ZN(N749), .A(N107) );
  BUF_X1 BUFF1_17( .Z(N753), .A(N116) );
  INV_X1 NOT1_18( .ZN(N763), .A(N116) );
  OR2_X1 OR2_19( .ZN(N768), .A1(N257), .A2(N264) );
  INV_X1 NOT1_20( .ZN(N769), .A(N1) );
  BUF_X1 BUFF1_21( .Z(N772), .A(N1) );
  INV_X1 NOT1_22( .ZN(N779), .A(N1) );
  BUF_X1 BUFF1_23( .Z(N782), .A(N13) );
  INV_X1 NOT1_24( .ZN(N786), .A(N13) );
  AND2_X1 AND2_25( .ZN(N793), .A1(N13), .A2(N20) );
  INV_X1 NOT1_26( .ZN(N794), .A(N20) );
  BUF_X1 BUFF1_27( .Z(N798), .A(N20) );
  INV_X1 NOT1_28( .ZN(N803), .A(N20) );
  INV_X1 NOT1_29( .ZN(N820), .A(N33) );
  BUF_X1 BUFF1_30( .Z(N821), .A(N33) );
  INV_X1 NOT1_31( .ZN(N825), .A(N33) );
  AND2_X1 AND2_32( .ZN(N829), .A1(N33), .A2(N41) );
  INV_X1 NOT1_33( .ZN(N832), .A(N41) );
  OR2_X1 OR2_34( .ZN(N835), .A1(N41), .A2(N45) );
  BUF_X1 BUFF1_35( .Z(N836), .A(N45) );
  INV_X1 NOT1_36( .ZN(N839), .A(N45) );
  INV_X1 NOT1_37( .ZN(N842), .A(N50) );
  BUF_X1 BUFF1_38( .Z(N845), .A(N58) );
  INV_X1 NOT1_39( .ZN(N848), .A(N58) );
  BUF_X1 BUFF1_40( .Z(N851), .A(N68) );
  INV_X1 NOT1_41( .ZN(N854), .A(N68) );
  BUF_X1 BUFF1_42( .Z(N858), .A(N87) );
  INV_X1 NOT1_43( .ZN(N861), .A(N87) );
  BUF_X1 BUFF1_44( .Z(N864), .A(N97) );
  INV_X1 NOT1_45( .ZN(N867), .A(N97) );
  INV_X1 NOT1_46( .ZN(N870), .A(N107) );
  BUF_X1 BUFF1_47( .Z(N874), .A(N1) );
  BUF_X1 BUFF1_48( .Z(N877), .A(N68) );
  BUF_X1 BUFF1_49( .Z(N880), .A(N107) );
  INV_X1 NOT1_50( .ZN(N883), .A(N20) );
  BUF_X1 BUFF1_51( .Z(N886), .A(N190) );
  INV_X1 NOT1_52( .ZN(N889), .A(N200) );
  AND2_X1 AND2_53( .ZN(N890), .A1(N20), .A2(N200) );
  NAND2_X1 NAND2_54( .ZN(N891), .A1(N20), .A2(N200) );
  AND2_X1 AND2_55( .ZN(N892), .A1(N20), .A2(N179) );
  INV_X1 NOT1_56( .ZN(N895), .A(N20) );
  OR2_X1 OR2_57( .ZN(N896), .A1(N349), .A2(N33) );
  NAND2_X1 NAND2_58( .ZN(N913), .A1(N1), .A2(N13) );
  NAND3_X1 NAND3_59( .ZN(N914), .A1(N1), .A2(N20), .A3(N33) );
  INV_X1 NOT1_60( .ZN(N915), .A(N20) );
  INV_X1 NOT1_61( .ZN(N916), .A(N33) );
  BUF_X1 BUFF1_62( .Z(N917), .A(N179) );
  INV_X1 NOT1_63( .ZN(N920), .A(N213) );
  BUF_X1 BUFF1_64( .Z(N923), .A(N343) );
  BUF_X1 BUFF1_65( .Z(N926), .A(N226) );
  BUF_X1 BUFF1_66( .Z(N929), .A(N232) );
  BUF_X1 BUFF1_67( .Z(N932), .A(N238) );
  BUF_X1 BUFF1_68( .Z(N935), .A(N244) );
  BUF_X1 BUFF1_69( .Z(N938), .A(N250) );
  BUF_X1 BUFF1_70( .Z(N941), .A(N257) );
  BUF_X1 BUFF1_71( .Z(N944), .A(N264) );
  BUF_X1 BUFF1_72( .Z(N947), .A(N270) );
  BUF_X1 BUFF1_73( .Z(N950), .A(N50) );
  BUF_X1 BUFF1_74( .Z(N953), .A(N58) );
  BUF_X1 BUFF1_75( .Z(N956), .A(N58) );
  BUF_X1 BUFF1_76( .Z(N959), .A(N97) );
  BUF_X1 BUFF1_77( .Z(N962), .A(N97) );
  BUF_X1 BUFF1_78( .Z(N965), .A(N330) );
  AND2_X1 AND2_79( .ZN(N1067), .A1(N250), .A2(N768) );
  OR2_X1 OR2_80( .ZN(N1117), .A1(N820), .A2(N20) );
  OR2_X1 OR2_81( .ZN(N1179), .A1(N895), .A2(N169) );
  INV_X1 NOT1_82( .ZN(N1196), .A(N793) );
  OR2_X1 OR2_83( .ZN(N1197), .A1(N915), .A2(N1) );
  AND2_X1 AND2_84( .ZN(N1202), .A1(N913), .A2(N914) );
  OR2_X1 OR2_85( .ZN(N1219), .A1(N916), .A2(N1) );
  AND3_X1 AND3_86( .ZN(N1250), .A1(N842), .A2(N848), .A3(N854) );
  NAND2_X1 NAND2_87( .ZN(N1251), .A1(N226), .A2(N655) );
  NAND2_X1 NAND2_88( .ZN(N1252), .A1(N232), .A2(N670) );
  NAND2_X1 NAND2_89( .ZN(N1253), .A1(N238), .A2(N690) );
  NAND2_X1 NAND2_90( .ZN(N1254), .A1(N244), .A2(N706) );
  NAND2_X1 NAND2_91( .ZN(N1255), .A1(N250), .A2(N715) );
  NAND2_X1 NAND2_92( .ZN(N1256), .A1(N257), .A2(N727) );
  NAND2_X1 NAND2_93( .ZN(N1257), .A1(N264), .A2(N740) );
  NAND2_X1 NAND2_94( .ZN(N1258), .A1(N270), .A2(N753) );
  INV_X4 NOT1_95( .ZN(N1259), .A(N926) );
  INV_X4 NOT1_96( .ZN(N1260), .A(N929) );
  INV_X4 NOT1_97( .ZN(N1261), .A(N932) );
  INV_X4 NOT1_98( .ZN(N1262), .A(N935) );
  NAND2_X1 NAND2_99( .ZN(N1263), .A1(N679), .A2(N686) );
  NAND2_X1 NAND2_100( .ZN(N1264), .A1(N736), .A2(N749) );
  NAND2_X1 NAND2_101( .ZN(N1267), .A1(N683), .A2(N699) );
  BUF_X1 BUFF1_102( .Z(N1268), .A(N665) );
  INV_X4 NOT1_103( .ZN(N1271), .A(N953) );
  INV_X4 NOT1_104( .ZN(N1272), .A(N959) );
  BUF_X1 BUFF1_105( .Z(N1273), .A(N839) );
  BUF_X1 BUFF1_106( .Z(N1276), .A(N839) );
  BUF_X1 BUFF1_107( .Z(N1279), .A(N782) );
  BUF_X1 BUFF1_108( .Z(N1298), .A(N825) );
  BUF_X1 BUFF1_109( .Z(N1302), .A(N832) );
  AND2_X1 AND2_110( .ZN(N1306), .A1(N779), .A2(N835) );
  AND3_X1 AND3_111( .ZN(N1315), .A1(N779), .A2(N836), .A3(N832) );
  AND2_X1 AND2_112( .ZN(N1322), .A1(N769), .A2(N836) );
  AND3_X1 AND3_113( .ZN(N1325), .A1(N772), .A2(N786), .A3(N798) );
  NAND3_X1 NAND3_114( .ZN(N1328), .A1(N772), .A2(N786), .A3(N798) );
  NAND2_X1 NAND2_115( .ZN(N1331), .A1(N772), .A2(N786) );
  BUF_X1 BUFF1_116( .Z(N1334), .A(N874) );
  NAND3_X1 NAND3_117( .ZN(N1337), .A1(N782), .A2(N794), .A3(N45) );
  NAND3_X1 NAND3_118( .ZN(N1338), .A1(N842), .A2(N848), .A3(N854) );
  INV_X1 NOT1_119( .ZN(N1339), .A(N956) );
  AND3_X1 AND3_120( .ZN(N1340), .A1(N861), .A2(N867), .A3(N870) );
  NAND3_X1 NAND3_121( .ZN(N1343), .A1(N861), .A2(N867), .A3(N870) );
  INV_X1 NOT1_122( .ZN(N1344), .A(N962) );
  INV_X1 NOT1_123( .ZN(N1345), .A(N803) );
  INV_X1 NOT1_124( .ZN(N1346), .A(N803) );
  INV_X1 NOT1_125( .ZN(N1347), .A(N803) );
  INV_X1 NOT1_126( .ZN(N1348), .A(N803) );
  INV_X1 NOT1_127( .ZN(N1349), .A(N803) );
  INV_X1 NOT1_128( .ZN(N1350), .A(N803) );
  INV_X1 NOT1_129( .ZN(N1351), .A(N803) );
  INV_X1 NOT1_130( .ZN(N1352), .A(N803) );
  OR2_X1 OR2_131( .ZN(N1353), .A1(N883), .A2(N886) );
  NOR2_X1 NOR2_132( .ZN(N1358), .A1(N883), .A2(N886) );
  BUF_X1 BUFF1_133( .Z(N1363), .A(N892) );
  INV_X1 NOT1_134( .ZN(N1366), .A(N892) );
  BUF_X1 BUFF1_135( .Z(N1369), .A(N821) );
  BUF_X1 BUFF1_136( .Z(N1384), .A(N825) );
  INV_X1 NOT1_137( .ZN(N1401), .A(N896) );
  INV_X1 NOT1_138( .ZN(N1402), .A(N896) );
  INV_X1 NOT1_139( .ZN(N1403), .A(N896) );
  INV_X1 NOT1_140( .ZN(N1404), .A(N896) );
  INV_X1 NOT1_141( .ZN(N1405), .A(N896) );
  INV_X1 NOT1_142( .ZN(N1406), .A(N896) );
  INV_X1 NOT1_143( .ZN(N1407), .A(N896) );
  INV_X1 NOT1_144( .ZN(N1408), .A(N896) );
  OR2_X1 OR2_145( .ZN(N1409), .A1(N1), .A2(N1196) );
  INV_X4 NOT1_146( .ZN(N1426), .A(N829) );
  INV_X4 NOT1_147( .ZN(N1427), .A(N829) );
  AND3_X1 AND3_148( .ZN(N1452), .A1(N769), .A2(N782), .A3(N794) );
  INV_X4 NOT1_149( .ZN(N1459), .A(N917) );
  INV_X1 NOT1_150( .ZN(N1460), .A(N965) );
  OR2_X1 OR2_151( .ZN(N1461), .A1(N920), .A2(N923) );
  NOR2_X1 NOR2_152( .ZN(N1464), .A1(N920), .A2(N923) );
  INV_X1 NOT1_153( .ZN(N1467), .A(N938) );
  INV_X1 NOT1_154( .ZN(N1468), .A(N941) );
  INV_X1 NOT1_155( .ZN(N1469), .A(N944) );
  INV_X1 NOT1_156( .ZN(N1470), .A(N947) );
  BUF_X1 BUFF1_157( .Z(N1471), .A(N679) );
  INV_X1 NOT1_158( .ZN(N1474), .A(N950) );
  BUF_X1 BUFF1_159( .Z(N1475), .A(N686) );
  BUF_X1 BUFF1_160( .Z(N1478), .A(N702) );
  BUF_X1 BUFF1_161( .Z(N1481), .A(N724) );
  BUF_X1 BUFF1_162( .Z(N1484), .A(N736) );
  BUF_X1 BUFF1_163( .Z(N1487), .A(N749) );
  BUF_X1 BUFF1_164( .Z(N1490), .A(N763) );
  BUF_X1 BUFF1_165( .Z(N1493), .A(N877) );
  BUF_X1 BUFF1_166( .Z(N1496), .A(N877) );
  BUF_X1 BUFF1_167( .Z(N1499), .A(N880) );
  BUF_X1 BUFF1_168( .Z(N1502), .A(N880) );
  NAND2_X1 NAND2_169( .ZN(N1505), .A1(N702), .A2(N1250) );
  AND4_X1 AND4_170( .ZN(N1507), .A1(N1251), .A2(N1252), .A3(N1253), .A4(N1254) );
  AND4_X1 AND4_171( .ZN(N1508), .A1(N1255), .A2(N1256), .A3(N1257), .A4(N1258) );
  NAND2_X1 NAND2_172( .ZN(N1509), .A1(N929), .A2(N1259) );
  NAND2_X1 NAND2_173( .ZN(N1510), .A1(N926), .A2(N1260) );
  NAND2_X1 NAND2_174( .ZN(N1511), .A1(N935), .A2(N1261) );
  NAND2_X1 NAND2_175( .ZN(N1512), .A1(N932), .A2(N1262) );
  AND2_X1 AND2_176( .ZN(N1520), .A1(N655), .A2(N1263) );
  AND2_X1 AND2_177( .ZN(N1562), .A1(N874), .A2(N1337) );
  INV_X1 NOT1_178( .ZN(N1579), .A(N1117) );
  AND2_X1 AND2_179( .ZN(N1580), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_180( .ZN(N1581), .A1(N1338), .A2(N1345) );
  INV_X1 NOT1_181( .ZN(N1582), .A(N1117) );
  AND2_X1 AND2_182( .ZN(N1583), .A1(N803), .A2(N1117) );
  INV_X1 NOT1_183( .ZN(N1584), .A(N1117) );
  AND2_X1 AND2_184( .ZN(N1585), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_185( .ZN(N1586), .A1(N854), .A2(N1347) );
  INV_X1 NOT1_186( .ZN(N1587), .A(N1117) );
  AND2_X1 AND2_187( .ZN(N1588), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_188( .ZN(N1589), .A1(N77), .A2(N1348) );
  INV_X1 NOT1_189( .ZN(N1590), .A(N1117) );
  AND2_X1 AND2_190( .ZN(N1591), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_191( .ZN(N1592), .A1(N1343), .A2(N1349) );
  INV_X1 NOT1_192( .ZN(N1593), .A(N1117) );
  AND2_X1 AND2_193( .ZN(N1594), .A1(N803), .A2(N1117) );
  INV_X1 NOT1_194( .ZN(N1595), .A(N1117) );
  AND2_X1 AND2_195( .ZN(N1596), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_196( .ZN(N1597), .A1(N870), .A2(N1351) );
  INV_X1 NOT1_197( .ZN(N1598), .A(N1117) );
  AND2_X1 AND2_198( .ZN(N1599), .A1(N803), .A2(N1117) );
  AND2_X1 AND2_199( .ZN(N1600), .A1(N116), .A2(N1352) );
  AND2_X1 AND2_200( .ZN(N1643), .A1(N222), .A2(N1401) );
  AND2_X1 AND2_201( .ZN(N1644), .A1(N223), .A2(N1402) );
  AND2_X1 AND2_202( .ZN(N1645), .A1(N226), .A2(N1403) );
  AND2_X1 AND2_203( .ZN(N1646), .A1(N232), .A2(N1404) );
  AND2_X1 AND2_204( .ZN(N1647), .A1(N238), .A2(N1405) );
  AND2_X1 AND2_205( .ZN(N1648), .A1(N244), .A2(N1406) );
  AND2_X1 AND2_206( .ZN(N1649), .A1(N250), .A2(N1407) );
  AND2_X1 AND2_207( .ZN(N1650), .A1(N257), .A2(N1408) );
  AND3_X1 AND3_208( .ZN(N1667), .A1(N1), .A2(N13), .A3(N1426) );
  AND3_X1 AND3_209( .ZN(N1670), .A1(N1), .A2(N13), .A3(N1427) );
  INV_X1 NOT1_210( .ZN(N1673), .A(N1202) );
  INV_X4 NOT1_211( .ZN(N1674), .A(N1202) );
  INV_X4 NOT1_212( .ZN(N1675), .A(N1202) );
  INV_X1 NOT1_213( .ZN(N1676), .A(N1202) );
  INV_X1 NOT1_214( .ZN(N1677), .A(N1202) );
  INV_X1 NOT1_215( .ZN(N1678), .A(N1202) );
  INV_X1 NOT1_216( .ZN(N1679), .A(N1202) );
  INV_X1 NOT1_217( .ZN(N1680), .A(N1202) );
  NAND2_X1 NAND2_218( .ZN(N1691), .A1(N941), .A2(N1467) );
  NAND2_X1 NAND2_219( .ZN(N1692), .A1(N938), .A2(N1468) );
  NAND2_X1 NAND2_220( .ZN(N1693), .A1(N947), .A2(N1469) );
  NAND2_X1 NAND2_221( .ZN(N1694), .A1(N944), .A2(N1470) );
  INV_X1 NOT1_222( .ZN(N1713), .A(N1505) );
  AND2_X1 AND2_223( .ZN(N1714), .A1(N87), .A2(N1264) );
  NAND2_X1 NAND2_224( .ZN(N1715), .A1(N1509), .A2(N1510) );
  NAND2_X1 NAND2_225( .ZN(N1718), .A1(N1511), .A2(N1512) );
  NAND2_X1 NAND2_226( .ZN(N1721), .A1(N1507), .A2(N1508) );
  AND2_X1 AND2_227( .ZN(N1722), .A1(N763), .A2(N1340) );
  NAND2_X1 NAND2_228( .ZN(N1725), .A1(N763), .A2(N1340) );
  INV_X1 NOT1_229( .ZN(N1726), .A(N1268) );
  NAND2_X1 NAND2_230( .ZN(N1727), .A1(N1493), .A2(N1271) );
  INV_X1 NOT1_231( .ZN(N1728), .A(N1493) );
  AND2_X1 AND2_232( .ZN(N1729), .A1(N683), .A2(N1268) );
  NAND2_X1 NAND2_233( .ZN(N1730), .A1(N1499), .A2(N1272) );
  INV_X1 NOT1_234( .ZN(N1731), .A(N1499) );
  NAND2_X1 NAND2_235( .ZN(N1735), .A1(N87), .A2(N1264) );
  INV_X1 NOT1_236( .ZN(N1736), .A(N1273) );
  INV_X1 NOT1_237( .ZN(N1737), .A(N1276) );
  NAND2_X1 NAND2_238( .ZN(N1738), .A1(N1325), .A2(N821) );
  NAND2_X1 NAND2_239( .ZN(N1747), .A1(N1325), .A2(N825) );
  NAND3_X1 NAND3_240( .ZN(N1756), .A1(N772), .A2(N1279), .A3(N798) );
  NAND4_X1 NAND4_241( .ZN(N1761), .A1(N772), .A2(N786), .A3(N798), .A4(N1302) );
  NAND2_X1 NAND2_242( .ZN(N1764), .A1(N1496), .A2(N1339) );
  INV_X1 NOT1_243( .ZN(N1765), .A(N1496) );
  NAND2_X1 NAND2_244( .ZN(N1766), .A1(N1502), .A2(N1344) );
  INV_X1 NOT1_245( .ZN(N1767), .A(N1502) );
  INV_X1 NOT1_246( .ZN(N1768), .A(N1328) );
  INV_X1 NOT1_247( .ZN(N1769), .A(N1334) );
  INV_X1 NOT1_248( .ZN(N1770), .A(N1331) );
  AND2_X1 AND2_249( .ZN(N1787), .A1(N845), .A2(N1579) );
  AND2_X1 AND2_250( .ZN(N1788), .A1(N150), .A2(N1580) );
  AND2_X1 AND2_251( .ZN(N1789), .A1(N851), .A2(N1582) );
  AND2_X1 AND2_252( .ZN(N1790), .A1(N159), .A2(N1583) );
  AND2_X1 AND2_253( .ZN(N1791), .A1(N77), .A2(N1584) );
  AND2_X1 AND2_254( .ZN(N1792), .A1(N50), .A2(N1585) );
  AND2_X1 AND2_255( .ZN(N1793), .A1(N858), .A2(N1587) );
  AND2_X1 AND2_256( .ZN(N1794), .A1(N845), .A2(N1588) );
  AND2_X1 AND2_257( .ZN(N1795), .A1(N864), .A2(N1590) );
  AND2_X1 AND2_258( .ZN(N1796), .A1(N851), .A2(N1591) );
  AND2_X1 AND2_259( .ZN(N1797), .A1(N107), .A2(N1593) );
  AND2_X1 AND2_260( .ZN(N1798), .A1(N77), .A2(N1594) );
  AND2_X1 AND2_261( .ZN(N1799), .A1(N116), .A2(N1595) );
  AND2_X1 AND2_262( .ZN(N1800), .A1(N858), .A2(N1596) );
  AND2_X1 AND2_263( .ZN(N1801), .A1(N283), .A2(N1598) );
  AND2_X1 AND2_264( .ZN(N1802), .A1(N864), .A2(N1599) );
  AND2_X1 AND2_265( .ZN(N1803), .A1(N200), .A2(N1363) );
  AND2_X1 AND2_266( .ZN(N1806), .A1(N889), .A2(N1363) );
  AND2_X1 AND2_267( .ZN(N1809), .A1(N890), .A2(N1366) );
  AND2_X1 AND2_268( .ZN(N1812), .A1(N891), .A2(N1366) );
  NAND2_X1 NAND2_269( .ZN(N1815), .A1(N1298), .A2(N1302) );
  NAND2_X1 NAND2_270( .ZN(N1818), .A1(N821), .A2(N1302) );
  NAND3_X1 NAND3_271( .ZN(N1821), .A1(N772), .A2(N1279), .A3(N1179) );
  NAND3_X1 NAND3_272( .ZN(N1824), .A1(N786), .A2(N794), .A3(N1298) );
  NAND2_X1 NAND2_273( .ZN(N1833), .A1(N786), .A2(N1298) );
  INV_X1 NOT1_274( .ZN(N1842), .A(N1369) );
  INV_X1 NOT1_275( .ZN(N1843), .A(N1369) );
  INV_X1 NOT1_276( .ZN(N1844), .A(N1369) );
  INV_X1 NOT1_277( .ZN(N1845), .A(N1369) );
  INV_X1 NOT1_278( .ZN(N1846), .A(N1369) );
  INV_X1 NOT1_279( .ZN(N1847), .A(N1369) );
  INV_X1 NOT1_280( .ZN(N1848), .A(N1369) );
  INV_X1 NOT1_281( .ZN(N1849), .A(N1384) );
  AND2_X1 AND2_282( .ZN(N1850), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_283( .ZN(N1851), .A(N1384) );
  AND2_X1 AND2_284( .ZN(N1852), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_285( .ZN(N1853), .A(N1384) );
  AND2_X1 AND2_286( .ZN(N1854), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_287( .ZN(N1855), .A(N1384) );
  AND2_X1 AND2_288( .ZN(N1856), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_289( .ZN(N1857), .A(N1384) );
  AND2_X1 AND2_290( .ZN(N1858), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_291( .ZN(N1859), .A(N1384) );
  AND2_X1 AND2_292( .ZN(N1860), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_293( .ZN(N1861), .A(N1384) );
  AND2_X1 AND2_294( .ZN(N1862), .A1(N1384), .A2(N896) );
  INV_X1 NOT1_295( .ZN(N1863), .A(N1384) );
  AND2_X1 AND2_296( .ZN(N1864), .A1(N1384), .A2(N896) );
  AND2_X1 AND2_297( .ZN(N1869), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_298( .ZN(N1870), .A1(N50), .A2(N1409) );
  INV_X1 NOT1_299( .ZN(N1873), .A(N1306) );
  AND2_X1 AND2_300( .ZN(N1874), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_301( .ZN(N1875), .A1(N58), .A2(N1409) );
  INV_X1 NOT1_302( .ZN(N1878), .A(N1306) );
  AND2_X1 AND2_303( .ZN(N1879), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_304( .ZN(N1880), .A1(N68), .A2(N1409) );
  INV_X1 NOT1_305( .ZN(N1883), .A(N1306) );
  AND2_X1 AND2_306( .ZN(N1884), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_307( .ZN(N1885), .A1(N77), .A2(N1409) );
  INV_X1 NOT1_308( .ZN(N1888), .A(N1306) );
  AND2_X1 AND2_309( .ZN(N1889), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_310( .ZN(N1890), .A1(N87), .A2(N1409) );
  INV_X1 NOT1_311( .ZN(N1893), .A(N1322) );
  AND2_X1 AND2_312( .ZN(N1894), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_313( .ZN(N1895), .A1(N97), .A2(N1409) );
  INV_X1 NOT1_314( .ZN(N1898), .A(N1315) );
  AND2_X1 AND2_315( .ZN(N1899), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_316( .ZN(N1900), .A1(N107), .A2(N1409) );
  INV_X1 NOT1_317( .ZN(N1903), .A(N1315) );
  AND2_X1 AND2_318( .ZN(N1904), .A1(N1202), .A2(N1409) );
  NOR2_X1 NOR2_319( .ZN(N1905), .A1(N116), .A2(N1409) );
  INV_X1 NOT1_320( .ZN(N1908), .A(N1315) );
  AND2_X1 AND2_321( .ZN(N1909), .A1(N1452), .A2(N213) );
  NAND2_X1 NAND2_322( .ZN(N1912), .A1(N1452), .A2(N213) );
  AND3_X1 AND3_323( .ZN(N1913), .A1(N1452), .A2(N213), .A3(N343) );
  NAND3_X1 NAND3_324( .ZN(N1917), .A1(N1452), .A2(N213), .A3(N343) );
  AND3_X1 AND3_325( .ZN(N1922), .A1(N1452), .A2(N213), .A3(N343) );
  NAND3_X1 NAND3_326( .ZN(N1926), .A1(N1452), .A2(N213), .A3(N343) );
  BUF_X1 BUFF1_327( .Z(N1930), .A(N1464) );
  NAND2_X1 NAND2_328( .ZN(N1933), .A1(N1691), .A2(N1692) );
  NAND2_X1 NAND2_329( .ZN(N1936), .A1(N1693), .A2(N1694) );
  INV_X1 NOT1_330( .ZN(N1939), .A(N1471) );
  NAND2_X1 NAND2_331( .ZN(N1940), .A1(N1471), .A2(N1474) );
  INV_X1 NOT1_332( .ZN(N1941), .A(N1475) );
  INV_X1 NOT1_333( .ZN(N1942), .A(N1478) );
  INV_X1 NOT1_334( .ZN(N1943), .A(N1481) );
  INV_X1 NOT1_335( .ZN(N1944), .A(N1484) );
  INV_X1 NOT1_336( .ZN(N1945), .A(N1487) );
  INV_X1 NOT1_337( .ZN(N1946), .A(N1490) );
  INV_X1 NOT1_338( .ZN(N1947), .A(N1714) );
  NAND2_X1 NAND2_339( .ZN(N1960), .A1(N953), .A2(N1728) );
  NAND2_X1 NAND2_340( .ZN(N1961), .A1(N959), .A2(N1731) );
  AND2_X1 AND2_341( .ZN(N1966), .A1(N1520), .A2(N1276) );
  NAND2_X1 NAND2_342( .ZN(N1981), .A1(N956), .A2(N1765) );
  NAND2_X1 NAND2_343( .ZN(N1982), .A1(N962), .A2(N1767) );
  AND2_X1 AND2_344( .ZN(N1983), .A1(N1067), .A2(N1768) );
  OR3_X1 OR3_345( .ZN(N1986), .A1(N1581), .A2(N1787), .A3(N1788) );
  OR3_X1 OR3_346( .ZN(N1987), .A1(N1586), .A2(N1791), .A3(N1792) );
  OR3_X1 OR3_347( .ZN(N1988), .A1(N1589), .A2(N1793), .A3(N1794) );
  OR3_X1 OR3_348( .ZN(N1989), .A1(N1592), .A2(N1795), .A3(N1796) );
  OR3_X1 OR3_349( .ZN(N1990), .A1(N1597), .A2(N1799), .A3(N1800) );
  OR3_X1 OR3_350( .ZN(N1991), .A1(N1600), .A2(N1801), .A3(N1802) );
  AND2_X1 AND2_351( .ZN(N2022), .A1(N77), .A2(N1849) );
  AND2_X1 AND2_352( .ZN(N2023), .A1(N223), .A2(N1850) );
  AND2_X1 AND2_353( .ZN(N2024), .A1(N87), .A2(N1851) );
  AND2_X1 AND2_354( .ZN(N2025), .A1(N226), .A2(N1852) );
  AND2_X1 AND2_355( .ZN(N2026), .A1(N97), .A2(N1853) );
  AND2_X1 AND2_356( .ZN(N2027), .A1(N232), .A2(N1854) );
  AND2_X1 AND2_357( .ZN(N2028), .A1(N107), .A2(N1855) );
  AND2_X1 AND2_358( .ZN(N2029), .A1(N238), .A2(N1856) );
  AND2_X1 AND2_359( .ZN(N2030), .A1(N116), .A2(N1857) );
  AND2_X1 AND2_360( .ZN(N2031), .A1(N244), .A2(N1858) );
  AND2_X1 AND2_361( .ZN(N2032), .A1(N283), .A2(N1859) );
  AND2_X1 AND2_362( .ZN(N2033), .A1(N250), .A2(N1860) );
  AND2_X1 AND2_363( .ZN(N2034), .A1(N294), .A2(N1861) );
  AND2_X1 AND2_364( .ZN(N2035), .A1(N257), .A2(N1862) );
  AND2_X1 AND2_365( .ZN(N2036), .A1(N303), .A2(N1863) );
  AND2_X1 AND2_366( .ZN(N2037), .A1(N264), .A2(N1864) );
  BUF_X1 BUFF1_367( .Z(N2038), .A(N1667) );
  INV_X1 NOT1_368( .ZN(N2043), .A(N1667) );
  BUF_X1 BUFF1_369( .Z(N2052), .A(N1670) );
  INV_X1 NOT1_370( .ZN(N2057), .A(N1670) );
  AND3_X1 AND3_371( .ZN(N2068), .A1(N50), .A2(N1197), .A3(N1869) );
  AND3_X1 AND3_372( .ZN(N2073), .A1(N58), .A2(N1197), .A3(N1874) );
  AND3_X1 AND3_373( .ZN(N2078), .A1(N68), .A2(N1197), .A3(N1879) );
  AND3_X1 AND3_374( .ZN(N2083), .A1(N77), .A2(N1197), .A3(N1884) );
  AND3_X1 AND3_375( .ZN(N2088), .A1(N87), .A2(N1219), .A3(N1889) );
  AND3_X1 AND3_376( .ZN(N2093), .A1(N97), .A2(N1219), .A3(N1894) );
  AND3_X1 AND3_377( .ZN(N2098), .A1(N107), .A2(N1219), .A3(N1899) );
  AND3_X1 AND3_378( .ZN(N2103), .A1(N116), .A2(N1219), .A3(N1904) );
  INV_X1 NOT1_379( .ZN(N2121), .A(N1562) );
  INV_X1 NOT1_380( .ZN(N2122), .A(N1562) );
  INV_X1 NOT1_381( .ZN(N2123), .A(N1562) );
  INV_X1 NOT1_382( .ZN(N2124), .A(N1562) );
  INV_X1 NOT1_383( .ZN(N2125), .A(N1562) );
  INV_X1 NOT1_384( .ZN(N2126), .A(N1562) );
  INV_X1 NOT1_385( .ZN(N2127), .A(N1562) );
  INV_X1 NOT1_386( .ZN(N2128), .A(N1562) );
  NAND2_X1 NAND2_387( .ZN(N2133), .A1(N950), .A2(N1939) );
  NAND2_X1 NAND2_388( .ZN(N2134), .A1(N1478), .A2(N1941) );
  NAND2_X1 NAND2_389( .ZN(N2135), .A1(N1475), .A2(N1942) );
  NAND2_X1 NAND2_390( .ZN(N2136), .A1(N1484), .A2(N1943) );
  NAND2_X1 NAND2_391( .ZN(N2137), .A1(N1481), .A2(N1944) );
  NAND2_X1 NAND2_392( .ZN(N2138), .A1(N1490), .A2(N1945) );
  NAND2_X1 NAND2_393( .ZN(N2139), .A1(N1487), .A2(N1946) );
  INV_X1 NOT1_394( .ZN(N2141), .A(N1933) );
  INV_X1 NOT1_395( .ZN(N2142), .A(N1936) );
  INV_X1 NOT1_396( .ZN(N2143), .A(N1738) );
  AND2_X1 AND2_397( .ZN(N2144), .A1(N1738), .A2(N1747) );
  INV_X1 NOT1_398( .ZN(N2145), .A(N1747) );
  NAND2_X1 NAND2_399( .ZN(N2146), .A1(N1727), .A2(N1960) );
  NAND2_X1 NAND2_400( .ZN(N2147), .A1(N1730), .A2(N1961) );
  AND4_X1 AND4_401( .ZN(N2148), .A1(N1722), .A2(N1267), .A3(N665), .A4(N58) );
  INV_X1 NOT1_402( .ZN(N2149), .A(N1738) );
  AND2_X1 AND2_403( .ZN(N2150), .A1(N1738), .A2(N1747) );
  INV_X1 NOT1_404( .ZN(N2151), .A(N1747) );
  INV_X1 NOT1_405( .ZN(N2152), .A(N1738) );
  INV_X1 NOT1_406( .ZN(N2153), .A(N1747) );
  AND2_X1 AND2_407( .ZN(N2154), .A1(N1738), .A2(N1747) );
  INV_X1 NOT1_408( .ZN(N2155), .A(N1738) );
  INV_X1 NOT1_409( .ZN(N2156), .A(N1747) );
  AND2_X1 AND2_410( .ZN(N2157), .A1(N1738), .A2(N1747) );
  BUF_X1 BUFF1_411( .Z(N2158), .A(N1761) );
  BUF_X1 BUFF1_412( .Z(N2175), .A(N1761) );
  NAND2_X1 NAND2_413( .ZN(N2178), .A1(N1764), .A2(N1981) );
  NAND2_X1 NAND2_414( .ZN(N2179), .A1(N1766), .A2(N1982) );
  INV_X1 NOT1_415( .ZN(N2180), .A(N1756) );
  AND2_X1 AND2_416( .ZN(N2181), .A1(N1756), .A2(N1328) );
  INV_X1 NOT1_417( .ZN(N2183), .A(N1756) );
  AND2_X1 AND2_418( .ZN(N2184), .A1(N1331), .A2(N1756) );
  NAND2_X1 NAND2_419( .ZN(N2185), .A1(N1358), .A2(N1812) );
  NAND2_X1 NAND2_420( .ZN(N2188), .A1(N1358), .A2(N1809) );
  NAND2_X1 NAND2_421( .ZN(N2191), .A1(N1353), .A2(N1812) );
  NAND2_X1 NAND2_422( .ZN(N2194), .A1(N1353), .A2(N1809) );
  NAND2_X1 NAND2_423( .ZN(N2197), .A1(N1358), .A2(N1806) );
  NAND2_X1 NAND2_424( .ZN(N2200), .A1(N1358), .A2(N1803) );
  NAND2_X1 NAND2_425( .ZN(N2203), .A1(N1353), .A2(N1806) );
  NAND2_X1 NAND2_426( .ZN(N2206), .A1(N1353), .A2(N1803) );
  INV_X1 NOT1_427( .ZN(N2209), .A(N1815) );
  INV_X1 NOT1_428( .ZN(N2210), .A(N1818) );
  AND2_X1 AND2_429( .ZN(N2211), .A1(N1815), .A2(N1818) );
  BUF_X1 BUFF1_430( .Z(N2212), .A(N1821) );
  BUF_X1 BUFF1_431( .Z(N2221), .A(N1821) );
  INV_X1 NOT1_432( .ZN(N2230), .A(N1833) );
  INV_X1 NOT1_433( .ZN(N2231), .A(N1833) );
  INV_X1 NOT1_434( .ZN(N2232), .A(N1833) );
  INV_X1 NOT1_435( .ZN(N2233), .A(N1833) );
  INV_X1 NOT1_436( .ZN(N2234), .A(N1824) );
  INV_X1 NOT1_437( .ZN(N2235), .A(N1824) );
  INV_X1 NOT1_438( .ZN(N2236), .A(N1824) );
  INV_X1 NOT1_439( .ZN(N2237), .A(N1824) );
  OR3_X1 OR3_440( .ZN(N2238), .A1(N2022), .A2(N1643), .A3(N2023) );
  OR3_X1 OR3_441( .ZN(N2239), .A1(N2024), .A2(N1644), .A3(N2025) );
  OR3_X1 OR3_442( .ZN(N2240), .A1(N2026), .A2(N1645), .A3(N2027) );
  OR3_X1 OR3_443( .ZN(N2241), .A1(N2028), .A2(N1646), .A3(N2029) );
  OR3_X1 OR3_444( .ZN(N2242), .A1(N2030), .A2(N1647), .A3(N2031) );
  OR3_X1 OR3_445( .ZN(N2243), .A1(N2032), .A2(N1648), .A3(N2033) );
  OR3_X1 OR3_446( .ZN(N2244), .A1(N2034), .A2(N1649), .A3(N2035) );
  OR3_X1 OR3_447( .ZN(N2245), .A1(N2036), .A2(N1650), .A3(N2037) );
  AND2_X1 AND2_448( .ZN(N2270), .A1(N1986), .A2(N1673) );
  AND2_X1 AND2_449( .ZN(N2277), .A1(N1987), .A2(N1675) );
  AND2_X1 AND2_450( .ZN(N2282), .A1(N1988), .A2(N1676) );
  AND2_X1 AND2_451( .ZN(N2287), .A1(N1989), .A2(N1677) );
  AND2_X1 AND2_452( .ZN(N2294), .A1(N1990), .A2(N1679) );
  AND2_X1 AND2_453( .ZN(N2299), .A1(N1991), .A2(N1680) );
  BUF_X1 BUFF1_454( .Z(N2304), .A(N1917) );
  AND2_X1 AND2_455( .ZN(N2307), .A1(N1930), .A2(N350) );
  NAND2_X1 NAND2_456( .ZN(N2310), .A1(N1930), .A2(N350) );
  BUF_X1 BUFF1_457( .Z(N2313), .A(N1715) );
  BUF_X1 BUFF1_458( .Z(N2316), .A(N1718) );
  BUF_X1 BUFF1_459( .Z(N2319), .A(N1715) );
  BUF_X1 BUFF1_460( .Z(N2322), .A(N1718) );
  NAND2_X1 NAND2_461( .ZN(N2325), .A1(N1940), .A2(N2133) );
  NAND2_X1 NAND2_462( .ZN(N2328), .A1(N2134), .A2(N2135) );
  NAND2_X1 NAND2_463( .ZN(N2331), .A1(N2136), .A2(N2137) );
  NAND2_X1 NAND2_464( .ZN(N2334), .A1(N2138), .A2(N2139) );
  NAND2_X1 NAND2_465( .ZN(N2341), .A1(N1936), .A2(N2141) );
  NAND2_X1 NAND2_466( .ZN(N2342), .A1(N1933), .A2(N2142) );
  AND2_X1 AND2_467( .ZN(N2347), .A1(N724), .A2(N2144) );
  AND3_X1 AND3_468( .ZN(N2348), .A1(N2146), .A2(N699), .A3(N1726) );
  AND2_X1 AND2_469( .ZN(N2349), .A1(N753), .A2(N2147) );
  AND2_X1 AND2_470( .ZN(N2350), .A1(N2148), .A2(N1273) );
  AND2_X1 AND2_471( .ZN(N2351), .A1(N736), .A2(N2150) );
  AND2_X1 AND2_472( .ZN(N2352), .A1(N1735), .A2(N2153) );
  AND2_X1 AND2_473( .ZN(N2353), .A1(N763), .A2(N2154) );
  AND2_X1 AND2_474( .ZN(N2354), .A1(N1725), .A2(N2156) );
  AND2_X1 AND2_475( .ZN(N2355), .A1(N749), .A2(N2157) );
  INV_X1 NOT1_476( .ZN(N2374), .A(N2178) );
  INV_X1 NOT1_477( .ZN(N2375), .A(N2179) );
  AND2_X1 AND2_478( .ZN(N2376), .A1(N1520), .A2(N2180) );
  AND2_X1 AND2_479( .ZN(N2379), .A1(N1721), .A2(N2181) );
  AND2_X1 AND2_480( .ZN(N2398), .A1(N665), .A2(N2211) );
  AND3_X1 AND3_481( .ZN(N2417), .A1(N2057), .A2(N226), .A3(N1873) );
  AND3_X1 AND3_482( .ZN(N2418), .A1(N2057), .A2(N274), .A3(N1306) );
  AND2_X1 AND2_483( .ZN(N2419), .A1(N2052), .A2(N2238) );
  AND3_X1 AND3_484( .ZN(N2420), .A1(N2057), .A2(N232), .A3(N1878) );
  AND3_X1 AND3_485( .ZN(N2421), .A1(N2057), .A2(N274), .A3(N1306) );
  AND2_X1 AND2_486( .ZN(N2422), .A1(N2052), .A2(N2239) );
  AND3_X1 AND3_487( .ZN(N2425), .A1(N2057), .A2(N238), .A3(N1883) );
  AND3_X1 AND3_488( .ZN(N2426), .A1(N2057), .A2(N274), .A3(N1306) );
  AND2_X1 AND2_489( .ZN(N2427), .A1(N2052), .A2(N2240) );
  AND3_X1 AND3_490( .ZN(N2430), .A1(N2057), .A2(N244), .A3(N1888) );
  AND3_X1 AND3_491( .ZN(N2431), .A1(N2057), .A2(N274), .A3(N1306) );
  AND2_X1 AND2_492( .ZN(N2432), .A1(N2052), .A2(N2241) );
  AND3_X1 AND3_493( .ZN(N2435), .A1(N2043), .A2(N250), .A3(N1893) );
  AND3_X1 AND3_494( .ZN(N2436), .A1(N2043), .A2(N274), .A3(N1322) );
  AND2_X1 AND2_495( .ZN(N2437), .A1(N2038), .A2(N2242) );
  AND3_X1 AND3_496( .ZN(N2438), .A1(N2043), .A2(N257), .A3(N1898) );
  AND3_X1 AND3_497( .ZN(N2439), .A1(N2043), .A2(N274), .A3(N1315) );
  AND2_X1 AND2_498( .ZN(N2440), .A1(N2038), .A2(N2243) );
  AND3_X1 AND3_499( .ZN(N2443), .A1(N2043), .A2(N264), .A3(N1903) );
  AND3_X1 AND3_500( .ZN(N2444), .A1(N2043), .A2(N274), .A3(N1315) );
  AND2_X1 AND2_501( .ZN(N2445), .A1(N2038), .A2(N2244) );
  AND3_X1 AND3_502( .ZN(N2448), .A1(N2043), .A2(N270), .A3(N1908) );
  AND3_X1 AND3_503( .ZN(N2449), .A1(N2043), .A2(N274), .A3(N1315) );
  AND2_X1 AND2_504( .ZN(N2450), .A1(N2038), .A2(N2245) );
  INV_X1 NOT1_505( .ZN(N2467), .A(N2313) );
  INV_X1 NOT1_506( .ZN(N2468), .A(N2316) );
  INV_X1 NOT1_507( .ZN(N2469), .A(N2319) );
  INV_X1 NOT1_508( .ZN(N2470), .A(N2322) );
  NAND2_X1 NAND2_509( .ZN(N2471), .A1(N2341), .A2(N2342) );
  INV_X1 NOT1_510( .ZN(N2474), .A(N2325) );
  INV_X1 NOT1_511( .ZN(N2475), .A(N2328) );
  INV_X1 NOT1_512( .ZN(N2476), .A(N2331) );
  INV_X1 NOT1_513( .ZN(N2477), .A(N2334) );
  OR2_X1 OR2_514( .ZN(N2478), .A1(N2348), .A2(N1729) );
  INV_X1 NOT1_515( .ZN(N2481), .A(N2175) );
  AND2_X1 AND2_516( .ZN(N2482), .A1(N2175), .A2(N1334) );
  AND2_X1 AND2_517( .ZN(N2483), .A1(N2349), .A2(N2183) );
  AND2_X1 AND2_518( .ZN(N2486), .A1(N2374), .A2(N1346) );
  AND2_X1 AND2_519( .ZN(N2487), .A1(N2375), .A2(N1350) );
  BUF_X1 BUFF1_520( .Z(N2488), .A(N2185) );
  BUF_X1 BUFF1_521( .Z(N2497), .A(N2188) );
  BUF_X1 BUFF1_522( .Z(N2506), .A(N2191) );
  BUF_X1 BUFF1_523( .Z(N2515), .A(N2194) );
  BUF_X1 BUFF1_524( .Z(N2524), .A(N2197) );
  BUF_X1 BUFF1_525( .Z(N2533), .A(N2200) );
  BUF_X1 BUFF1_526( .Z(N2542), .A(N2203) );
  BUF_X1 BUFF1_527( .Z(N2551), .A(N2206) );
  BUF_X1 BUFF1_528( .Z(N2560), .A(N2185) );
  BUF_X1 BUFF1_529( .Z(N2569), .A(N2188) );
  BUF_X1 BUFF1_530( .Z(N2578), .A(N2191) );
  BUF_X1 BUFF1_531( .Z(N2587), .A(N2194) );
  BUF_X1 BUFF1_532( .Z(N2596), .A(N2197) );
  BUF_X1 BUFF1_533( .Z(N2605), .A(N2200) );
  BUF_X1 BUFF1_534( .Z(N2614), .A(N2203) );
  BUF_X1 BUFF1_535( .Z(N2623), .A(N2206) );
  INV_X1 NOT1_536( .ZN(N2632), .A(N2212) );
  AND2_X1 AND2_537( .ZN(N2633), .A1(N2212), .A2(N1833) );
  INV_X1 NOT1_538( .ZN(N2634), .A(N2212) );
  AND2_X1 AND2_539( .ZN(N2635), .A1(N2212), .A2(N1833) );
  INV_X1 NOT1_540( .ZN(N2636), .A(N2212) );
  AND2_X1 AND2_541( .ZN(N2637), .A1(N2212), .A2(N1833) );
  INV_X1 NOT1_542( .ZN(N2638), .A(N2212) );
  AND2_X1 AND2_543( .ZN(N2639), .A1(N2212), .A2(N1833) );
  INV_X1 NOT1_544( .ZN(N2640), .A(N2221) );
  AND2_X1 AND2_545( .ZN(N2641), .A1(N2221), .A2(N1824) );
  INV_X1 NOT1_546( .ZN(N2642), .A(N2221) );
  AND2_X1 AND2_547( .ZN(N2643), .A1(N2221), .A2(N1824) );
  INV_X1 NOT1_548( .ZN(N2644), .A(N2221) );
  AND2_X1 AND2_549( .ZN(N2645), .A1(N2221), .A2(N1824) );
  INV_X1 NOT1_550( .ZN(N2646), .A(N2221) );
  AND2_X1 AND2_551( .ZN(N2647), .A1(N2221), .A2(N1824) );
  OR3_X1 OR3_552( .ZN(N2648), .A1(N2270), .A2(N1870), .A3(N2068) );
  NOR3_X1 NOR3_553( .ZN(N2652), .A1(N2270), .A2(N1870), .A3(N2068) );
  OR3_X1 OR3_554( .ZN(N2656), .A1(N2417), .A2(N2418), .A3(N2419) );
  OR3_X1 OR3_555( .ZN(N2659), .A1(N2420), .A2(N2421), .A3(N2422) );
  OR3_X1 OR3_556( .ZN(N2662), .A1(N2277), .A2(N1880), .A3(N2078) );
  NOR3_X1 NOR3_557( .ZN(N2666), .A1(N2277), .A2(N1880), .A3(N2078) );
  OR3_X1 OR3_558( .ZN(N2670), .A1(N2425), .A2(N2426), .A3(N2427) );
  OR3_X1 OR3_559( .ZN(N2673), .A1(N2282), .A2(N1885), .A3(N2083) );
  NOR3_X1 NOR3_560( .ZN(N2677), .A1(N2282), .A2(N1885), .A3(N2083) );
  OR3_X1 OR3_561( .ZN(N2681), .A1(N2430), .A2(N2431), .A3(N2432) );
  OR3_X1 OR3_562( .ZN(N2684), .A1(N2287), .A2(N1890), .A3(N2088) );
  NOR3_X1 NOR3_563( .ZN(N2688), .A1(N2287), .A2(N1890), .A3(N2088) );
  OR3_X1 OR3_564( .ZN(N2692), .A1(N2435), .A2(N2436), .A3(N2437) );
  OR3_X1 OR3_565( .ZN(N2697), .A1(N2438), .A2(N2439), .A3(N2440) );
  OR3_X1 OR3_566( .ZN(N2702), .A1(N2294), .A2(N1900), .A3(N2098) );
  NOR3_X1 NOR3_567( .ZN(N2706), .A1(N2294), .A2(N1900), .A3(N2098) );
  OR3_X1 OR3_568( .ZN(N2710), .A1(N2443), .A2(N2444), .A3(N2445) );
  OR3_X1 OR3_569( .ZN(N2715), .A1(N2299), .A2(N1905), .A3(N2103) );
  NOR3_X1 NOR3_570( .ZN(N2719), .A1(N2299), .A2(N1905), .A3(N2103) );
  OR3_X1 OR3_571( .ZN(N2723), .A1(N2448), .A2(N2449), .A3(N2450) );
  INV_X1 NOT1_572( .ZN(N2728), .A(N2304) );
  INV_X1 NOT1_573( .ZN(N2729), .A(N2158) );
  AND2_X1 AND2_574( .ZN(N2730), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_575( .ZN(N2731), .A(N2158) );
  AND2_X1 AND2_576( .ZN(N2732), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_577( .ZN(N2733), .A(N2158) );
  AND2_X1 AND2_578( .ZN(N2734), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_579( .ZN(N2735), .A(N2158) );
  AND2_X1 AND2_580( .ZN(N2736), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_581( .ZN(N2737), .A(N2158) );
  AND2_X1 AND2_582( .ZN(N2738), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_583( .ZN(N2739), .A(N2158) );
  AND2_X1 AND2_584( .ZN(N2740), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_585( .ZN(N2741), .A(N2158) );
  AND2_X1 AND2_586( .ZN(N2742), .A1(N1562), .A2(N2158) );
  INV_X1 NOT1_587( .ZN(N2743), .A(N2158) );
  AND2_X1 AND2_588( .ZN(N2744), .A1(N1562), .A2(N2158) );
  OR3_X1 OR3_589( .ZN(N2745), .A1(N2376), .A2(N1983), .A3(N2379) );
  NOR3_X1 NOR3_590( .ZN(N2746), .A1(N2376), .A2(N1983), .A3(N2379) );
  NAND2_X1 NAND2_591( .ZN(N2748), .A1(N2316), .A2(N2467) );
  NAND2_X1 NAND2_592( .ZN(N2749), .A1(N2313), .A2(N2468) );
  NAND2_X1 NAND2_593( .ZN(N2750), .A1(N2322), .A2(N2469) );
  NAND2_X1 NAND2_594( .ZN(N2751), .A1(N2319), .A2(N2470) );
  NAND2_X1 NAND2_595( .ZN(N2754), .A1(N2328), .A2(N2474) );
  NAND2_X1 NAND2_596( .ZN(N2755), .A1(N2325), .A2(N2475) );
  NAND2_X1 NAND2_597( .ZN(N2756), .A1(N2334), .A2(N2476) );
  NAND2_X1 NAND2_598( .ZN(N2757), .A1(N2331), .A2(N2477) );
  AND2_X1 AND2_599( .ZN(N2758), .A1(N1520), .A2(N2481) );
  AND2_X1 AND2_600( .ZN(N2761), .A1(N1722), .A2(N2482) );
  AND2_X1 AND2_601( .ZN(N2764), .A1(N2478), .A2(N1770) );
  OR3_X1 OR3_602( .ZN(N2768), .A1(N2486), .A2(N1789), .A3(N1790) );
  OR3_X1 OR3_603( .ZN(N2769), .A1(N2487), .A2(N1797), .A3(N1798) );
  AND2_X1 AND2_604( .ZN(N2898), .A1(N665), .A2(N2633) );
  AND2_X1 AND2_605( .ZN(N2899), .A1(N679), .A2(N2635) );
  AND2_X1 AND2_606( .ZN(N2900), .A1(N686), .A2(N2637) );
  AND2_X1 AND2_607( .ZN(N2901), .A1(N702), .A2(N2639) );
  INV_X1 NOT1_608( .ZN(N2962), .A(N2746) );
  NAND2_X1 NAND2_609( .ZN(N2966), .A1(N2748), .A2(N2749) );
  NAND2_X1 NAND2_610( .ZN(N2967), .A1(N2750), .A2(N2751) );
  BUF_X1 BUFF1_611( .Z(N2970), .A(N2471) );
  NAND2_X1 NAND2_612( .ZN(N2973), .A1(N2754), .A2(N2755) );
  NAND2_X1 NAND2_613( .ZN(N2977), .A1(N2756), .A2(N2757) );
  AND2_X1 AND2_614( .ZN(N2980), .A1(N2471), .A2(N2143) );
  INV_X1 NOT1_615( .ZN(N2984), .A(N2488) );
  INV_X1 NOT1_616( .ZN(N2985), .A(N2497) );
  INV_X1 NOT1_617( .ZN(N2986), .A(N2506) );
  INV_X1 NOT1_618( .ZN(N2987), .A(N2515) );
  INV_X1 NOT1_619( .ZN(N2988), .A(N2524) );
  INV_X1 NOT1_620( .ZN(N2989), .A(N2533) );
  INV_X1 NOT1_621( .ZN(N2990), .A(N2542) );
  INV_X1 NOT1_622( .ZN(N2991), .A(N2551) );
  INV_X1 NOT1_623( .ZN(N2992), .A(N2488) );
  INV_X1 NOT1_624( .ZN(N2993), .A(N2497) );
  INV_X1 NOT1_625( .ZN(N2994), .A(N2506) );
  INV_X1 NOT1_626( .ZN(N2995), .A(N2515) );
  INV_X1 NOT1_627( .ZN(N2996), .A(N2524) );
  INV_X1 NOT1_628( .ZN(N2997), .A(N2533) );
  INV_X1 NOT1_629( .ZN(N2998), .A(N2542) );
  INV_X1 NOT1_630( .ZN(N2999), .A(N2551) );
  INV_X1 NOT1_631( .ZN(N3000), .A(N2488) );
  INV_X1 NOT1_632( .ZN(N3001), .A(N2497) );
  INV_X1 NOT1_633( .ZN(N3002), .A(N2506) );
  INV_X1 NOT1_634( .ZN(N3003), .A(N2515) );
  INV_X1 NOT1_635( .ZN(N3004), .A(N2524) );
  INV_X1 NOT1_636( .ZN(N3005), .A(N2533) );
  INV_X1 NOT1_637( .ZN(N3006), .A(N2542) );
  INV_X1 NOT1_638( .ZN(N3007), .A(N2551) );
  INV_X1 NOT1_639( .ZN(N3008), .A(N2488) );
  INV_X1 NOT1_640( .ZN(N3009), .A(N2497) );
  INV_X1 NOT1_641( .ZN(N3010), .A(N2506) );
  INV_X1 NOT1_642( .ZN(N3011), .A(N2515) );
  INV_X1 NOT1_643( .ZN(N3012), .A(N2524) );
  INV_X1 NOT1_644( .ZN(N3013), .A(N2533) );
  INV_X1 NOT1_645( .ZN(N3014), .A(N2542) );
  INV_X1 NOT1_646( .ZN(N3015), .A(N2551) );
  INV_X1 NOT1_647( .ZN(N3016), .A(N2488) );
  INV_X1 NOT1_648( .ZN(N3017), .A(N2497) );
  INV_X1 NOT1_649( .ZN(N3018), .A(N2506) );
  INV_X1 NOT1_650( .ZN(N3019), .A(N2515) );
  INV_X1 NOT1_651( .ZN(N3020), .A(N2524) );
  INV_X1 NOT1_652( .ZN(N3021), .A(N2533) );
  INV_X1 NOT1_653( .ZN(N3022), .A(N2542) );
  INV_X1 NOT1_654( .ZN(N3023), .A(N2551) );
  INV_X1 NOT1_655( .ZN(N3024), .A(N2488) );
  INV_X1 NOT1_656( .ZN(N3025), .A(N2497) );
  INV_X1 NOT1_657( .ZN(N3026), .A(N2506) );
  INV_X1 NOT1_658( .ZN(N3027), .A(N2515) );
  INV_X1 NOT1_659( .ZN(N3028), .A(N2524) );
  INV_X1 NOT1_660( .ZN(N3029), .A(N2533) );
  INV_X1 NOT1_661( .ZN(N3030), .A(N2542) );
  INV_X1 NOT1_662( .ZN(N3031), .A(N2551) );
  INV_X1 NOT1_663( .ZN(N3032), .A(N2488) );
  INV_X1 NOT1_664( .ZN(N3033), .A(N2497) );
  INV_X1 NOT1_665( .ZN(N3034), .A(N2506) );
  INV_X1 NOT1_666( .ZN(N3035), .A(N2515) );
  INV_X1 NOT1_667( .ZN(N3036), .A(N2524) );
  INV_X1 NOT1_668( .ZN(N3037), .A(N2533) );
  INV_X1 NOT1_669( .ZN(N3038), .A(N2542) );
  INV_X1 NOT1_670( .ZN(N3039), .A(N2551) );
  INV_X1 NOT1_671( .ZN(N3040), .A(N2488) );
  INV_X1 NOT1_672( .ZN(N3041), .A(N2497) );
  INV_X1 NOT1_673( .ZN(N3042), .A(N2506) );
  INV_X1 NOT1_674( .ZN(N3043), .A(N2515) );
  INV_X1 NOT1_675( .ZN(N3044), .A(N2524) );
  INV_X1 NOT1_676( .ZN(N3045), .A(N2533) );
  INV_X1 NOT1_677( .ZN(N3046), .A(N2542) );
  INV_X1 NOT1_678( .ZN(N3047), .A(N2551) );
  INV_X1 NOT1_679( .ZN(N3048), .A(N2560) );
  INV_X1 NOT1_680( .ZN(N3049), .A(N2569) );
  INV_X1 NOT1_681( .ZN(N3050), .A(N2578) );
  INV_X1 NOT1_682( .ZN(N3051), .A(N2587) );
  INV_X1 NOT1_683( .ZN(N3052), .A(N2596) );
  INV_X1 NOT1_684( .ZN(N3053), .A(N2605) );
  INV_X1 NOT1_685( .ZN(N3054), .A(N2614) );
  INV_X1 NOT1_686( .ZN(N3055), .A(N2623) );
  INV_X1 NOT1_687( .ZN(N3056), .A(N2560) );
  INV_X1 NOT1_688( .ZN(N3057), .A(N2569) );
  INV_X1 NOT1_689( .ZN(N3058), .A(N2578) );
  INV_X1 NOT1_690( .ZN(N3059), .A(N2587) );
  INV_X1 NOT1_691( .ZN(N3060), .A(N2596) );
  INV_X1 NOT1_692( .ZN(N3061), .A(N2605) );
  INV_X1 NOT1_693( .ZN(N3062), .A(N2614) );
  INV_X1 NOT1_694( .ZN(N3063), .A(N2623) );
  INV_X1 NOT1_695( .ZN(N3064), .A(N2560) );
  INV_X1 NOT1_696( .ZN(N3065), .A(N2569) );
  INV_X1 NOT1_697( .ZN(N3066), .A(N2578) );
  INV_X1 NOT1_698( .ZN(N3067), .A(N2587) );
  INV_X1 NOT1_699( .ZN(N3068), .A(N2596) );
  INV_X1 NOT1_700( .ZN(N3069), .A(N2605) );
  INV_X1 NOT1_701( .ZN(N3070), .A(N2614) );
  INV_X1 NOT1_702( .ZN(N3071), .A(N2623) );
  INV_X1 NOT1_703( .ZN(N3072), .A(N2560) );
  INV_X1 NOT1_704( .ZN(N3073), .A(N2569) );
  INV_X1 NOT1_705( .ZN(N3074), .A(N2578) );
  INV_X1 NOT1_706( .ZN(N3075), .A(N2587) );
  INV_X1 NOT1_707( .ZN(N3076), .A(N2596) );
  INV_X1 NOT1_708( .ZN(N3077), .A(N2605) );
  INV_X1 NOT1_709( .ZN(N3078), .A(N2614) );
  INV_X1 NOT1_710( .ZN(N3079), .A(N2623) );
  INV_X1 NOT1_711( .ZN(N3080), .A(N2560) );
  INV_X1 NOT1_712( .ZN(N3081), .A(N2569) );
  INV_X1 NOT1_713( .ZN(N3082), .A(N2578) );
  INV_X1 NOT1_714( .ZN(N3083), .A(N2587) );
  INV_X1 NOT1_715( .ZN(N3084), .A(N2596) );
  INV_X1 NOT1_716( .ZN(N3085), .A(N2605) );
  INV_X1 NOT1_717( .ZN(N3086), .A(N2614) );
  INV_X1 NOT1_718( .ZN(N3087), .A(N2623) );
  INV_X1 NOT1_719( .ZN(N3088), .A(N2560) );
  INV_X1 NOT1_720( .ZN(N3089), .A(N2569) );
  INV_X1 NOT1_721( .ZN(N3090), .A(N2578) );
  INV_X1 NOT1_722( .ZN(N3091), .A(N2587) );
  INV_X1 NOT1_723( .ZN(N3092), .A(N2596) );
  INV_X1 NOT1_724( .ZN(N3093), .A(N2605) );
  INV_X1 NOT1_725( .ZN(N3094), .A(N2614) );
  INV_X1 NOT1_726( .ZN(N3095), .A(N2623) );
  INV_X1 NOT1_727( .ZN(N3096), .A(N2560) );
  INV_X1 NOT1_728( .ZN(N3097), .A(N2569) );
  INV_X1 NOT1_729( .ZN(N3098), .A(N2578) );
  INV_X1 NOT1_730( .ZN(N3099), .A(N2587) );
  INV_X1 NOT1_731( .ZN(N3100), .A(N2596) );
  INV_X1 NOT1_732( .ZN(N3101), .A(N2605) );
  INV_X1 NOT1_733( .ZN(N3102), .A(N2614) );
  INV_X1 NOT1_734( .ZN(N3103), .A(N2623) );
  INV_X1 NOT1_735( .ZN(N3104), .A(N2560) );
  INV_X1 NOT1_736( .ZN(N3105), .A(N2569) );
  INV_X1 NOT1_737( .ZN(N3106), .A(N2578) );
  INV_X1 NOT1_738( .ZN(N3107), .A(N2587) );
  INV_X1 NOT1_739( .ZN(N3108), .A(N2596) );
  INV_X1 NOT1_740( .ZN(N3109), .A(N2605) );
  INV_X1 NOT1_741( .ZN(N3110), .A(N2614) );
  INV_X1 NOT1_742( .ZN(N3111), .A(N2623) );
  BUF_X1 BUFF1_743( .Z(N3112), .A(N2656) );
  INV_X1 NOT1_744( .ZN(N3115), .A(N2656) );
  INV_X1 NOT1_745( .ZN(N3118), .A(N2652) );
  AND2_X1 AND2_746( .ZN(N3119), .A1(N2768), .A2(N1674) );
  BUF_X1 BUFF1_747( .Z(N3122), .A(N2659) );
  INV_X1 NOT1_748( .ZN(N3125), .A(N2659) );
  BUF_X1 BUFF1_749( .Z(N3128), .A(N2670) );
  INV_X1 NOT1_750( .ZN(N3131), .A(N2670) );
  INV_X1 NOT1_751( .ZN(N3134), .A(N2666) );
  BUF_X1 BUFF1_752( .Z(N3135), .A(N2681) );
  INV_X1 NOT1_753( .ZN(N3138), .A(N2681) );
  INV_X1 NOT1_754( .ZN(N3141), .A(N2677) );
  BUF_X1 BUFF1_755( .Z(N3142), .A(N2692) );
  INV_X1 NOT1_756( .ZN(N3145), .A(N2692) );
  INV_X1 NOT1_757( .ZN(N3148), .A(N2688) );
  AND2_X1 AND2_758( .ZN(N3149), .A1(N2769), .A2(N1678) );
  BUF_X1 BUFF1_759( .Z(N3152), .A(N2697) );
  INV_X1 NOT1_760( .ZN(N3155), .A(N2697) );
  BUF_X1 BUFF1_761( .Z(N3158), .A(N2710) );
  INV_X1 NOT1_762( .ZN(N3161), .A(N2710) );
  INV_X1 NOT1_763( .ZN(N3164), .A(N2706) );
  BUF_X1 BUFF1_764( .Z(N3165), .A(N2723) );
  INV_X1 NOT1_765( .ZN(N3168), .A(N2723) );
  INV_X1 NOT1_766( .ZN(N3171), .A(N2719) );
  AND2_X1 AND2_767( .ZN(N3172), .A1(N1909), .A2(N2648) );
  AND2_X1 AND2_768( .ZN(N3175), .A1(N1913), .A2(N2662) );
  AND2_X1 AND2_769( .ZN(N3178), .A1(N1913), .A2(N2673) );
  AND2_X1 AND2_770( .ZN(N3181), .A1(N1913), .A2(N2684) );
  AND2_X1 AND2_771( .ZN(N3184), .A1(N1922), .A2(N2702) );
  AND2_X1 AND2_772( .ZN(N3187), .A1(N1922), .A2(N2715) );
  INV_X1 NOT1_773( .ZN(N3190), .A(N2692) );
  INV_X1 NOT1_774( .ZN(N3191), .A(N2697) );
  INV_X1 NOT1_775( .ZN(N3192), .A(N2710) );
  INV_X1 NOT1_776( .ZN(N3193), .A(N2723) );
  AND4_X1 AND5_777_A( .ZN(extra0), .A1(N2692), .A2(N2697), .A3(N2710), .A4(N2723) );
  AND2_X1 AND5_777( .ZN(N3194), .A1(extra0), .A2(N1459) );
  NAND2_X1 NAND2_778( .ZN(N3195), .A1(N2745), .A2(N2962) );
  INV_X1 NOT1_779( .ZN(N3196), .A(N2966) );
  OR3_X1 OR3_780( .ZN(N3206), .A1(N2980), .A2(N2145), .A3(N2347) );
  AND2_X1 AND2_781( .ZN(N3207), .A1(N124), .A2(N2984) );
  AND2_X1 AND2_782( .ZN(N3208), .A1(N159), .A2(N2985) );
  AND2_X1 AND2_783( .ZN(N3209), .A1(N150), .A2(N2986) );
  AND2_X1 AND2_784( .ZN(N3210), .A1(N143), .A2(N2987) );
  AND2_X1 AND2_785( .ZN(N3211), .A1(N137), .A2(N2988) );
  AND2_X1 AND2_786( .ZN(N3212), .A1(N132), .A2(N2989) );
  AND2_X1 AND2_787( .ZN(N3213), .A1(N128), .A2(N2990) );
  AND2_X1 AND2_788( .ZN(N3214), .A1(N125), .A2(N2991) );
  AND2_X1 AND2_789( .ZN(N3215), .A1(N125), .A2(N2992) );
  AND2_X1 AND2_790( .ZN(N3216), .A1(N655), .A2(N2993) );
  AND2_X1 AND2_791( .ZN(N3217), .A1(N159), .A2(N2994) );
  AND2_X1 AND2_792( .ZN(N3218), .A1(N150), .A2(N2995) );
  AND2_X1 AND2_793( .ZN(N3219), .A1(N143), .A2(N2996) );
  AND2_X1 AND2_794( .ZN(N3220), .A1(N137), .A2(N2997) );
  AND2_X1 AND2_795( .ZN(N3221), .A1(N132), .A2(N2998) );
  AND2_X1 AND2_796( .ZN(N3222), .A1(N128), .A2(N2999) );
  AND2_X1 AND2_797( .ZN(N3223), .A1(N128), .A2(N3000) );
  AND2_X1 AND2_798( .ZN(N3224), .A1(N670), .A2(N3001) );
  AND2_X1 AND2_799( .ZN(N3225), .A1(N655), .A2(N3002) );
  AND2_X1 AND2_800( .ZN(N3226), .A1(N159), .A2(N3003) );
  AND2_X1 AND2_801( .ZN(N3227), .A1(N150), .A2(N3004) );
  AND2_X1 AND2_802( .ZN(N3228), .A1(N143), .A2(N3005) );
  AND2_X1 AND2_803( .ZN(N3229), .A1(N137), .A2(N3006) );
  AND2_X1 AND2_804( .ZN(N3230), .A1(N132), .A2(N3007) );
  AND2_X1 AND2_805( .ZN(N3231), .A1(N132), .A2(N3008) );
  AND2_X1 AND2_806( .ZN(N3232), .A1(N690), .A2(N3009) );
  AND2_X1 AND2_807( .ZN(N3233), .A1(N670), .A2(N3010) );
  AND2_X1 AND2_808( .ZN(N3234), .A1(N655), .A2(N3011) );
  AND2_X1 AND2_809( .ZN(N3235), .A1(N159), .A2(N3012) );
  AND2_X1 AND2_810( .ZN(N3236), .A1(N150), .A2(N3013) );
  AND2_X1 AND2_811( .ZN(N3237), .A1(N143), .A2(N3014) );
  AND2_X1 AND2_812( .ZN(N3238), .A1(N137), .A2(N3015) );
  AND2_X1 AND2_813( .ZN(N3239), .A1(N137), .A2(N3016) );
  AND2_X1 AND2_814( .ZN(N3240), .A1(N706), .A2(N3017) );
  AND2_X1 AND2_815( .ZN(N3241), .A1(N690), .A2(N3018) );
  AND2_X1 AND2_816( .ZN(N3242), .A1(N670), .A2(N3019) );
  AND2_X1 AND2_817( .ZN(N3243), .A1(N655), .A2(N3020) );
  AND2_X1 AND2_818( .ZN(N3244), .A1(N159), .A2(N3021) );
  AND2_X1 AND2_819( .ZN(N3245), .A1(N150), .A2(N3022) );
  AND2_X1 AND2_820( .ZN(N3246), .A1(N143), .A2(N3023) );
  AND2_X1 AND2_821( .ZN(N3247), .A1(N143), .A2(N3024) );
  AND2_X1 AND2_822( .ZN(N3248), .A1(N715), .A2(N3025) );
  AND2_X1 AND2_823( .ZN(N3249), .A1(N706), .A2(N3026) );
  AND2_X1 AND2_824( .ZN(N3250), .A1(N690), .A2(N3027) );
  AND2_X1 AND2_825( .ZN(N3251), .A1(N670), .A2(N3028) );
  AND2_X1 AND2_826( .ZN(N3252), .A1(N655), .A2(N3029) );
  AND2_X1 AND2_827( .ZN(N3253), .A1(N159), .A2(N3030) );
  AND2_X1 AND2_828( .ZN(N3254), .A1(N150), .A2(N3031) );
  AND2_X1 AND2_829( .ZN(N3255), .A1(N150), .A2(N3032) );
  AND2_X1 AND2_830( .ZN(N3256), .A1(N727), .A2(N3033) );
  AND2_X1 AND2_831( .ZN(N3257), .A1(N715), .A2(N3034) );
  AND2_X1 AND2_832( .ZN(N3258), .A1(N706), .A2(N3035) );
  AND2_X1 AND2_833( .ZN(N3259), .A1(N690), .A2(N3036) );
  AND2_X1 AND2_834( .ZN(N3260), .A1(N670), .A2(N3037) );
  AND2_X1 AND2_835( .ZN(N3261), .A1(N655), .A2(N3038) );
  AND2_X1 AND2_836( .ZN(N3262), .A1(N159), .A2(N3039) );
  AND2_X1 AND2_837( .ZN(N3263), .A1(N159), .A2(N3040) );
  AND2_X1 AND2_838( .ZN(N3264), .A1(N740), .A2(N3041) );
  AND2_X1 AND2_839( .ZN(N3265), .A1(N727), .A2(N3042) );
  AND2_X1 AND2_840( .ZN(N3266), .A1(N715), .A2(N3043) );
  AND2_X1 AND2_841( .ZN(N3267), .A1(N706), .A2(N3044) );
  AND2_X1 AND2_842( .ZN(N3268), .A1(N690), .A2(N3045) );
  AND2_X1 AND2_843( .ZN(N3269), .A1(N670), .A2(N3046) );
  AND2_X1 AND2_844( .ZN(N3270), .A1(N655), .A2(N3047) );
  AND2_X1 AND2_845( .ZN(N3271), .A1(N283), .A2(N3048) );
  AND2_X1 AND2_846( .ZN(N3272), .A1(N670), .A2(N3049) );
  AND2_X1 AND2_847( .ZN(N3273), .A1(N690), .A2(N3050) );
  AND2_X1 AND2_848( .ZN(N3274), .A1(N706), .A2(N3051) );
  AND2_X1 AND2_849( .ZN(N3275), .A1(N715), .A2(N3052) );
  AND2_X1 AND2_850( .ZN(N3276), .A1(N727), .A2(N3053) );
  AND2_X1 AND2_851( .ZN(N3277), .A1(N740), .A2(N3054) );
  AND2_X1 AND2_852( .ZN(N3278), .A1(N753), .A2(N3055) );
  AND2_X1 AND2_853( .ZN(N3279), .A1(N294), .A2(N3056) );
  AND2_X1 AND2_854( .ZN(N3280), .A1(N690), .A2(N3057) );
  AND2_X1 AND2_855( .ZN(N3281), .A1(N706), .A2(N3058) );
  AND2_X1 AND2_856( .ZN(N3282), .A1(N715), .A2(N3059) );
  AND2_X1 AND2_857( .ZN(N3283), .A1(N727), .A2(N3060) );
  AND2_X1 AND2_858( .ZN(N3284), .A1(N740), .A2(N3061) );
  AND2_X1 AND2_859( .ZN(N3285), .A1(N753), .A2(N3062) );
  AND2_X1 AND2_860( .ZN(N3286), .A1(N283), .A2(N3063) );
  AND2_X1 AND2_861( .ZN(N3287), .A1(N303), .A2(N3064) );
  AND2_X1 AND2_862( .ZN(N3288), .A1(N706), .A2(N3065) );
  AND2_X1 AND2_863( .ZN(N3289), .A1(N715), .A2(N3066) );
  AND2_X1 AND2_864( .ZN(N3290), .A1(N727), .A2(N3067) );
  AND2_X1 AND2_865( .ZN(N3291), .A1(N740), .A2(N3068) );
  AND2_X1 AND2_866( .ZN(N3292), .A1(N753), .A2(N3069) );
  AND2_X1 AND2_867( .ZN(N3293), .A1(N283), .A2(N3070) );
  AND2_X1 AND2_868( .ZN(N3294), .A1(N294), .A2(N3071) );
  AND2_X1 AND2_869( .ZN(N3295), .A1(N311), .A2(N3072) );
  AND2_X1 AND2_870( .ZN(N3296), .A1(N715), .A2(N3073) );
  AND2_X1 AND2_871( .ZN(N3297), .A1(N727), .A2(N3074) );
  AND2_X1 AND2_872( .ZN(N3298), .A1(N740), .A2(N3075) );
  AND2_X1 AND2_873( .ZN(N3299), .A1(N753), .A2(N3076) );
  AND2_X1 AND2_874( .ZN(N3300), .A1(N283), .A2(N3077) );
  AND2_X1 AND2_875( .ZN(N3301), .A1(N294), .A2(N3078) );
  AND2_X1 AND2_876( .ZN(N3302), .A1(N303), .A2(N3079) );
  AND2_X1 AND2_877( .ZN(N3303), .A1(N317), .A2(N3080) );
  AND2_X1 AND2_878( .ZN(N3304), .A1(N727), .A2(N3081) );
  AND2_X1 AND2_879( .ZN(N3305), .A1(N740), .A2(N3082) );
  AND2_X1 AND2_880( .ZN(N3306), .A1(N753), .A2(N3083) );
  AND2_X1 AND2_881( .ZN(N3307), .A1(N283), .A2(N3084) );
  AND2_X1 AND2_882( .ZN(N3308), .A1(N294), .A2(N3085) );
  AND2_X1 AND2_883( .ZN(N3309), .A1(N303), .A2(N3086) );
  AND2_X1 AND2_884( .ZN(N3310), .A1(N311), .A2(N3087) );
  AND2_X1 AND2_885( .ZN(N3311), .A1(N322), .A2(N3088) );
  AND2_X1 AND2_886( .ZN(N3312), .A1(N740), .A2(N3089) );
  AND2_X1 AND2_887( .ZN(N3313), .A1(N753), .A2(N3090) );
  AND2_X1 AND2_888( .ZN(N3314), .A1(N283), .A2(N3091) );
  AND2_X1 AND2_889( .ZN(N3315), .A1(N294), .A2(N3092) );
  AND2_X1 AND2_890( .ZN(N3316), .A1(N303), .A2(N3093) );
  AND2_X1 AND2_891( .ZN(N3317), .A1(N311), .A2(N3094) );
  AND2_X1 AND2_892( .ZN(N3318), .A1(N317), .A2(N3095) );
  AND2_X1 AND2_893( .ZN(N3319), .A1(N326), .A2(N3096) );
  AND2_X1 AND2_894( .ZN(N3320), .A1(N753), .A2(N3097) );
  AND2_X1 AND2_895( .ZN(N3321), .A1(N283), .A2(N3098) );
  AND2_X1 AND2_896( .ZN(N3322), .A1(N294), .A2(N3099) );
  AND2_X1 AND2_897( .ZN(N3323), .A1(N303), .A2(N3100) );
  AND2_X1 AND2_898( .ZN(N3324), .A1(N311), .A2(N3101) );
  AND2_X1 AND2_899( .ZN(N3325), .A1(N317), .A2(N3102) );
  AND2_X1 AND2_900( .ZN(N3326), .A1(N322), .A2(N3103) );
  AND2_X1 AND2_901( .ZN(N3327), .A1(N329), .A2(N3104) );
  AND2_X1 AND2_902( .ZN(N3328), .A1(N283), .A2(N3105) );
  AND2_X1 AND2_903( .ZN(N3329), .A1(N294), .A2(N3106) );
  AND2_X1 AND2_904( .ZN(N3330), .A1(N303), .A2(N3107) );
  AND2_X1 AND2_905( .ZN(N3331), .A1(N311), .A2(N3108) );
  AND2_X1 AND2_906( .ZN(N3332), .A1(N317), .A2(N3109) );
  AND2_X1 AND2_907( .ZN(N3333), .A1(N322), .A2(N3110) );
  AND2_X1 AND2_908( .ZN(N3334), .A1(N326), .A2(N3111) );
  AND4_X1 AND5_909_A( .ZN(extra1), .A1(N3190), .A2(N3191), .A3(N3192), .A4(N3193) );
  AND2_X1 AND5_909( .ZN(N3383), .A1(extra1), .A2(N917) );
  BUF_X1 BUFF1_910( .Z(N3384), .A(N2977) );
  AND2_X1 AND2_911( .ZN(N3387), .A1(N3196), .A2(N1736) );
  AND2_X1 AND2_912( .ZN(N3388), .A1(N2977), .A2(N2149) );
  AND2_X1 AND2_913( .ZN(N3389), .A1(N2973), .A2(N1737) );
  NOR3_X1 NOR8_914_A( .ZN(extra2), .A1(N3207), .A2(N3208), .A3(N3209) );
  NOR3_X1 NOR8_914_B( .ZN(extra3), .A1(extra2), .A2(N3210), .A3(N3211) );
  NOR3_X1 NOR8_914_C( .ZN(extra4), .A1(extra3), .A2(N3212), .A3(N3213) );
  NOR2_X1 NOR8_914( .ZN(N3390), .A1(extra4), .A2(N3214) );
  NOR3_X1 NOR8_915_A( .ZN(extra5), .A1(N3215), .A2(N3216), .A3(N3217) );
  NOR3_X1 NOR8_915_B( .ZN(extra6), .A1(extra5), .A2(N3218), .A3(N3219) );
  NOR3_X1 NOR8_915_C( .ZN(extra7), .A1(extra6), .A2(N3220), .A3(N3221) );
  NOR2_X1 NOR8_915( .ZN(N3391), .A1(extra7), .A2(N3222) );
  NOR3_X1 NOR8_916_A( .ZN(extra8), .A1(N3223), .A2(N3224), .A3(N3225) );
  NOR3_X1 NOR8_916_B( .ZN(extra9), .A1(extra8), .A2(N3226), .A3(N3227) );
  NOR3_X1 NOR8_916_C( .ZN(extra10), .A1(extra9), .A2(N3228), .A3(N3229) );
  NOR2_X1 NOR8_916( .ZN(N3392), .A1(extra10), .A2(N3230) );
  NOR3_X1 NOR8_917_A( .ZN(extra11), .A1(N3231), .A2(N3232), .A3(N3233) );
  NOR3_X1 NOR8_917_B( .ZN(extra12), .A1(extra11), .A2(N3234), .A3(N3235) );
  NOR3_X1 NOR8_917_C( .ZN(extra13), .A1(extra12), .A2(N3236), .A3(N3237) );
  NOR2_X1 NOR8_917( .ZN(N3393), .A1(extra13), .A2(N3238) );
  NOR3_X1 NOR8_918_A( .ZN(extra14), .A1(N3239), .A2(N3240), .A3(N3241) );
  NOR3_X1 NOR8_918_B( .ZN(extra15), .A1(extra14), .A2(N3242), .A3(N3243) );
  NOR3_X1 NOR8_918_C( .ZN(extra16), .A1(extra15), .A2(N3244), .A3(N3245) );
  NOR2_X1 NOR8_918( .ZN(N3394), .A1(extra16), .A2(N3246) );
  NOR3_X1 NOR8_919_A( .ZN(extra17), .A1(N3247), .A2(N3248), .A3(N3249) );
  NOR3_X1 NOR8_919_B( .ZN(extra18), .A1(extra17), .A2(N3250), .A3(N3251) );
  NOR3_X1 NOR8_919_C( .ZN(extra19), .A1(extra18), .A2(N3252), .A3(N3253) );
  NOR2_X1 NOR8_919( .ZN(N3395), .A1(extra19), .A2(N3254) );
  NOR3_X1 NOR8_920_A( .ZN(extra20), .A1(N3255), .A2(N3256), .A3(N3257) );
  NOR3_X1 NOR8_920_B( .ZN(extra21), .A1(extra20), .A2(N3258), .A3(N3259) );
  NOR3_X1 NOR8_920_C( .ZN(extra22), .A1(extra21), .A2(N3260), .A3(N3261) );
  NOR2_X1 NOR8_920( .ZN(N3396), .A1(extra22), .A2(N3262) );
  NOR3_X1 NOR8_921_A( .ZN(extra23), .A1(N3263), .A2(N3264), .A3(N3265) );
  NOR3_X1 NOR8_921_B( .ZN(extra24), .A1(extra23), .A2(N3266), .A3(N3267) );
  NOR3_X1 NOR8_921_C( .ZN(extra25), .A1(extra24), .A2(N3268), .A3(N3269) );
  NOR2_X1 NOR8_921( .ZN(N3397), .A1(extra25), .A2(N3270) );
  NOR3_X1 NOR8_922_A( .ZN(extra26), .A1(N3271), .A2(N3272), .A3(N3273) );
  NOR3_X1 NOR8_922_B( .ZN(extra27), .A1(extra26), .A2(N3274), .A3(N3275) );
  NOR3_X1 NOR8_922_C( .ZN(extra28), .A1(extra27), .A2(N3276), .A3(N3277) );
  NOR2_X1 NOR8_922( .ZN(N3398), .A1(extra28), .A2(N3278) );
  NOR3_X1 NOR8_923_A( .ZN(extra29), .A1(N3279), .A2(N3280), .A3(N3281) );
  NOR3_X1 NOR8_923_B( .ZN(extra30), .A1(extra29), .A2(N3282), .A3(N3283) );
  NOR3_X1 NOR8_923_C( .ZN(extra31), .A1(extra30), .A2(N3284), .A3(N3285) );
  NOR2_X1 NOR8_923( .ZN(N3399), .A1(extra31), .A2(N3286) );
  NOR3_X1 NOR8_924_A( .ZN(extra32), .A1(N3287), .A2(N3288), .A3(N3289) );
  NOR3_X1 NOR8_924_B( .ZN(extra33), .A1(extra32), .A2(N3290), .A3(N3291) );
  NOR3_X1 NOR8_924_C( .ZN(extra34), .A1(extra33), .A2(N3292), .A3(N3293) );
  NOR2_X1 NOR8_924( .ZN(N3400), .A1(extra34), .A2(N3294) );
  NOR3_X1 NOR8_925_A( .ZN(extra35), .A1(N3295), .A2(N3296), .A3(N3297) );
  NOR3_X1 NOR8_925_B( .ZN(extra36), .A1(extra35), .A2(N3298), .A3(N3299) );
  NOR3_X1 NOR8_925_C( .ZN(extra37), .A1(extra36), .A2(N3300), .A3(N3301) );
  NOR2_X1 NOR8_925( .ZN(N3401), .A1(extra37), .A2(N3302) );
  NOR3_X1 NOR8_926_A( .ZN(extra38), .A1(N3303), .A2(N3304), .A3(N3305) );
  NOR3_X1 NOR8_926_B( .ZN(extra39), .A1(extra38), .A2(N3306), .A3(N3307) );
  NOR3_X1 NOR8_926_C( .ZN(extra40), .A1(extra39), .A2(N3308), .A3(N3309) );
  NOR2_X1 NOR8_926( .ZN(N3402), .A1(extra40), .A2(N3310) );
  NOR3_X1 NOR8_927_A( .ZN(extra41), .A1(N3311), .A2(N3312), .A3(N3313) );
  NOR3_X1 NOR8_927_B( .ZN(extra42), .A1(extra41), .A2(N3314), .A3(N3315) );
  NOR3_X1 NOR8_927_C( .ZN(extra43), .A1(extra42), .A2(N3316), .A3(N3317) );
  NOR2_X1 NOR8_927( .ZN(N3403), .A1(extra43), .A2(N3318) );
  NOR3_X1 NOR8_928_A( .ZN(extra44), .A1(N3319), .A2(N3320), .A3(N3321) );
  NOR3_X1 NOR8_928_B( .ZN(extra45), .A1(extra44), .A2(N3322), .A3(N3323) );
  NOR3_X1 NOR8_928_C( .ZN(extra46), .A1(extra45), .A2(N3324), .A3(N3325) );
  NOR2_X1 NOR8_928( .ZN(N3404), .A1(extra46), .A2(N3326) );
  NOR3_X1 NOR8_929_A( .ZN(extra47), .A1(N3327), .A2(N3328), .A3(N3329) );
  NOR3_X1 NOR8_929_B( .ZN(extra48), .A1(extra47), .A2(N3330), .A3(N3331) );
  NOR3_X1 NOR8_929_C( .ZN(extra49), .A1(extra48), .A2(N3332), .A3(N3333) );
  NOR2_X1 NOR8_929( .ZN(N3405), .A1(extra49), .A2(N3334) );
  AND2_X1 AND2_930( .ZN(N3406), .A1(N3206), .A2(N2641) );
  AND3_X1 AND3_931( .ZN(N3407), .A1(N169), .A2(N2648), .A3(N3112) );
  AND3_X1 AND3_932( .ZN(N3410), .A1(N179), .A2(N2648), .A3(N3115) );
  AND3_X1 AND3_933( .ZN(N3413), .A1(N190), .A2(N2652), .A3(N3115) );
  AND3_X1 AND3_934( .ZN(N3414), .A1(N200), .A2(N2652), .A3(N3112) );
  OR3_X1 OR3_935( .ZN(N3415), .A1(N3119), .A2(N1875), .A3(N2073) );
  NOR3_X1 NOR3_936( .ZN(N3419), .A1(N3119), .A2(N1875), .A3(N2073) );
  AND3_X1 AND3_937( .ZN(N3423), .A1(N169), .A2(N2662), .A3(N3128) );
  AND3_X1 AND3_938( .ZN(N3426), .A1(N179), .A2(N2662), .A3(N3131) );
  AND3_X1 AND3_939( .ZN(N3429), .A1(N190), .A2(N2666), .A3(N3131) );
  AND3_X1 AND3_940( .ZN(N3430), .A1(N200), .A2(N2666), .A3(N3128) );
  AND3_X1 AND3_941( .ZN(N3431), .A1(N169), .A2(N2673), .A3(N3135) );
  AND3_X1 AND3_942( .ZN(N3434), .A1(N179), .A2(N2673), .A3(N3138) );
  AND3_X1 AND3_943( .ZN(N3437), .A1(N190), .A2(N2677), .A3(N3138) );
  AND3_X1 AND3_944( .ZN(N3438), .A1(N200), .A2(N2677), .A3(N3135) );
  AND3_X1 AND3_945( .ZN(N3439), .A1(N169), .A2(N2684), .A3(N3142) );
  AND3_X1 AND3_946( .ZN(N3442), .A1(N179), .A2(N2684), .A3(N3145) );
  AND3_X1 AND3_947( .ZN(N3445), .A1(N190), .A2(N2688), .A3(N3145) );
  AND3_X1 AND3_948( .ZN(N3446), .A1(N200), .A2(N2688), .A3(N3142) );
  OR3_X1 OR3_949( .ZN(N3447), .A1(N3149), .A2(N1895), .A3(N2093) );
  NOR3_X1 NOR3_950( .ZN(N3451), .A1(N3149), .A2(N1895), .A3(N2093) );
  AND3_X1 AND3_951( .ZN(N3455), .A1(N169), .A2(N2702), .A3(N3158) );
  AND3_X1 AND3_952( .ZN(N3458), .A1(N179), .A2(N2702), .A3(N3161) );
  AND3_X1 AND3_953( .ZN(N3461), .A1(N190), .A2(N2706), .A3(N3161) );
  AND3_X1 AND3_954( .ZN(N3462), .A1(N200), .A2(N2706), .A3(N3158) );
  AND3_X1 AND3_955( .ZN(N3463), .A1(N169), .A2(N2715), .A3(N3165) );
  AND3_X1 AND3_956( .ZN(N3466), .A1(N179), .A2(N2715), .A3(N3168) );
  AND3_X1 AND3_957( .ZN(N3469), .A1(N190), .A2(N2719), .A3(N3168) );
  AND3_X1 AND3_958( .ZN(N3470), .A1(N200), .A2(N2719), .A3(N3165) );
  OR2_X1 OR2_959( .ZN(N3471), .A1(N3194), .A2(N3383) );
  BUF_X1 BUFF1_960( .Z(N3472), .A(N2967) );
  BUF_X1 BUFF1_961( .Z(N3475), .A(N2970) );
  BUF_X1 BUFF1_962( .Z(N3478), .A(N2967) );
  BUF_X1 BUFF1_963( .Z(N3481), .A(N2970) );
  BUF_X1 BUFF1_964( .Z(N3484), .A(N2973) );
  BUF_X1 BUFF1_965( .Z(N3487), .A(N2973) );
  BUF_X1 BUFF1_966( .Z(N3490), .A(N3172) );
  BUF_X1 BUFF1_967( .Z(N3493), .A(N3172) );
  BUF_X1 BUFF1_968( .Z(N3496), .A(N3175) );
  BUF_X1 BUFF1_969( .Z(N3499), .A(N3175) );
  BUF_X1 BUFF1_970( .Z(N3502), .A(N3178) );
  BUF_X1 BUFF1_971( .Z(N3505), .A(N3178) );
  BUF_X1 BUFF1_972( .Z(N3508), .A(N3181) );
  BUF_X1 BUFF1_973( .Z(N3511), .A(N3181) );
  BUF_X1 BUFF1_974( .Z(N3514), .A(N3184) );
  BUF_X1 BUFF1_975( .Z(N3517), .A(N3184) );
  BUF_X1 BUFF1_976( .Z(N3520), .A(N3187) );
  BUF_X1 BUFF1_977( .Z(N3523), .A(N3187) );
  NOR2_X1 NOR2_978( .ZN(N3534), .A1(N3387), .A2(N2350) );
  OR3_X1 OR3_979( .ZN(N3535), .A1(N3388), .A2(N2151), .A3(N2351) );
  NOR2_X1 NOR2_980( .ZN(N3536), .A1(N3389), .A2(N1966) );
  AND2_X1 AND2_981( .ZN(N3537), .A1(N3390), .A2(N2209) );
  AND2_X1 AND2_982( .ZN(N3538), .A1(N3398), .A2(N2210) );
  AND2_X1 AND2_983( .ZN(N3539), .A1(N3391), .A2(N1842) );
  AND2_X1 AND2_984( .ZN(N3540), .A1(N3399), .A2(N1369) );
  AND2_X1 AND2_985( .ZN(N3541), .A1(N3392), .A2(N1843) );
  AND2_X1 AND2_986( .ZN(N3542), .A1(N3400), .A2(N1369) );
  AND2_X1 AND2_987( .ZN(N3543), .A1(N3393), .A2(N1844) );
  AND2_X1 AND2_988( .ZN(N3544), .A1(N3401), .A2(N1369) );
  AND2_X1 AND2_989( .ZN(N3545), .A1(N3394), .A2(N1845) );
  AND2_X1 AND2_990( .ZN(N3546), .A1(N3402), .A2(N1369) );
  AND2_X1 AND2_991( .ZN(N3547), .A1(N3395), .A2(N1846) );
  AND2_X1 AND2_992( .ZN(N3548), .A1(N3403), .A2(N1369) );
  AND2_X1 AND2_993( .ZN(N3549), .A1(N3396), .A2(N1847) );
  AND2_X1 AND2_994( .ZN(N3550), .A1(N3404), .A2(N1369) );
  AND2_X1 AND2_995( .ZN(N3551), .A1(N3397), .A2(N1848) );
  AND2_X1 AND2_996( .ZN(N3552), .A1(N3405), .A2(N1369) );
  OR3_X1 OR3_997( .ZN(N3557), .A1(N3413), .A2(N3414), .A3(N3118) );
  OR3_X1 OR3_998( .ZN(N3568), .A1(N3429), .A2(N3430), .A3(N3134) );
  OR3_X1 OR3_999( .ZN(N3573), .A1(N3437), .A2(N3438), .A3(N3141) );
  OR3_X1 OR3_1000( .ZN(N3578), .A1(N3445), .A2(N3446), .A3(N3148) );
  OR3_X1 OR3_1001( .ZN(N3589), .A1(N3461), .A2(N3462), .A3(N3164) );
  OR3_X1 OR3_1002( .ZN(N3594), .A1(N3469), .A2(N3470), .A3(N3171) );
  AND2_X1 AND2_1003( .ZN(N3605), .A1(N3471), .A2(N2728) );
  INV_X32 NOT1_1004( .ZN(N3626), .A(N3478) );
  INV_X32 NOT1_1005( .ZN(N3627), .A(N3481) );
  INV_X32 NOT1_1006( .ZN(N3628), .A(N3487) );
  INV_X1 NOT1_1007( .ZN(N3629), .A(N3484) );
  INV_X1 NOT1_1008( .ZN(N3630), .A(N3472) );
  INV_X1 NOT1_1009( .ZN(N3631), .A(N3475) );
  AND2_X1 AND2_1010( .ZN(N3632), .A1(N3536), .A2(N2152) );
  AND2_X1 AND2_1011( .ZN(N3633), .A1(N3534), .A2(N2155) );
  OR3_X1 OR3_1012( .ZN(N3634), .A1(N3537), .A2(N3538), .A3(N2398) );
  OR2_X1 OR2_1013( .ZN(N3635), .A1(N3539), .A2(N3540) );
  OR2_X1 OR2_1014( .ZN(N3636), .A1(N3541), .A2(N3542) );
  OR2_X1 OR2_1015( .ZN(N3637), .A1(N3543), .A2(N3544) );
  OR2_X1 OR2_1016( .ZN(N3638), .A1(N3545), .A2(N3546) );
  OR2_X1 OR2_1017( .ZN(N3639), .A1(N3547), .A2(N3548) );
  OR2_X1 OR2_1018( .ZN(N3640), .A1(N3549), .A2(N3550) );
  OR2_X1 OR2_1019( .ZN(N3641), .A1(N3551), .A2(N3552) );
  AND2_X1 AND2_1020( .ZN(N3642), .A1(N3535), .A2(N2643) );
  OR2_X1 OR2_1021( .ZN(N3643), .A1(N3407), .A2(N3410) );
  NOR2_X1 NOR2_1022( .ZN(N3644), .A1(N3407), .A2(N3410) );
  AND3_X1 AND3_1023( .ZN(N3645), .A1(N169), .A2(N3415), .A3(N3122) );
  AND3_X1 AND3_1024( .ZN(N3648), .A1(N179), .A2(N3415), .A3(N3125) );
  AND3_X1 AND3_1025( .ZN(N3651), .A1(N190), .A2(N3419), .A3(N3125) );
  AND3_X1 AND3_1026( .ZN(N3652), .A1(N200), .A2(N3419), .A3(N3122) );
  INV_X1 NOT1_1027( .ZN(N3653), .A(N3419) );
  OR2_X1 OR2_1028( .ZN(N3654), .A1(N3423), .A2(N3426) );
  NOR2_X1 NOR2_1029( .ZN(N3657), .A1(N3423), .A2(N3426) );
  OR2_X1 OR2_1030( .ZN(N3658), .A1(N3431), .A2(N3434) );
  NOR2_X1 NOR2_1031( .ZN(N3661), .A1(N3431), .A2(N3434) );
  OR2_X1 OR2_1032( .ZN(N3662), .A1(N3439), .A2(N3442) );
  NOR2_X1 NOR2_1033( .ZN(N3663), .A1(N3439), .A2(N3442) );
  AND3_X1 AND3_1034( .ZN(N3664), .A1(N169), .A2(N3447), .A3(N3152) );
  AND3_X1 AND3_1035( .ZN(N3667), .A1(N179), .A2(N3447), .A3(N3155) );
  AND3_X1 AND3_1036( .ZN(N3670), .A1(N190), .A2(N3451), .A3(N3155) );
  AND3_X1 AND3_1037( .ZN(N3671), .A1(N200), .A2(N3451), .A3(N3152) );
  INV_X1 NOT1_1038( .ZN(N3672), .A(N3451) );
  OR2_X1 OR2_1039( .ZN(N3673), .A1(N3455), .A2(N3458) );
  NOR2_X1 NOR2_1040( .ZN(N3676), .A1(N3455), .A2(N3458) );
  OR2_X1 OR2_1041( .ZN(N3677), .A1(N3463), .A2(N3466) );
  NOR2_X1 NOR2_1042( .ZN(N3680), .A1(N3463), .A2(N3466) );
  INV_X1 NOT1_1043( .ZN(N3681), .A(N3493) );
  AND2_X1 AND2_1044( .ZN(N3682), .A1(N1909), .A2(N3415) );
  INV_X1 NOT1_1045( .ZN(N3685), .A(N3496) );
  INV_X1 NOT1_1046( .ZN(N3686), .A(N3499) );
  INV_X1 NOT1_1047( .ZN(N3687), .A(N3502) );
  INV_X1 NOT1_1048( .ZN(N3688), .A(N3505) );
  INV_X1 NOT1_1049( .ZN(N3689), .A(N3511) );
  AND2_X1 AND2_1050( .ZN(N3690), .A1(N1922), .A2(N3447) );
  INV_X1 NOT1_1051( .ZN(N3693), .A(N3517) );
  INV_X1 NOT1_1052( .ZN(N3694), .A(N3520) );
  INV_X1 NOT1_1053( .ZN(N3695), .A(N3523) );
  INV_X1 NOT1_1054( .ZN(N3696), .A(N3514) );
  BUF_X1 BUFF1_1055( .Z(N3697), .A(N3384) );
  BUF_X1 BUFF1_1056( .Z(N3700), .A(N3384) );
  INV_X1 NOT1_1057( .ZN(N3703), .A(N3490) );
  INV_X1 NOT1_1058( .ZN(N3704), .A(N3508) );
  NAND2_X1 NAND2_1059( .ZN(N3705), .A1(N3475), .A2(N3630) );
  NAND2_X1 NAND2_1060( .ZN(N3706), .A1(N3472), .A2(N3631) );
  NAND2_X1 NAND2_1061( .ZN(N3707), .A1(N3481), .A2(N3626) );
  NAND2_X1 NAND2_1062( .ZN(N3708), .A1(N3478), .A2(N3627) );
  OR3_X1 OR3_1063( .ZN(N3711), .A1(N3632), .A2(N2352), .A3(N2353) );
  OR3_X1 OR3_1064( .ZN(N3712), .A1(N3633), .A2(N2354), .A3(N2355) );
  AND2_X1 AND2_1065( .ZN(N3713), .A1(N3634), .A2(N2632) );
  AND2_X1 AND2_1066( .ZN(N3714), .A1(N3635), .A2(N2634) );
  AND2_X1 AND2_1067( .ZN(N3715), .A1(N3636), .A2(N2636) );
  AND2_X1 AND2_1068( .ZN(N3716), .A1(N3637), .A2(N2638) );
  AND2_X1 AND2_1069( .ZN(N3717), .A1(N3638), .A2(N2640) );
  AND2_X1 AND2_1070( .ZN(N3718), .A1(N3639), .A2(N2642) );
  AND2_X1 AND2_1071( .ZN(N3719), .A1(N3640), .A2(N2644) );
  AND2_X1 AND2_1072( .ZN(N3720), .A1(N3641), .A2(N2646) );
  AND2_X1 AND2_1073( .ZN(N3721), .A1(N3644), .A2(N3557) );
  OR3_X1 OR3_1074( .ZN(N3731), .A1(N3651), .A2(N3652), .A3(N3653) );
  AND2_X1 AND2_1075( .ZN(N3734), .A1(N3657), .A2(N3568) );
  AND2_X1 AND2_1076( .ZN(N3740), .A1(N3661), .A2(N3573) );
  AND2_X1 AND2_1077( .ZN(N3743), .A1(N3663), .A2(N3578) );
  OR3_X1 OR3_1078( .ZN(N3753), .A1(N3670), .A2(N3671), .A3(N3672) );
  AND2_X1 AND2_1079( .ZN(N3756), .A1(N3676), .A2(N3589) );
  AND2_X1 AND2_1080( .ZN(N3762), .A1(N3680), .A2(N3594) );
  INV_X1 NOT1_1081( .ZN(N3765), .A(N3643) );
  INV_X1 NOT1_1082( .ZN(N3766), .A(N3662) );
  NAND2_X1 NAND2_1083( .ZN(N3773), .A1(N3705), .A2(N3706) );
  NAND2_X1 NAND2_1084( .ZN(N3774), .A1(N3707), .A2(N3708) );
  NAND2_X1 NAND2_1085( .ZN(N3775), .A1(N3700), .A2(N3628) );
  INV_X1 NOT1_1086( .ZN(N3776), .A(N3700) );
  NAND2_X1 NAND2_1087( .ZN(N3777), .A1(N3697), .A2(N3629) );
  INV_X1 NOT1_1088( .ZN(N3778), .A(N3697) );
  AND2_X1 AND2_1089( .ZN(N3779), .A1(N3712), .A2(N2645) );
  AND2_X1 AND2_1090( .ZN(N3780), .A1(N3711), .A2(N2647) );
  OR2_X1 OR2_1091( .ZN(N3786), .A1(N3645), .A2(N3648) );
  NOR2_X1 NOR2_1092( .ZN(N3789), .A1(N3645), .A2(N3648) );
  OR2_X1 OR2_1093( .ZN(N3800), .A1(N3664), .A2(N3667) );
  NOR2_X1 NOR2_1094( .ZN(N3803), .A1(N3664), .A2(N3667) );
  AND2_X1 AND2_1095( .ZN(N3809), .A1(N3654), .A2(N1917) );
  AND2_X1 AND2_1096( .ZN(N3812), .A1(N3658), .A2(N1917) );
  AND2_X1 AND2_1097( .ZN(N3815), .A1(N3673), .A2(N1926) );
  AND2_X1 AND2_1098( .ZN(N3818), .A1(N3677), .A2(N1926) );
  BUF_X1 BUFF1_1099( .Z(N3821), .A(N3682) );
  BUF_X1 BUFF1_1100( .Z(N3824), .A(N3682) );
  BUF_X1 BUFF1_1101( .Z(N3827), .A(N3690) );
  BUF_X1 BUFF1_1102( .Z(N3830), .A(N3690) );
  NAND2_X1 NAND2_1103( .ZN(N3833), .A1(N3773), .A2(N3774) );
  NAND2_X1 NAND2_1104( .ZN(N3834), .A1(N3487), .A2(N3776) );
  NAND2_X1 NAND2_1105( .ZN(N3835), .A1(N3484), .A2(N3778) );
  AND2_X1 AND2_1106( .ZN(N3838), .A1(N3789), .A2(N3731) );
  AND2_X1 AND2_1107( .ZN(N3845), .A1(N3803), .A2(N3753) );
  BUF_X1 BUFF1_1108( .Z(N3850), .A(N3721) );
  BUF_X1 BUFF1_1109( .Z(N3855), .A(N3734) );
  BUF_X1 BUFF1_1110( .Z(N3858), .A(N3740) );
  BUF_X1 BUFF1_1111( .Z(N3861), .A(N3743) );
  BUF_X1 BUFF1_1112( .Z(N3865), .A(N3756) );
  BUF_X1 BUFF1_1113( .Z(N3868), .A(N3762) );
  NAND2_X1 NAND2_1114( .ZN(N3884), .A1(N3775), .A2(N3834) );
  NAND2_X1 NAND2_1115( .ZN(N3885), .A1(N3777), .A2(N3835) );
  NAND2_X1 NAND2_1116( .ZN(N3894), .A1(N3721), .A2(N3786) );
  NAND2_X1 NAND2_1117( .ZN(N3895), .A1(N3743), .A2(N3800) );
  INV_X1 NOT1_1118( .ZN(N3898), .A(N3821) );
  INV_X1 NOT1_1119( .ZN(N3899), .A(N3824) );
  INV_X1 NOT1_1120( .ZN(N3906), .A(N3830) );
  INV_X1 NOT1_1121( .ZN(N3911), .A(N3827) );
  AND2_X1 AND2_1122( .ZN(N3912), .A1(N3786), .A2(N1912) );
  BUF_X1 BUFF1_1123( .Z(N3913), .A(N3812) );
  AND2_X1 AND2_1124( .ZN(N3916), .A1(N3800), .A2(N1917) );
  BUF_X1 BUFF1_1125( .Z(N3917), .A(N3818) );
  INV_X1 NOT1_1126( .ZN(N3920), .A(N3809) );
  BUF_X1 BUFF1_1127( .Z(N3921), .A(N3818) );
  INV_X1 NOT1_1128( .ZN(N3924), .A(N3884) );
  INV_X1 NOT1_1129( .ZN(N3925), .A(N3885) );
  AND4_X1 AND4_1130( .ZN(N3926), .A1(N3721), .A2(N3838), .A3(N3734), .A4(N3740) );
  NAND3_X1 NAND3_1131( .ZN(N3930), .A1(N3721), .A2(N3838), .A3(N3654) );
  NAND4_X1 NAND4_1132( .ZN(N3931), .A1(N3658), .A2(N3838), .A3(N3734), .A4(N3721) );
  AND4_X1 AND4_1133( .ZN(N3932), .A1(N3743), .A2(N3845), .A3(N3756), .A4(N3762) );
  NAND3_X1 NAND3_1134( .ZN(N3935), .A1(N3743), .A2(N3845), .A3(N3673) );
  NAND4_X1 NAND4_1135( .ZN(N3936), .A1(N3677), .A2(N3845), .A3(N3756), .A4(N3743) );
  BUF_X1 BUFF1_1136( .Z(N3937), .A(N3838) );
  BUF_X1 BUFF1_1137( .Z(N3940), .A(N3845) );
  INV_X1 NOT1_1138( .ZN(N3947), .A(N3912) );
  INV_X1 NOT1_1139( .ZN(N3948), .A(N3916) );
  BUF_X1 BUFF1_1140( .Z(N3950), .A(N3850) );
  BUF_X1 BUFF1_1141( .Z(N3953), .A(N3850) );
  BUF_X1 BUFF1_1142( .Z(N3956), .A(N3855) );
  BUF_X1 BUFF1_1143( .Z(N3959), .A(N3855) );
  BUF_X1 BUFF1_1144( .Z(N3962), .A(N3858) );
  BUF_X1 BUFF1_1145( .Z(N3965), .A(N3858) );
  BUF_X1 BUFF1_1146( .Z(N3968), .A(N3861) );
  BUF_X1 BUFF1_1147( .Z(N3971), .A(N3861) );
  BUF_X1 BUFF1_1148( .Z(N3974), .A(N3865) );
  BUF_X1 BUFF1_1149( .Z(N3977), .A(N3865) );
  BUF_X1 BUFF1_1150( .Z(N3980), .A(N3868) );
  BUF_X1 BUFF1_1151( .Z(N3983), .A(N3868) );
  NAND2_X1 NAND2_1152( .ZN(N3987), .A1(N3924), .A2(N3925) );
  NAND4_X1 NAND4_1153( .ZN(N3992), .A1(N3765), .A2(N3894), .A3(N3930), .A4(N3931) );
  NAND4_X1 NAND4_1154( .ZN(N3996), .A1(N3766), .A2(N3895), .A3(N3935), .A4(N3936) );
  INV_X1 NOT1_1155( .ZN(N4013), .A(N3921) );
  AND2_X1 AND2_1156( .ZN(N4028), .A1(N3932), .A2(N3926) );
  NAND2_X1 NAND2_1157( .ZN(N4029), .A1(N3953), .A2(N3681) );
  NAND2_X1 NAND2_1158( .ZN(N4030), .A1(N3959), .A2(N3686) );
  NAND2_X1 NAND2_1159( .ZN(N4031), .A1(N3965), .A2(N3688) );
  NAND2_X1 NAND2_1160( .ZN(N4032), .A1(N3971), .A2(N3689) );
  NAND2_X1 NAND2_1161( .ZN(N4033), .A1(N3977), .A2(N3693) );
  NAND2_X1 NAND2_1162( .ZN(N4034), .A1(N3983), .A2(N3695) );
  BUF_X1 BUFF1_1163( .Z(N4035), .A(N3926) );
  INV_X1 NOT1_1164( .ZN(N4042), .A(N3953) );
  INV_X1 NOT1_1165( .ZN(N4043), .A(N3956) );
  NAND2_X1 NAND2_1166( .ZN(N4044), .A1(N3956), .A2(N3685) );
  INV_X1 NOT1_1167( .ZN(N4045), .A(N3959) );
  INV_X1 NOT1_1168( .ZN(N4046), .A(N3962) );
  NAND2_X1 NAND2_1169( .ZN(N4047), .A1(N3962), .A2(N3687) );
  INV_X1 NOT1_1170( .ZN(N4048), .A(N3965) );
  INV_X1 NOT1_1171( .ZN(N4049), .A(N3971) );
  INV_X1 NOT1_1172( .ZN(N4050), .A(N3977) );
  INV_X1 NOT1_1173( .ZN(N4051), .A(N3980) );
  NAND2_X1 NAND2_1174( .ZN(N4052), .A1(N3980), .A2(N3694) );
  INV_X1 NOT1_1175( .ZN(N4053), .A(N3983) );
  INV_X1 NOT1_1176( .ZN(N4054), .A(N3974) );
  NAND2_X1 NAND2_1177( .ZN(N4055), .A1(N3974), .A2(N3696) );
  AND2_X1 AND2_1178( .ZN(N4056), .A1(N3932), .A2(N2304) );
  INV_X1 NOT1_1179( .ZN(N4057), .A(N3950) );
  NAND2_X1 NAND2_1180( .ZN(N4058), .A1(N3950), .A2(N3703) );
  BUF_X1 BUFF1_1181( .Z(N4059), .A(N3937) );
  BUF_X1 BUFF1_1182( .Z(N4062), .A(N3937) );
  INV_X1 NOT1_1183( .ZN(N4065), .A(N3968) );
  NAND2_X1 NAND2_1184( .ZN(N4066), .A1(N3968), .A2(N3704) );
  BUF_X1 BUFF1_1185( .Z(N4067), .A(N3940) );
  BUF_X1 BUFF1_1186( .Z(N4070), .A(N3940) );
  NAND2_X1 NAND2_1187( .ZN(N4073), .A1(N3926), .A2(N3996) );
  INV_X1 NOT1_1188( .ZN(N4074), .A(N3992) );
  NAND2_X1 NAND2_1189( .ZN(N4075), .A1(N3493), .A2(N4042) );
  NAND2_X1 NAND2_1190( .ZN(N4076), .A1(N3499), .A2(N4045) );
  NAND2_X1 NAND2_1191( .ZN(N4077), .A1(N3505), .A2(N4048) );
  NAND2_X1 NAND2_1192( .ZN(N4078), .A1(N3511), .A2(N4049) );
  NAND2_X1 NAND2_1193( .ZN(N4079), .A1(N3517), .A2(N4050) );
  NAND2_X1 NAND2_1194( .ZN(N4080), .A1(N3523), .A2(N4053) );
  NAND2_X1 NAND2_1195( .ZN(N4085), .A1(N3496), .A2(N4043) );
  NAND2_X1 NAND2_1196( .ZN(N4086), .A1(N3502), .A2(N4046) );
  NAND2_X1 NAND2_1197( .ZN(N4088), .A1(N3520), .A2(N4051) );
  NAND2_X1 NAND2_1198( .ZN(N4090), .A1(N3514), .A2(N4054) );
  AND2_X1 AND2_1199( .ZN(N4091), .A1(N3996), .A2(N1926) );
  OR2_X1 OR2_1200( .ZN(N4094), .A1(N3605), .A2(N4056) );
  NAND2_X1 NAND2_1201( .ZN(N4098), .A1(N3490), .A2(N4057) );
  NAND2_X1 NAND2_1202( .ZN(N4101), .A1(N3508), .A2(N4065) );
  AND2_X1 AND2_1203( .ZN(N4104), .A1(N4073), .A2(N4074) );
  NAND2_X2 NAND2_1204( .ZN(N4105), .A1(N4075), .A2(N4029) );
  NAND2_X1 NAND2_1205( .ZN(N4106), .A1(N4062), .A2(N3899) );
  NAND2_X1 NAND2_1206( .ZN(N4107), .A1(N4076), .A2(N4030) );
  NAND2_X1 NAND2_1207( .ZN(N4108), .A1(N4077), .A2(N4031) );
  NAND2_X1 NAND2_1208( .ZN(N4109), .A1(N4078), .A2(N4032) );
  NAND2_X1 NAND2_1209( .ZN(N4110), .A1(N4070), .A2(N3906) );
  NAND2_X1 NAND2_1210( .ZN(N4111), .A1(N4079), .A2(N4033) );
  NAND2_X1 NAND2_1211( .ZN(N4112), .A1(N4080), .A2(N4034) );
  INV_X1 NOT1_1212( .ZN(N4113), .A(N4059) );
  NAND2_X1 NAND2_1213( .ZN(N4114), .A1(N4059), .A2(N3898) );
  INV_X1 NOT1_1214( .ZN(N4115), .A(N4062) );
  NAND2_X1 NAND2_1215( .ZN(N4116), .A1(N4085), .A2(N4044) );
  NAND2_X1 NAND2_1216( .ZN(N4119), .A1(N4086), .A2(N4047) );
  INV_X1 NOT1_1217( .ZN(N4122), .A(N4070) );
  NAND2_X1 NAND2_1218( .ZN(N4123), .A1(N4088), .A2(N4052) );
  INV_X1 NOT1_1219( .ZN(N4126), .A(N4067) );
  NAND2_X1 NAND2_1220( .ZN(N4127), .A1(N4067), .A2(N3911) );
  NAND2_X1 NAND2_1221( .ZN(N4128), .A1(N4090), .A2(N4055) );
  NAND2_X1 NAND2_1222( .ZN(N4139), .A1(N4098), .A2(N4058) );
  NAND2_X1 NAND2_1223( .ZN(N4142), .A1(N4101), .A2(N4066) );
  INV_X1 NOT1_1224( .ZN(N4145), .A(N4104) );
  INV_X1 NOT1_1225( .ZN(N4146), .A(N4105) );
  NAND2_X1 NAND2_1226( .ZN(N4147), .A1(N3824), .A2(N4115) );
  INV_X1 NOT1_1227( .ZN(N4148), .A(N4107) );
  INV_X1 NOT1_1228( .ZN(N4149), .A(N4108) );
  INV_X1 NOT1_1229( .ZN(N4150), .A(N4109) );
  NAND2_X1 NAND2_1230( .ZN(N4151), .A1(N3830), .A2(N4122) );
  INV_X1 NOT1_1231( .ZN(N4152), .A(N4111) );
  INV_X1 NOT1_1232( .ZN(N4153), .A(N4112) );
  NAND2_X1 NAND2_1233( .ZN(N4154), .A1(N3821), .A2(N4113) );
  NAND2_X1 NAND2_1234( .ZN(N4161), .A1(N3827), .A2(N4126) );
  BUF_X1 BUFF1_1235( .Z(N4167), .A(N4091) );
  BUF_X1 BUFF1_1236( .Z(N4174), .A(N4094) );
  BUF_X1 BUFF1_1237( .Z(N4182), .A(N4091) );
  AND2_X2 AND2_1238( .ZN(N4186), .A1(N330), .A2(N4094) );
  AND2_X2 AND2_1239( .ZN(N4189), .A1(N4146), .A2(N2230) );
  NAND2_X1 NAND2_1240( .ZN(N4190), .A1(N4147), .A2(N4106) );
  AND2_X1 AND2_1241( .ZN(N4191), .A1(N4148), .A2(N2232) );
  AND2_X1 AND2_1242( .ZN(N4192), .A1(N4149), .A2(N2233) );
  AND2_X1 AND2_1243( .ZN(N4193), .A1(N4150), .A2(N2234) );
  NAND2_X1 NAND2_1244( .ZN(N4194), .A1(N4151), .A2(N4110) );
  AND2_X1 AND2_1245( .ZN(N4195), .A1(N4152), .A2(N2236) );
  AND2_X1 AND2_1246( .ZN(N4196), .A1(N4153), .A2(N2237) );
  NAND2_X1 NAND2_1247( .ZN(N4197), .A1(N4154), .A2(N4114) );
  BUF_X1 BUFF1_1248( .Z(N4200), .A(N4116) );
  BUF_X1 BUFF1_1249( .Z(N4203), .A(N4116) );
  BUF_X1 BUFF1_1250( .Z(N4209), .A(N4119) );
  BUF_X1 BUFF1_1251( .Z(N4213), .A(N4119) );
  NAND2_X1 NAND2_1252( .ZN(N4218), .A1(N4161), .A2(N4127) );
  BUF_X1 BUFF1_1253( .Z(N4223), .A(N4123) );
  AND2_X1 AND2_1254( .ZN(N4238), .A1(N4128), .A2(N3917) );
  INV_X1 NOT1_1255( .ZN(N4239), .A(N4139) );
  INV_X1 NOT1_1256( .ZN(N4241), .A(N4142) );
  AND2_X1 AND2_1257( .ZN(N4242), .A1(N330), .A2(N4123) );
  BUF_X1 BUFF1_1258( .Z(N4247), .A(N4128) );
  NOR3_X1 NOR3_1259( .ZN(N4251), .A1(N3713), .A2(N4189), .A3(N2898) );
  INV_X1 NOT1_1260( .ZN(N4252), .A(N4190) );
  NOR3_X1 NOR3_1261( .ZN(N4253), .A1(N3715), .A2(N4191), .A3(N2900) );
  NOR3_X1 NOR3_1262( .ZN(N4254), .A1(N3716), .A2(N4192), .A3(N2901) );
  NOR3_X1 NOR3_1263( .ZN(N4255), .A1(N3717), .A2(N4193), .A3(N3406) );
  INV_X1 NOT1_1264( .ZN(N4256), .A(N4194) );
  NOR3_X1 NOR3_1265( .ZN(N4257), .A1(N3719), .A2(N4195), .A3(N3779) );
  NOR3_X1 NOR3_1266( .ZN(N4258), .A1(N3720), .A2(N4196), .A3(N3780) );
  AND2_X1 AND2_1267( .ZN(N4283), .A1(N4167), .A2(N4035) );
  AND2_X1 AND2_1268( .ZN(N4284), .A1(N4174), .A2(N4035) );
  OR2_X1 OR2_1269( .ZN(N4287), .A1(N3815), .A2(N4238) );
  INV_X1 NOT1_1270( .ZN(N4291), .A(N4186) );
  INV_X1 NOT1_1271( .ZN(N4295), .A(N4167) );
  BUF_X1 BUFF1_1272( .Z(N4296), .A(N4167) );
  INV_X1 NOT1_1273( .ZN(N4299), .A(N4182) );
  AND2_X1 AND2_1274( .ZN(N4303), .A1(N4252), .A2(N2231) );
  AND2_X1 AND2_1275( .ZN(N4304), .A1(N4256), .A2(N2235) );
  BUF_X1 BUFF1_1276( .Z(N4305), .A(N4197) );
  OR2_X1 OR2_1277( .ZN(N4310), .A1(N3992), .A2(N4283) );
  AND3_X1 AND3_1278( .ZN(N4316), .A1(N4174), .A2(N4213), .A3(N4203) );
  AND2_X1 AND2_1279( .ZN(N4317), .A1(N4174), .A2(N4209) );
  AND3_X1 AND3_1280( .ZN(N4318), .A1(N4223), .A2(N4128), .A3(N4218) );
  AND2_X2 AND2_1281( .ZN(N4319), .A1(N4223), .A2(N4128) );
  AND2_X2 AND2_1282( .ZN(N4322), .A1(N4167), .A2(N4209) );
  NAND2_X1 NAND2_1283( .ZN(N4325), .A1(N4203), .A2(N3913) );
  NAND3_X1 NAND3_1284( .ZN(N4326), .A1(N4203), .A2(N4213), .A3(N4167) );
  NAND2_X1 NAND2_1285( .ZN(N4327), .A1(N4218), .A2(N3815) );
  NAND3_X1 NAND3_1286( .ZN(N4328), .A1(N4218), .A2(N4128), .A3(N3917) );
  NAND2_X1 NAND2_1287( .ZN(N4329), .A1(N4247), .A2(N4013) );
  INV_X1 NOT1_1288( .ZN(N4330), .A(N4247) );
  AND3_X1 AND3_1289( .ZN(N4331), .A1(N330), .A2(N4094), .A3(N4295) );
  AND2_X1 AND2_1290( .ZN(N4335), .A1(N4251), .A2(N2730) );
  AND2_X1 AND2_1291( .ZN(N4338), .A1(N4253), .A2(N2734) );
  AND2_X1 AND2_1292( .ZN(N4341), .A1(N4254), .A2(N2736) );
  AND2_X1 AND2_1293( .ZN(N4344), .A1(N4255), .A2(N2738) );
  AND2_X1 AND2_1294( .ZN(N4347), .A1(N4257), .A2(N2742) );
  AND2_X1 AND2_1295( .ZN(N4350), .A1(N4258), .A2(N2744) );
  BUF_X1 BUFF1_1296( .Z(N4353), .A(N4197) );
  BUF_X1 BUFF1_1297( .Z(N4356), .A(N4203) );
  BUF_X1 BUFF1_1298( .Z(N4359), .A(N4209) );
  BUF_X1 BUFF1_1299( .Z(N4362), .A(N4218) );
  BUF_X1 BUFF1_1300( .Z(N4365), .A(N4242) );
  BUF_X1 BUFF1_1301( .Z(N4368), .A(N4242) );
  AND2_X1 AND2_1302( .ZN(N4371), .A1(N4223), .A2(N4223) );
  NOR3_X1 NOR3_1303( .ZN(N4376), .A1(N3714), .A2(N4303), .A3(N2899) );
  NOR3_X1 NOR3_1304( .ZN(N4377), .A1(N3718), .A2(N4304), .A3(N3642) );
  AND2_X1 AND2_1305( .ZN(N4387), .A1(N330), .A2(N4317) );
  AND2_X1 AND2_1306( .ZN(N4390), .A1(N330), .A2(N4318) );
  NAND2_X1 NAND2_1307( .ZN(N4393), .A1(N3921), .A2(N4330) );
  BUF_X1 BUFF1_1308( .Z(N4398), .A(N4287) );
  BUF_X1 BUFF1_1309( .Z(N4413), .A(N4284) );
  NAND3_X1 NAND3_1310( .ZN(N4416), .A1(N3920), .A2(N4325), .A3(N4326) );
  OR2_X1 OR2_1311( .ZN(N4421), .A1(N3812), .A2(N4322) );
  NAND3_X1 NAND3_1312( .ZN(N4427), .A1(N3948), .A2(N4327), .A3(N4328) );
  BUF_X1 BUFF1_1313( .Z(N4430), .A(N4287) );
  AND2_X1 AND2_1314( .ZN(N4435), .A1(N330), .A2(N4316) );
  OR2_X1 OR2_1315( .ZN(N4442), .A1(N4331), .A2(N4296) );
  AND4_X1 AND4_1316( .ZN(N4443), .A1(N4174), .A2(N4305), .A3(N4203), .A4(N4213) );
  NAND2_X1 NAND2_1317( .ZN(N4446), .A1(N4305), .A2(N3809) );
  NAND3_X1 NAND3_1318( .ZN(N4447), .A1(N4305), .A2(N4200), .A3(N3913) );
  NAND4_X1 NAND4_1319( .ZN(N4448), .A1(N4305), .A2(N4200), .A3(N4213), .A4(N4167) );
  INV_X1 NOT1_1320( .ZN(N4452), .A(N4356) );
  NAND2_X1 NAND2_1321( .ZN(N4458), .A1(N4329), .A2(N4393) );
  INV_X1 NOT1_1322( .ZN(N4461), .A(N4365) );
  INV_X1 NOT1_1323( .ZN(N4462), .A(N4368) );
  NAND2_X1 NAND2_1324( .ZN(N4463), .A1(N4371), .A2(N1460) );
  INV_X1 NOT1_1325( .ZN(N4464), .A(N4371) );
  BUF_X1 BUFF1_1326( .Z(N4465), .A(N4310) );
  NOR2_X1 NOR2_1327( .ZN(N4468), .A1(N4331), .A2(N4296) );
  AND2_X1 AND2_1328( .ZN(N4472), .A1(N4376), .A2(N2732) );
  AND2_X1 AND2_1329( .ZN(N4475), .A1(N4377), .A2(N2740) );
  BUF_X1 BUFF1_1330( .Z(N4479), .A(N4310) );
  INV_X1 NOT1_1331( .ZN(N4484), .A(N4353) );
  INV_X1 NOT1_1332( .ZN(N4486), .A(N4359) );
  NAND2_X1 NAND2_1333( .ZN(N4487), .A1(N4359), .A2(N4299) );
  INV_X1 NOT1_1334( .ZN(N4491), .A(N4362) );
  AND2_X1 AND2_1335( .ZN(N4493), .A1(N330), .A2(N4319) );
  INV_X1 NOT1_1336( .ZN(N4496), .A(N4398) );
  AND2_X1 AND2_1337( .ZN(N4497), .A1(N4287), .A2(N4398) );
  AND2_X1 AND2_1338( .ZN(N4498), .A1(N4442), .A2(N1769) );
  NAND4_X1 NAND4_1339( .ZN(N4503), .A1(N3947), .A2(N4446), .A3(N4447), .A4(N4448) );
  INV_X1 NOT1_1340( .ZN(N4506), .A(N4413) );
  INV_X1 NOT1_1341( .ZN(N4507), .A(N4435) );
  INV_X1 NOT1_1342( .ZN(N4508), .A(N4421) );
  NAND2_X2 NAND2_1343( .ZN(N4509), .A1(N4421), .A2(N4452) );
  INV_X1 NOT1_1344( .ZN(N4510), .A(N4427) );
  NAND2_X2 NAND2_1345( .ZN(N4511), .A1(N4427), .A2(N4241) );
  NAND2_X2 NAND2_1346( .ZN(N4515), .A1(N965), .A2(N4464) );
  INV_X1 NOT1_1347( .ZN(N4526), .A(N4416) );
  NAND2_X1 NAND2_1348( .ZN(N4527), .A1(N4416), .A2(N4484) );
  NAND2_X1 NAND2_1349( .ZN(N4528), .A1(N4182), .A2(N4486) );
  INV_X1 NOT1_1350( .ZN(N4529), .A(N4430) );
  NAND2_X1 NAND2_1351( .ZN(N4530), .A1(N4430), .A2(N4491) );
  BUF_X1 BUFF1_1352( .Z(N4531), .A(N4387) );
  BUF_X1 BUFF1_1353( .Z(N4534), .A(N4387) );
  BUF_X1 BUFF1_1354( .Z(N4537), .A(N4390) );
  BUF_X1 BUFF1_1355( .Z(N4540), .A(N4390) );
  AND3_X1 AND3_1356( .ZN(N4545), .A1(N330), .A2(N4319), .A3(N4496) );
  AND2_X1 AND2_1357( .ZN(N4549), .A1(N330), .A2(N4443) );
  NAND2_X1 NAND2_1358( .ZN(N4552), .A1(N4356), .A2(N4508) );
  NAND2_X1 NAND2_1359( .ZN(N4555), .A1(N4142), .A2(N4510) );
  INV_X1 NOT1_1360( .ZN(N4558), .A(N4493) );
  NAND2_X1 NAND2_1361( .ZN(N4559), .A1(N4463), .A2(N4515) );
  INV_X1 NOT1_1362( .ZN(N4562), .A(N4465) );
  AND2_X1 AND2_1363( .ZN(N4563), .A1(N4310), .A2(N4465) );
  BUF_X1 BUFF1_1364( .Z(N4564), .A(N4468) );
  INV_X1 NOT1_1365( .ZN(N4568), .A(N4479) );
  BUF_X1 BUFF1_1366( .Z(N4569), .A(N4443) );
  NAND2_X1 NAND2_1367( .ZN(N4572), .A1(N4353), .A2(N4526) );
  NAND2_X1 NAND2_1368( .ZN(N4573), .A1(N4362), .A2(N4529) );
  NAND2_X1 NAND2_1369( .ZN(N4576), .A1(N4487), .A2(N4528) );
  BUF_X1 BUFF1_1370( .Z(N4581), .A(N4458) );
  BUF_X1 BUFF1_1371( .Z(N4584), .A(N4458) );
  OR3_X1 OR3_1372( .ZN(N4587), .A1(N2758), .A2(N4498), .A3(N2761) );
  NOR3_X1 NOR3_1373( .ZN(N4588), .A1(N2758), .A2(N4498), .A3(N2761) );
  OR2_X1 OR2_1374( .ZN(N4589), .A1(N4545), .A2(N4497) );
  NAND2_X1 NAND2_1375( .ZN(N4593), .A1(N4552), .A2(N4509) );
  INV_X1 NOT1_1376( .ZN(N4596), .A(N4531) );
  INV_X1 NOT1_1377( .ZN(N4597), .A(N4534) );
  NAND2_X1 NAND2_1378( .ZN(N4599), .A1(N4555), .A2(N4511) );
  INV_X1 NOT1_1379( .ZN(N4602), .A(N4537) );
  INV_X1 NOT1_1380( .ZN(N4603), .A(N4540) );
  AND3_X1 AND3_1381( .ZN(N4608), .A1(N330), .A2(N4284), .A3(N4562) );
  BUF_X1 BUFF1_1382( .Z(N4613), .A(N4503) );
  BUF_X1 BUFF1_1383( .Z(N4616), .A(N4503) );
  NAND2_X1 NAND2_1384( .ZN(N4619), .A1(N4572), .A2(N4527) );
  NAND2_X1 NAND2_1385( .ZN(N4623), .A1(N4573), .A2(N4530) );
  INV_X1 NOT1_1386( .ZN(N4628), .A(N4588) );
  NAND2_X1 NAND2_1387( .ZN(N4629), .A1(N4569), .A2(N4506) );
  INV_X1 NOT1_1388( .ZN(N4630), .A(N4569) );
  INV_X1 NOT1_1389( .ZN(N4635), .A(N4576) );
  NAND2_X1 NAND2_1390( .ZN(N4636), .A1(N4576), .A2(N4291) );
  INV_X1 NOT1_1391( .ZN(N4640), .A(N4581) );
  NAND2_X1 NAND2_1392( .ZN(N4641), .A1(N4581), .A2(N4461) );
  INV_X1 NOT1_1393( .ZN(N4642), .A(N4584) );
  NAND2_X1 NAND2_1394( .ZN(N4643), .A1(N4584), .A2(N4462) );
  NOR2_X1 NOR2_1395( .ZN(N4644), .A1(N4608), .A2(N4563) );
  AND2_X1 AND2_1396( .ZN(N4647), .A1(N4559), .A2(N2128) );
  AND2_X1 AND2_1397( .ZN(N4650), .A1(N4559), .A2(N2743) );
  BUF_X1 BUFF1_1398( .Z(N4656), .A(N4549) );
  BUF_X1 BUFF1_1399( .Z(N4659), .A(N4549) );
  BUF_X1 BUFF1_1400( .Z(N4664), .A(N4564) );
  AND2_X1 AND2_1401( .ZN(N4667), .A1(N4587), .A2(N4628) );
  NAND2_X2 NAND2_1402( .ZN(N4668), .A1(N4413), .A2(N4630) );
  INV_X1 NOT1_1403( .ZN(N4669), .A(N4616) );
  NAND2_X2 NAND2_1404( .ZN(N4670), .A1(N4616), .A2(N4239) );
  INV_X1 NOT1_1405( .ZN(N4673), .A(N4619) );
  NAND2_X1 NAND2_1406( .ZN(N4674), .A1(N4619), .A2(N4507) );
  NAND2_X1 NAND2_1407( .ZN(N4675), .A1(N4186), .A2(N4635) );
  INV_X1 NOT1_1408( .ZN(N4676), .A(N4623) );
  NAND2_X1 NAND2_1409( .ZN(N4677), .A1(N4623), .A2(N4558) );
  NAND2_X1 NAND2_1410( .ZN(N4678), .A1(N4365), .A2(N4640) );
  NAND2_X1 NAND2_1411( .ZN(N4679), .A1(N4368), .A2(N4642) );
  INV_X1 NOT1_1412( .ZN(N4687), .A(N4613) );
  NAND2_X1 NAND2_1413( .ZN(N4688), .A1(N4613), .A2(N4568) );
  BUF_X1 BUFF1_1414( .Z(N4691), .A(N4593) );
  BUF_X1 BUFF1_1415( .Z(N4694), .A(N4593) );
  BUF_X1 BUFF1_1416( .Z(N4697), .A(N4599) );
  BUF_X1 BUFF1_1417( .Z(N4700), .A(N4599) );
  NAND2_X1 NAND2_1418( .ZN(N4704), .A1(N4629), .A2(N4668) );
  NAND2_X1 NAND2_1419( .ZN(N4705), .A1(N4139), .A2(N4669) );
  INV_X1 NOT1_1420( .ZN(N4706), .A(N4656) );
  INV_X1 NOT1_1421( .ZN(N4707), .A(N4659) );
  NAND2_X1 NAND2_1422( .ZN(N4708), .A1(N4435), .A2(N4673) );
  NAND2_X1 NAND2_1423( .ZN(N4711), .A1(N4675), .A2(N4636) );
  NAND2_X1 NAND2_1424( .ZN(N4716), .A1(N4493), .A2(N4676) );
  NAND2_X1 NAND2_1425( .ZN(N4717), .A1(N4678), .A2(N4641) );
  NAND2_X1 NAND2_1426( .ZN(N4721), .A1(N4679), .A2(N4643) );
  BUF_X1 BUFF1_1427( .Z(N4722), .A(N4644) );
  INV_X1 NOT1_1428( .ZN(N4726), .A(N4664) );
  OR3_X1 OR3_1429( .ZN(N4727), .A1(N4647), .A2(N4650), .A3(N4350) );
  NOR3_X1 NOR3_1430( .ZN(N4730), .A1(N4647), .A2(N4650), .A3(N4350) );
  NAND2_X1 NAND2_1431( .ZN(N4733), .A1(N4479), .A2(N4687) );
  NAND2_X1 NAND2_1432( .ZN(N4740), .A1(N4705), .A2(N4670) );
  NAND2_X1 NAND2_1433( .ZN(N4743), .A1(N4708), .A2(N4674) );
  INV_X1 NOT1_1434( .ZN(N4747), .A(N4691) );
  NAND2_X1 NAND2_1435( .ZN(N4748), .A1(N4691), .A2(N4596) );
  INV_X1 NOT1_1436( .ZN(N4749), .A(N4694) );
  NAND2_X1 NAND2_1437( .ZN(N4750), .A1(N4694), .A2(N4597) );
  INV_X1 NOT1_1438( .ZN(N4753), .A(N4697) );
  NAND2_X1 NAND2_1439( .ZN(N4754), .A1(N4697), .A2(N4602) );
  INV_X1 NOT1_1440( .ZN(N4755), .A(N4700) );
  NAND2_X1 NAND2_1441( .ZN(N4756), .A1(N4700), .A2(N4603) );
  NAND2_X1 NAND2_1442( .ZN(N4757), .A1(N4716), .A2(N4677) );
  NAND2_X1 NAND2_1443( .ZN(N4769), .A1(N4733), .A2(N4688) );
  AND2_X1 AND2_1444( .ZN(N4772), .A1(N330), .A2(N4704) );
  INV_X1 NOT1_1445( .ZN(N4775), .A(N4721) );
  INV_X1 NOT1_1446( .ZN(N4778), .A(N4730) );
  NAND2_X1 NAND2_1447( .ZN(N4786), .A1(N4531), .A2(N4747) );
  NAND2_X1 NAND2_1448( .ZN(N4787), .A1(N4534), .A2(N4749) );
  NAND2_X1 NAND2_1449( .ZN(N4788), .A1(N4537), .A2(N4753) );
  NAND2_X1 NAND2_1450( .ZN(N4789), .A1(N4540), .A2(N4755) );
  AND2_X1 AND2_1451( .ZN(N4794), .A1(N4711), .A2(N2124) );
  AND2_X1 AND2_1452( .ZN(N4797), .A1(N4711), .A2(N2735) );
  AND2_X1 AND2_1453( .ZN(N4800), .A1(N4717), .A2(N2127) );
  BUF_X1 BUFF1_1454( .Z(N4805), .A(N4722) );
  AND2_X1 AND2_1455( .ZN(N4808), .A1(N4717), .A2(N4468) );
  BUF_X1 BUFF1_1456( .Z(N4812), .A(N4727) );
  AND2_X1 AND2_1457( .ZN(N4815), .A1(N4727), .A2(N4778) );
  INV_X1 NOT1_1458( .ZN(N4816), .A(N4769) );
  INV_X1 NOT1_1459( .ZN(N4817), .A(N4772) );
  NAND2_X1 NAND2_1460( .ZN(N4818), .A1(N4786), .A2(N4748) );
  NAND2_X1 NAND2_1461( .ZN(N4822), .A1(N4787), .A2(N4750) );
  NAND2_X1 NAND2_1462( .ZN(N4823), .A1(N4788), .A2(N4754) );
  NAND2_X1 NAND2_1463( .ZN(N4826), .A1(N4789), .A2(N4756) );
  NAND2_X1 NAND2_1464( .ZN(N4829), .A1(N4775), .A2(N4726) );
  INV_X1 NOT1_1465( .ZN(N4830), .A(N4775) );
  AND2_X1 AND2_1466( .ZN(N4831), .A1(N4743), .A2(N2122) );
  AND2_X1 AND2_1467( .ZN(N4838), .A1(N4757), .A2(N2126) );
  BUF_X1 BUFF1_1468( .Z(N4844), .A(N4740) );
  BUF_X1 BUFF1_1469( .Z(N4847), .A(N4740) );
  BUF_X1 BUFF1_1470( .Z(N4850), .A(N4743) );
  BUF_X1 BUFF1_1471( .Z(N4854), .A(N4757) );
  NAND2_X1 NAND2_1472( .ZN(N4859), .A1(N4772), .A2(N4816) );
  NAND2_X1 NAND2_1473( .ZN(N4860), .A1(N4769), .A2(N4817) );
  INV_X1 NOT1_1474( .ZN(N4868), .A(N4826) );
  INV_X1 NOT1_1475( .ZN(N4870), .A(N4805) );
  INV_X1 NOT1_1476( .ZN(N4872), .A(N4808) );
  NAND2_X1 NAND2_1477( .ZN(N4873), .A1(N4664), .A2(N4830) );
  OR3_X1 OR3_1478( .ZN(N4876), .A1(N4794), .A2(N4797), .A3(N4341) );
  NOR3_X1 NOR3_1479( .ZN(N4880), .A1(N4794), .A2(N4797), .A3(N4341) );
  INV_X1 NOT1_1480( .ZN(N4885), .A(N4812) );
  INV_X1 NOT1_1481( .ZN(N4889), .A(N4822) );
  NAND2_X1 NAND2_1482( .ZN(N4895), .A1(N4859), .A2(N4860) );
  INV_X1 NOT1_1483( .ZN(N4896), .A(N4844) );
  NAND2_X1 NAND2_1484( .ZN(N4897), .A1(N4844), .A2(N4706) );
  INV_X1 NOT1_1485( .ZN(N4898), .A(N4847) );
  NAND2_X1 NAND2_1486( .ZN(N4899), .A1(N4847), .A2(N4707) );
  NOR2_X1 NOR2_1487( .ZN(N4900), .A1(N4868), .A2(N4564) );
  AND4_X1 AND4_1488( .ZN(N4901), .A1(N4717), .A2(N4757), .A3(N4823), .A4(N4564) );
  INV_X1 NOT1_1489( .ZN(N4902), .A(N4850) );
  INV_X1 NOT1_1490( .ZN(N4904), .A(N4854) );
  NAND2_X1 NAND2_1491( .ZN(N4905), .A1(N4854), .A2(N4872) );
  NAND2_X1 NAND2_1492( .ZN(N4906), .A1(N4873), .A2(N4829) );
  AND2_X1 AND2_1493( .ZN(N4907), .A1(N4818), .A2(N2123) );
  AND2_X1 AND2_1494( .ZN(N4913), .A1(N4823), .A2(N2125) );
  AND2_X1 AND2_1495( .ZN(N4916), .A1(N4818), .A2(N4644) );
  INV_X1 NOT1_1496( .ZN(N4920), .A(N4880) );
  AND2_X1 AND2_1497( .ZN(N4921), .A1(N4895), .A2(N2184) );
  NAND2_X1 NAND2_1498( .ZN(N4924), .A1(N4656), .A2(N4896) );
  NAND2_X1 NAND2_1499( .ZN(N4925), .A1(N4659), .A2(N4898) );
  OR2_X1 OR2_1500( .ZN(N4926), .A1(N4900), .A2(N4901) );
  NAND2_X1 NAND2_1501( .ZN(N4928), .A1(N4889), .A2(N4870) );
  INV_X1 NOT1_1502( .ZN(N4929), .A(N4889) );
  NAND2_X1 NAND2_1503( .ZN(N4930), .A1(N4808), .A2(N4904) );
  INV_X1 NOT1_1504( .ZN(N4931), .A(N4906) );
  BUF_X1 BUFF1_1505( .Z(N4937), .A(N4876) );
  BUF_X1 BUFF1_1506( .Z(N4940), .A(N4876) );
  AND2_X1 AND2_1507( .ZN(N4944), .A1(N4876), .A2(N4920) );
  NAND2_X1 NAND2_1508( .ZN(N4946), .A1(N4924), .A2(N4897) );
  NAND2_X1 NAND2_1509( .ZN(N4949), .A1(N4925), .A2(N4899) );
  NAND2_X1 NAND2_1510( .ZN(N4950), .A1(N4916), .A2(N4902) );
  INV_X1 NOT1_1511( .ZN(N4951), .A(N4916) );
  NAND2_X1 NAND2_1512( .ZN(N4952), .A1(N4805), .A2(N4929) );
  NAND2_X1 NAND2_1513( .ZN(N4953), .A1(N4930), .A2(N4905) );
  AND2_X1 AND2_1514( .ZN(N4954), .A1(N4926), .A2(N2737) );
  AND2_X1 AND2_1515( .ZN(N4957), .A1(N4931), .A2(N2741) );
  OR3_X1 OR3_1516( .ZN(N4964), .A1(N2764), .A2(N2483), .A3(N4921) );
  NOR3_X1 NOR3_1517( .ZN(N4965), .A1(N2764), .A2(N2483), .A3(N4921) );
  INV_X1 NOT1_1518( .ZN(N4968), .A(N4949) );
  NAND2_X1 NAND2_1519( .ZN(N4969), .A1(N4850), .A2(N4951) );
  NAND2_X1 NAND2_1520( .ZN(N4970), .A1(N4952), .A2(N4928) );
  AND2_X1 AND2_1521( .ZN(N4973), .A1(N4953), .A2(N2739) );
  INV_X1 NOT1_1522( .ZN(N4978), .A(N4937) );
  INV_X1 NOT1_1523( .ZN(N4979), .A(N4940) );
  INV_X1 NOT1_1524( .ZN(N4980), .A(N4965) );
  NOR2_X1 NOR2_1525( .ZN(N4981), .A1(N4968), .A2(N4722) );
  AND4_X1 AND4_1526( .ZN(N4982), .A1(N4818), .A2(N4743), .A3(N4946), .A4(N4722) );
  NAND2_X1 NAND2_1527( .ZN(N4983), .A1(N4950), .A2(N4969) );
  INV_X1 NOT1_1528( .ZN(N4984), .A(N4970) );
  AND2_X1 AND2_1529( .ZN(N4985), .A1(N4946), .A2(N2121) );
  OR3_X1 OR3_1530( .ZN(N4988), .A1(N4913), .A2(N4954), .A3(N4344) );
  NOR3_X1 NOR3_1531( .ZN(N4991), .A1(N4913), .A2(N4954), .A3(N4344) );
  OR3_X1 OR3_1532( .ZN(N4996), .A1(N4800), .A2(N4957), .A3(N4347) );
  NOR3_X1 NOR3_1533( .ZN(N4999), .A1(N4800), .A2(N4957), .A3(N4347) );
  AND2_X1 AND2_1534( .ZN(N5002), .A1(N4964), .A2(N4980) );
  OR2_X1 OR2_1535( .ZN(N5007), .A1(N4981), .A2(N4982) );
  AND2_X1 AND2_1536( .ZN(N5010), .A1(N4983), .A2(N2731) );
  AND2_X1 AND2_1537( .ZN(N5013), .A1(N4984), .A2(N2733) );
  OR3_X1 OR3_1538( .ZN(N5018), .A1(N4838), .A2(N4973), .A3(N4475) );
  NOR3_X1 NOR3_1539( .ZN(N5021), .A1(N4838), .A2(N4973), .A3(N4475) );
  INV_X1 NOT1_1540( .ZN(N5026), .A(N4991) );
  INV_X1 NOT1_1541( .ZN(N5029), .A(N4999) );
  AND2_X1 AND2_1542( .ZN(N5030), .A1(N5007), .A2(N2729) );
  BUF_X1 BUFF1_1543( .Z(N5039), .A(N4996) );
  BUF_X1 BUFF1_1544( .Z(N5042), .A(N4988) );
  AND2_X1 AND2_1545( .ZN(N5045), .A1(N4988), .A2(N5026) );
  INV_X1 NOT1_1546( .ZN(N5046), .A(N5021) );
  AND2_X1 AND2_1547( .ZN(N5047), .A1(N4996), .A2(N5029) );
  OR3_X1 OR3_1548( .ZN(N5050), .A1(N4831), .A2(N5010), .A3(N4472) );
  NOR3_X1 NOR3_1549( .ZN(N5055), .A1(N4831), .A2(N5010), .A3(N4472) );
  OR3_X1 OR3_1550( .ZN(N5058), .A1(N4907), .A2(N5013), .A3(N4338) );
  NOR3_X1 NOR3_1551( .ZN(N5061), .A1(N4907), .A2(N5013), .A3(N4338) );
  AND4_X1 AND4_1552( .ZN(N5066), .A1(N4730), .A2(N4999), .A3(N5021), .A4(N4991) );
  BUF_X1 BUFF1_1553( .Z(N5070), .A(N5018) );
  AND2_X1 AND2_1554( .ZN(N5078), .A1(N5018), .A2(N5046) );
  OR3_X1 OR3_1555( .ZN(N5080), .A1(N4985), .A2(N5030), .A3(N4335) );
  NOR3_X1 NOR3_1556( .ZN(N5085), .A1(N4985), .A2(N5030), .A3(N4335) );
  NAND2_X1 NAND2_1557( .ZN(N5094), .A1(N5039), .A2(N4885) );
  INV_X1 NOT1_1558( .ZN(N5095), .A(N5039) );
  INV_X1 NOT1_1559( .ZN(N5097), .A(N5042) );
  AND2_X1 AND2_1560( .ZN(N5102), .A1(N5050), .A2(N5050) );
  INV_X1 NOT1_1561( .ZN(N5103), .A(N5061) );
  NAND2_X1 NAND2_1562( .ZN(N5108), .A1(N4812), .A2(N5095) );
  INV_X1 NOT1_1563( .ZN(N5109), .A(N5070) );
  NAND2_X1 NAND2_1564( .ZN(N5110), .A1(N5070), .A2(N5097) );
  BUF_X1 BUFF1_1565( .Z(N5111), .A(N5058) );
  AND2_X1 AND2_1566( .ZN(N5114), .A1(N5050), .A2(N1461) );
  BUF_X1 BUFF1_1567( .Z(N5117), .A(N5050) );
  AND2_X1 AND2_1568( .ZN(N5120), .A1(N5080), .A2(N5080) );
  AND2_X1 AND2_1569( .ZN(N5121), .A1(N5058), .A2(N5103) );
  NAND2_X1 NAND2_1570( .ZN(N5122), .A1(N5094), .A2(N5108) );
  NAND2_X1 NAND2_1571( .ZN(N5125), .A1(N5042), .A2(N5109) );
  AND2_X1 AND2_1572( .ZN(N5128), .A1(N1461), .A2(N5080) );
  AND4_X1 AND4_1573( .ZN(N5133), .A1(N4880), .A2(N5061), .A3(N5055), .A4(N5085) );
  AND3_X1 AND3_1574( .ZN(N5136), .A1(N5055), .A2(N5085), .A3(N1464) );
  BUF_X1 BUFF1_1575( .Z(N5139), .A(N5080) );
  NAND2_X1 NAND2_1576( .ZN(N5145), .A1(N5125), .A2(N5110) );
  BUF_X1 BUFF1_1577( .Z(N5151), .A(N5111) );
  BUF_X1 BUFF1_1578( .Z(N5154), .A(N5111) );
  INV_X1 NOT1_1579( .ZN(N5159), .A(N5117) );
  BUF_X1 BUFF1_1580( .Z(N5160), .A(N5114) );
  BUF_X1 BUFF1_1581( .Z(N5163), .A(N5114) );
  AND2_X1 AND2_1582( .ZN(N5166), .A1(N5066), .A2(N5133) );
  AND2_X1 AND2_1583( .ZN(N5173), .A1(N5066), .A2(N5133) );
  BUF_X1 BUFF1_1584( .Z(N5174), .A(N5122) );
  BUF_X1 BUFF1_1585( .Z(N5177), .A(N5122) );
  INV_X1 NOT1_1586( .ZN(N5182), .A(N5139) );
  NAND2_X1 NAND2_1587( .ZN(N5183), .A1(N5139), .A2(N5159) );
  BUF_X1 BUFF1_1588( .Z(N5184), .A(N5128) );
  BUF_X1 BUFF1_1589( .Z(N5188), .A(N5128) );
  INV_X1 NOT1_1590( .ZN(N5192), .A(N5166) );
  NOR2_X1 NOR2_1591( .ZN(N5193), .A1(N5136), .A2(N5173) );
  NAND2_X1 NAND2_1592( .ZN(N5196), .A1(N5151), .A2(N4978) );
  INV_X1 NOT1_1593( .ZN(N5197), .A(N5151) );
  NAND2_X1 NAND2_1594( .ZN(N5198), .A1(N5154), .A2(N4979) );
  INV_X1 NOT1_1595( .ZN(N5199), .A(N5154) );
  INV_X1 NOT1_1596( .ZN(N5201), .A(N5160) );
  INV_X1 NOT1_1597( .ZN(N5203), .A(N5163) );
  BUF_X1 BUFF1_1598( .Z(N5205), .A(N5145) );
  BUF_X1 BUFF1_1599( .Z(N5209), .A(N5145) );
  NAND2_X1 NAND2_1600( .ZN(N5212), .A1(N5117), .A2(N5182) );
  AND2_X1 AND2_1601( .ZN(N5215), .A1(N213), .A2(N5193) );
  INV_X1 NOT1_1602( .ZN(N5217), .A(N5174) );
  INV_X1 NOT1_1603( .ZN(N5219), .A(N5177) );
  NAND2_X1 NAND2_1604( .ZN(N5220), .A1(N4937), .A2(N5197) );
  NAND2_X1 NAND2_1605( .ZN(N5221), .A1(N4940), .A2(N5199) );
  INV_X1 NOT1_1606( .ZN(N5222), .A(N5184) );
  NAND2_X1 NAND2_1607( .ZN(N5223), .A1(N5184), .A2(N5201) );
  NAND2_X1 NAND2_1608( .ZN(N5224), .A1(N5188), .A2(N5203) );
  INV_X1 NOT1_1609( .ZN(N5225), .A(N5188) );
  NAND2_X1 NAND2_1610( .ZN(N5228), .A1(N5183), .A2(N5212) );
  INV_X1 NOT1_1611( .ZN(N5231), .A(N5215) );
  NAND2_X1 NAND2_1612( .ZN(N5232), .A1(N5205), .A2(N5217) );
  INV_X1 NOT1_1613( .ZN(N5233), .A(N5205) );
  NAND2_X1 NAND2_1614( .ZN(N5234), .A1(N5209), .A2(N5219) );
  INV_X1 NOT1_1615( .ZN(N5235), .A(N5209) );
  NAND2_X1 NAND2_1616( .ZN(N5236), .A1(N5196), .A2(N5220) );
  NAND2_X1 NAND2_1617( .ZN(N5240), .A1(N5198), .A2(N5221) );
  NAND2_X1 NAND2_1618( .ZN(N5242), .A1(N5160), .A2(N5222) );
  NAND2_X1 NAND2_1619( .ZN(N5243), .A1(N5163), .A2(N5225) );
  NAND2_X1 NAND2_1620( .ZN(N5245), .A1(N5174), .A2(N5233) );
  NAND2_X2 NAND2_1621( .ZN(N5246), .A1(N5177), .A2(N5235) );
  INV_X1 NOT1_1622( .ZN(N5250), .A(N5240) );
  INV_X1 NOT1_1623( .ZN(N5253), .A(N5228) );
  NAND2_X1 NAND2_1624( .ZN(N5254), .A1(N5242), .A2(N5223) );
  NAND2_X1 NAND2_1625( .ZN(N5257), .A1(N5243), .A2(N5224) );
  NAND2_X1 NAND2_1626( .ZN(N5258), .A1(N5232), .A2(N5245) );
  NAND2_X1 NAND2_1627( .ZN(N5261), .A1(N5234), .A2(N5246) );
  INV_X1 NOT1_1628( .ZN(N5266), .A(N5257) );
  BUF_X1 BUFF1_1629( .Z(N5269), .A(N5236) );
  AND3_X1 AND3_1630( .ZN(N5277), .A1(N5236), .A2(N5254), .A3(N2307) );
  AND3_X1 AND3_1631( .ZN(N5278), .A1(N5250), .A2(N5254), .A3(N2310) );
  INV_X1 NOT1_1632( .ZN(N5279), .A(N5261) );
  INV_X1 NOT1_1633( .ZN(N5283), .A(N5269) );
  NAND2_X1 NAND2_1634( .ZN(N5284), .A1(N5269), .A2(N5253) );
  AND3_X1 AND3_1635( .ZN(N5285), .A1(N5236), .A2(N5266), .A3(N2310) );
  AND3_X1 AND3_1636( .ZN(N5286), .A1(N5250), .A2(N5266), .A3(N2307) );
  BUF_X1 BUFF1_1637( .Z(N5289), .A(N5258) );
  BUF_X1 BUFF1_1638( .Z(N5292), .A(N5258) );
  NAND2_X1 NAND2_1639( .ZN(N5295), .A1(N5228), .A2(N5283) );
  OR4_X1 OR4_1640( .ZN(N5298), .A1(N5277), .A2(N5285), .A3(N5278), .A4(N5286) );
  BUF_X1 BUFF1_1641( .Z(N5303), .A(N5279) );
  BUF_X1 BUFF1_1642( .Z(N5306), .A(N5279) );
  NAND2_X1 NAND2_1643( .ZN(N5309), .A1(N5295), .A2(N5284) );
  INV_X1 NOT1_1644( .ZN(N5312), .A(N5292) );
  INV_X1 NOT1_1645( .ZN(N5313), .A(N5289) );
  INV_X1 NOT1_1646( .ZN(N5322), .A(N5306) );
  INV_X1 NOT1_1647( .ZN(N5323), .A(N5303) );
  BUF_X1 BUFF1_1648( .Z(N5324), .A(N5298) );
  BUF_X1 BUFF1_1649( .Z(N5327), .A(N5298) );
  BUF_X1 BUFF1_1650( .Z(N5332), .A(N5309) );
  BUF_X1 BUFF1_1651( .Z(N5335), .A(N5309) );
  NAND2_X1 NAND2_1652( .ZN(N5340), .A1(N5324), .A2(N5323) );
  NAND2_X1 NAND2_1653( .ZN(N5341), .A1(N5327), .A2(N5322) );
  INV_X1 NOT1_1654( .ZN(N5344), .A(N5327) );
  INV_X1 NOT1_1655( .ZN(N5345), .A(N5324) );
  NAND2_X1 NAND2_1656( .ZN(N5348), .A1(N5332), .A2(N5313) );
  NAND2_X1 NAND2_1657( .ZN(N5349), .A1(N5335), .A2(N5312) );
  NAND2_X1 NAND2_1658( .ZN(N5350), .A1(N5303), .A2(N5345) );
  NAND2_X1 NAND2_1659( .ZN(N5351), .A1(N5306), .A2(N5344) );
  INV_X1 NOT1_1660( .ZN(N5352), .A(N5335) );
  INV_X1 NOT1_1661( .ZN(N5353), .A(N5332) );
  NAND2_X1 NAND2_1662( .ZN(N5354), .A1(N5289), .A2(N5353) );
  NAND2_X1 NAND2_1663( .ZN(N5355), .A1(N5292), .A2(N5352) );
  NAND2_X1 NAND2_1664( .ZN(N5356), .A1(N5350), .A2(N5340) );
  NAND2_X1 NAND2_1665( .ZN(N5357), .A1(N5351), .A2(N5341) );
  NAND2_X1 NAND2_1666( .ZN(N5358), .A1(N5348), .A2(N5354) );
  NAND2_X1 NAND2_1667( .ZN(N5359), .A1(N5349), .A2(N5355) );
  AND2_X1 AND2_1668( .ZN(N5360), .A1(N5356), .A2(N5357) );
  NAND2_X1 NAND2_1669( .ZN(N5361), .A1(N5358), .A2(N5359) );

endmodule
