// Verilog
// c5315
// Ninputs 178
// Noutputs 123
// NtotalGates 2307
// BUFF1 313
// AND2 319
// NOT1 581
// NAND2 454
// AND4 27
// OR2 95
// AND3 359
// OR3 50
// OR4 61
// NOR2 19
// AND5 11
// OR5 8
// NOR3 6
// NOR4 2
// AND9 2

module c5315(N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,N27,N31,N34,N37,N40,N43,N46,N49,
  N52,N53,N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,N82,N83,N86,N87,N88,N91,
  N94,N97,N100,N103,N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,
  N126,N127,N128,N129,N130,N131,N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,N155,N158,
  N161,N164,N167,N170,N173,N176,N179,N182,N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,
  N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,N251,N254,N257,N264,N265,N272,N273,N280,
  N281,N288,N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,N324,N331,N332,N335,N338,N341,
  N348,N351,N358,N361,N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,N435,N446,N457,N468,
  N479,N490,N503,N514,N523,N534,N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,N580,N583,
  N588,N591,N592,N595,N596,N597,N598,N599,N603,N607,N610,N613,N616,N619,N625,N631,N709,N816,
  N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,
  N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,
  N4279,N4737,N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,N6925,N6926,N6927,N7015,
  N7363,N7365,N7432,N7449,N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,N7506,N7511,
  N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,
  N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,
  N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,N8124,N8127,N8128);
input N1,N4,N11,N14,N17,N20,N23,N24,N25,N26,N27,N31,N34,N37,N40,N43,N46,N49,N52,N53,
  N54,N61,N64,N67,N70,N73,N76,N79,N80,N81,N82,N83,N86,N87,N88,N91,N94,N97,N100,N103,
  N106,N109,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N126,N127,N128,N129,N130,N131,
  N132,N135,N136,N137,N140,N141,N145,N146,N149,N152,N155,N158,N161,N164,N167,N170,N173,N176,N179,N182,
  N185,N188,N191,N194,N197,N200,N203,N206,N209,N210,N217,N218,N225,N226,N233,N234,N241,N242,N245,N248,
  N251,N254,N257,N264,N265,N272,N273,N280,N281,N288,N289,N292,N293,N299,N302,N307,N308,N315,N316,N323,
  N324,N331,N332,N335,N338,N341,N348,N351,N358,N361,N366,N369,N372,N373,N374,N386,N389,N400,N411,N422,
  N435,N446,N457,N468,N479,N490,N503,N514,N523,N534,N545,N549,N552,N556,N559,N562,N566,N571,N574,N577,
  N580,N583,N588,N591,N592,N595,N596,N597,N598,N599,N603,N607,N610,N613,N616,N619,N625,N631;
output N709,N816,N1066,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1147,N1152,N1153,N1154,N1155,N1972,N2054,N2060,
  N2061,N2139,N2142,N2309,N2387,N2527,N2584,N2590,N2623,N3357,N3358,N3359,N3360,N3604,N3613,N4272,N4275,N4278,N4279,N4737,
  N4738,N4739,N4740,N5240,N5388,N6641,N6643,N6646,N6648,N6716,N6877,N6924,N6925,N6926,N6927,N7015,N7363,N7365,N7432,N7449,
  N7465,N7466,N7467,N7469,N7470,N7471,N7472,N7473,N7474,N7476,N7503,N7504,N7506,N7511,N7515,N7516,N7517,N7518,N7519,N7520,
  N7521,N7522,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7626,N7698,N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,
  N7707,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N8075,N8076,N8123,
  N8124,N8127,N8128;

  wire N1042,N1043,N1067,N1080,N1092,N1104,N1146,N1148,N1149,N1150,N1151,N1156,N1157,N1161,N1173,N1185,
    N1197,N1209,N1213,N1216,N1219,N1223,N1235,N1247,N1259,N1271,N1280,N1292,N1303,N1315,N1327,N1339,
    N1351,N1363,N1375,N1378,N1381,N1384,N1387,N1390,N1393,N1396,N1415,N1418,N1421,N1424,N1427,N1430,
    N1433,N1436,N1455,N1462,N1469,N1475,N1479,N1482,N1492,N1495,N1498,N1501,N1504,N1507,N1510,N1513,
    N1516,N1519,N1522,N1525,N1542,N1545,N1548,N1551,N1554,N1557,N1560,N1563,N1566,N1573,N1580,N1583,
    N1588,N1594,N1597,N1600,N1603,N1606,N1609,N1612,N1615,N1618,N1621,N1624,N1627,N1630,N1633,N1636,
    N1639,N1642,N1645,N1648,N1651,N1654,N1657,N1660,N1663,N1675,N1685,N1697,N1709,N1721,N1727,N1731,
    N1743,N1755,N1758,N1761,N1769,N1777,N1785,N1793,N1800,N1807,N1814,N1821,N1824,N1827,N1830,N1833,
    N1836,N1839,N1842,N1845,N1848,N1851,N1854,N1857,N1860,N1863,N1866,N1869,N1872,N1875,N1878,N1881,
    N1884,N1887,N1890,N1893,N1896,N1899,N1902,N1905,N1908,N1911,N1914,N1917,N1920,N1923,N1926,N1929,
    N1932,N1935,N1938,N1941,N1944,N1947,N1950,N1953,N1956,N1959,N1962,N1965,N1968,N2349,N2350,N2585,
    N2586,N2587,N2588,N2589,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,
    N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
    N2619,N2620,N2621,N2622,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,
    N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2653,N2664,N2675,N2681,
    N2692,N2703,N2704,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,
    N2722,N2728,N2739,N2750,N2756,N2767,N2778,N2779,N2790,N2801,N2812,N2823,N2824,N2825,N2826,N2827,
    N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,
    N2844,N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2861,N2867,N2868,N2869,
    N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2882,N2891,N2901,N2902,N2903,N2904,N2905,N2906,
    N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,
    N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
    N2939,N2940,N2941,N2942,N2948,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,
    N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
    N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,
    N3003,N3006,N3007,N3010,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
    N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3038,N3041,N3052,N3063,N3068,
    N3071,N3072,N3073,N3074,N3075,N3086,N3097,N3108,N3119,N3130,N3141,N3142,N3143,N3144,N3145,N3146,
    N3147,N3158,N3169,N3180,N3191,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3203,N3401,N3402,N3403,
    N3404,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3444,N3445,N3446,
    N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3459,N3460,N3461,N3462,N3463,N3464,
    N3465,N3466,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3502,
    N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3558,N3559,N3560,
    N3561,N3562,N3563,N3605,N3606,N3607,N3608,N3609,N3610,N3614,N3615,N3616,N3617,N3618,N3619,N3620,
    N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,
    N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,
    N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,
    N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,
    N3685,N3686,N3687,N3688,N3689,N3691,N3700,N3701,N3702,N3703,N3704,N3705,N3708,N3709,N3710,N3711,
    N3712,N3713,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,
    N3729,N3730,N3731,N3732,N3738,N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,
    N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,
    N3766,N3767,N3768,N3769,N3770,N3771,N3775,N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,
    N3788,N3789,N3793,N3797,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,N3813,
    N3816,N3819,N3822,N3823,N3824,N3827,N3828,N3829,N3830,N3831,N3834,N3835,N3836,N3837,N3838,N3839,
    N3840,N3841,N3842,N3849,N3855,N3861,N3867,N3873,N3881,N3887,N3893,N3908,N3909,N3911,N3914,N3915,
    N3916,N3917,N3918,N3919,N3920,N3921,N3927,N3933,N3942,N3948,N3956,N3962,N3968,N3975,N3976,N3977,
    N3978,N3979,N3980,N3981,N3982,N3983,N3984,N3987,N3988,N3989,N3990,N3991,N3998,N4008,N4011,N4021,
    N4024,N4027,N4031,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4067,N4080,
    N4088,N4091,N4094,N4097,N4100,N4103,N4106,N4109,N4144,N4147,N4150,N4153,N4156,N4159,N4183,N4184,
    N4185,N4186,N4188,N4191,N4196,N4197,N4198,N4199,N4200,N4203,N4206,N4209,N4212,N4215,N4219,N4223,
    N4224,N4225,N4228,N4231,N4234,N4237,N4240,N4243,N4246,N4249,N4252,N4255,N4258,N4263,N4264,N4267,
    N4268,N4269,N4270,N4271,N4273,N4274,N4276,N4277,N4280,N4284,N4290,N4297,N4298,N4301,N4305,N4310,
    N4316,N4320,N4325,N4331,N4332,N4336,N4342,N4349,N4357,N4364,N4375,N4379,N4385,N4392,N4396,N4400,
    N4405,N4412,N4418,N4425,N4436,N4440,N4445,N4451,N4456,N4462,N4469,N4477,N4512,N4515,N4516,N4521,
    N4523,N4524,N4532,N4547,N4548,N4551,N4554,N4557,N4560,N4563,N4566,N4569,N4572,N4575,N4578,N4581,
    N4584,N4587,N4590,N4593,N4596,N4599,N4602,N4605,N4608,N4611,N4614,N4617,N4621,N4624,N4627,N4630,
    N4633,N4637,N4640,N4643,N4646,N4649,N4652,N4655,N4658,N4662,N4665,N4668,N4671,N4674,N4677,N4680,
    N4683,N4686,N4689,N4692,N4695,N4698,N4701,N4702,N4720,N4721,N4724,N4725,N4726,N4727,N4728,N4729,
    N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4741,N4855,N4856,N4908,N4909,N4939,N4942,N4947,N4953,
    N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4965,N4966,N4967,N4968,N4972,N4973,N4974,N4975,
    N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N5049,N5052,N5053,N5054,
    N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5065,N5066,N5067,N5068,N5069,N5070,N5071,
    N5072,N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,
    N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,
    N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,N5118,N5119,
    N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5135,N5136,
    N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5150,N5153,N5154,N5155,
    N5156,N5157,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5169,N5172,N5173,N5176,N5177,N5180,N5183,
    N5186,N5189,N5192,N5195,N5198,N5199,N5202,N5205,N5208,N5211,N5214,N5217,N5220,N5223,N5224,N5225,
    N5226,N5227,N5228,N5229,N5230,N5232,N5233,N5234,N5235,N5236,N5239,N5241,N5242,N5243,N5244,N5245,
    N5246,N5247,N5248,N5249,N5250,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,
    N5263,N5264,N5274,N5275,N5282,N5283,N5284,N5298,N5299,N5300,N5303,N5304,N5305,N5306,N5307,N5308,
    N5309,N5310,N5311,N5312,N5315,N5319,N5324,N5328,N5331,N5332,N5346,N5363,N5364,N5365,N5366,N5367,
    N5368,N5369,N5370,N5371,N5374,N5377,N5382,N5385,N5389,N5396,N5407,N5418,N5424,N5431,N5441,N5452,
    N5462,N5469,N5470,N5477,N5488,N5498,N5506,N5520,N5536,N5549,N5555,N5562,N5573,N5579,N5595,N5606,
    N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5624,N5634,N5655,N5671,N5684,N5690,N5691,N5692,N5696,
    N5700,N5703,N5707,N5711,N5726,N5727,N5728,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5739,N5742,
    N5745,N5755,N5756,N5954,N5955,N5956,N6005,N6006,N6023,N6024,N6025,N6028,N6031,N6034,N6037,N6040,
    N6044,N6045,N6048,N6051,N6054,N6065,N6066,N6067,N6068,N6069,N6071,N6072,N6073,N6074,N6075,N6076,
    N6077,N6078,N6079,N6080,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,N6091,N6094,N6095,N6096,
    N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6111,N6112,N6113,N6114,
    N6115,N6116,N6117,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,
    N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6152,
    N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6168,N6171,N6172,N6173,
    N6174,N6175,N6178,N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,
    N6192,N6193,N6194,N6197,N6200,N6203,N6206,N6209,N6212,N6215,N6218,N6221,N6234,N6235,N6238,N6241,
    N6244,N6247,N6250,N6253,N6256,N6259,N6262,N6265,N6268,N6271,N6274,N6277,N6280,N6283,N6286,N6289,
    N6292,N6295,N6298,N6301,N6304,N6307,N6310,N6313,N6316,N6319,N6322,N6325,N6328,N6331,N6335,N6338,
    N6341,N6344,N6347,N6350,N6353,N6356,N6359,N6364,N6367,N6370,N6373,N6374,N6375,N6376,N6377,N6378,
    N6382,N6386,N6388,N6392,N6397,N6411,N6415,N6419,N6427,N6434,N6437,N6441,N6445,N6448,N6449,N6466,
    N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6478,N6482,N6486,N6490,N6494,N6500,N6504,
    N6508,N6512,N6516,N6526,N6536,N6539,N6553,N6556,N6566,N6569,N6572,N6575,N6580,N6584,N6587,N6592,
    N6599,N6606,N6609,N6619,N6622,N6630,N6631,N6632,N6633,N6634,N6637,N6640,N6650,N6651,N6653,N6655,
    N6657,N6659,N6660,N6661,N6662,N6663,N6664,N6666,N6668,N6670,N6672,N6675,N6680,N6681,N6682,N6683,
    N6689,N6690,N6691,N6692,N6693,N6695,N6698,N6699,N6700,N6703,N6708,N6709,N6710,N6711,N6712,N6713,
    N6714,N6715,N6718,N6719,N6720,N6721,N6722,N6724,N6739,N6740,N6741,N6744,N6745,N6746,N6751,N6752,
    N6753,N6754,N6755,N6760,N6761,N6762,N6772,N6773,N6776,N6777,N6782,N6783,N6784,N6785,N6790,N6791,
    N6792,N6795,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,N6811,N6812,N6813,N6814,
    N6815,N6816,N6817,N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6834,N6835,N6836,N6837,
    N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6860,
    N6861,N6862,N6863,N6866,N6872,N6873,N6874,N6875,N6876,N6879,N6880,N6881,N6884,N6885,N6888,N6889,
    N6890,N6891,N6894,N6895,N6896,N6897,N6900,N6901,N6904,N6905,N6908,N6909,N6912,N6913,N6914,N6915,
    N6916,N6919,N6922,N6923,N6930,N6932,N6935,N6936,N6937,N6938,N6939,N6940,N6946,N6947,N6948,N6949,
    N6953,N6954,N6955,N6956,N6957,N6958,N6964,N6965,N6966,N6967,N6973,N6974,N6975,N6976,N6977,N6978,
    N6979,N6987,N6990,N6999,N7002,N7003,N7006,N7011,N7012,N7013,N7016,N7018,N7019,N7020,N7021,N7022,
    N7023,N7028,N7031,N7034,N7037,N7040,N7041,N7044,N7045,N7046,N7047,N7048,N7049,N7054,N7057,N7060,
    N7064,N7065,N7072,N7073,N7074,N7075,N7076,N7079,N7080,N7083,N7084,N7085,N7086,N7087,N7088,N7089,
    N7090,N7093,N7094,N7097,N7101,N7105,N7110,N7114,N7115,N7116,N7125,N7126,N7127,N7130,N7131,N7139,
    N7140,N7141,N7146,N7147,N7149,N7150,N7151,N7152,N7153,N7158,N7159,N7160,N7166,N7167,N7168,N7169,
    N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,N7185,
    N7186,N7187,N7188,N7189,N7190,N7196,N7197,N7198,N7204,N7205,N7206,N7207,N7208,N7209,N7212,N7215,
    N7216,N7217,N7218,N7219,N7222,N7225,N7228,N7229,N7236,N7239,N7242,N7245,N7250,N7257,N7260,N7263,
    N7268,N7269,N7270,N7276,N7282,N7288,N7294,N7300,N7301,N7304,N7310,N7320,N7321,N7328,N7338,N7339,
    N7340,N7341,N7342,N7349,N7357,N7364,N7394,N7397,N7402,N7405,N7406,N7407,N7408,N7409,N7412,N7415,
    N7416,N7417,N7418,N7419,N7420,N7421,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7433,N7434,
    N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7450,N7451,
    N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,N7464,N7468,N7479,N7481,
    N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,N7492,N7493,N7498,N7499,N7500,N7505,N7507,N7508,
    N7509,N7510,N7512,N7513,N7514,N7525,N7526,N7527,N7528,N7529,N7530,N7531,N7537,N7543,N7549,N7555,
    N7561,N7567,N7573,N7579,N7582,N7585,N7586,N7587,N7588,N7589,N7592,N7595,N7598,N7599,N7624,N7625,
    N7631,N7636,N7657,N7658,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,
    N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,
    N7693,N7694,N7695,N7696,N7697,N7708,N7709,N7710,N7711,N7712,N7715,N7718,N7719,N7720,N7721,N7722,
    N7723,N7724,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7743,N7744,N7749,N7750,N7751,N7762,
    N7765,N7768,N7769,N7770,N7771,N7772,N7775,N7778,N7781,N7782,N7787,N7788,N7795,N7796,N7797,N7798,
    N7799,N7800,N7803,N7806,N7807,N7808,N7809,N7810,N7811,N7812,N7815,N7816,N7821,N7822,N7823,N7826,
    N7829,N7832,N7833,N7834,N7835,N7836,N7839,N7842,N7845,N7846,N7851,N7852,N7859,N7860,N7861,N7862,
    N7863,N7864,N7867,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7879,N7880,N7885,N7886,N7887,N7890,
    N7893,N7896,N7897,N7898,N7899,N7900,N7903,N7906,N7909,N7910,N7917,N7918,N7923,N7924,N7925,N7926,
    N7927,N7928,N7929,N7930,N7931,N7932,N7935,N7938,N7939,N7940,N7943,N7944,N7945,N7946,N7951,N7954,
    N7957,N7960,N7963,N7966,N7967,N7968,N7969,N7970,N7973,N7974,N7984,N7985,N7987,N7988,N7989,N7990,
    N7991,N7992,N7993,N7994,N7995,N7996,N7997,N7998,N8001,N8004,N8009,N8013,N8017,N8020,N8021,N8022,
    N8023,N8025,N8026,N8027,N8031,N8032,N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,
    N8043,N8044,N8045,N8048,N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8064,N8071,N8072,N8073,N8074,
    N8077,N8078,N8079,N8082,N8089,N8090,N8091,N8092,N8093,N8096,N8099,N8102,N8113,N8114,N8115,N8116,
    N8117,N8118,N8119,N8120,N8121,N8122,N8125,N8126,extra0,extra1,extra2,extra3,extra4,extra5,extra6,extra7,
    extra8,extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,extra17,extra18,extra19,extra20,extra21,extra22,extra23,
    extra24;

  BUF_X1 BUFF1_1( .Z(N709), .A(N141) );
  BUF_X1 BUFF1_2( .Z(N816), .A(N293) );
  AND2_X1 AND2_3( .ZN(N1042), .A1(N135), .A2(N631) );
  INV_X1 NOT1_4( .ZN(N1043), .A(N591) );
  BUF_X1 BUFF1_5( .Z(N1066), .A(N592) );
  INV_X1 NOT1_6( .ZN(N1067), .A(N595) );
  INV_X1 NOT1_7( .ZN(N1080), .A(N596) );
  INV_X1 NOT1_8( .ZN(N1092), .A(N597) );
  INV_X1 NOT1_9( .ZN(N1104), .A(N598) );
  INV_X1 NOT1_10( .ZN(N1137), .A(N545) );
  INV_X1 NOT1_11( .ZN(N1138), .A(N348) );
  INV_X1 NOT1_12( .ZN(N1139), .A(N366) );
  AND2_X1 AND2_13( .ZN(N1140), .A1(N552), .A2(N562) );
  INV_X1 NOT1_14( .ZN(N1141), .A(N549) );
  INV_X2 NOT1_15( .ZN(N1142), .A(N545) );
  INV_X1 NOT1_16( .ZN(N1143), .A(N545) );
  INV_X1 NOT1_17( .ZN(N1144), .A(N338) );
  INV_X1 NOT1_18( .ZN(N1145), .A(N358) );
  NAND2_X1 NAND2_19( .ZN(N1146), .A1(N373), .A2(N1) );
  AND2_X1 AND2_20( .ZN(N1147), .A1(N141), .A2(N145) );
  INV_X1 NOT1_21( .ZN(N1148), .A(N592) );
  INV_X1 NOT1_22( .ZN(N1149), .A(N1042) );
  AND2_X1 AND2_23( .ZN(N1150), .A1(N1043), .A2(N27) );
  AND2_X1 AND2_24( .ZN(N1151), .A1(N386), .A2(N556) );
  INV_X1 NOT1_25( .ZN(N1152), .A(N245) );
  INV_X1 NOT1_26( .ZN(N1153), .A(N552) );
  INV_X1 NOT1_27( .ZN(N1154), .A(N562) );
  INV_X1 NOT1_28( .ZN(N1155), .A(N559) );
  AND4_X1 AND4_29( .ZN(N1156), .A1(N386), .A2(N559), .A3(N556), .A4(N552) );
  INV_X1 NOT1_30( .ZN(N1157), .A(N566) );
  BUF_X1 BUFF1_31( .Z(N1161), .A(N571) );
  BUF_X1 BUFF1_32( .Z(N1173), .A(N574) );
  BUF_X1 BUFF1_33( .Z(N1185), .A(N571) );
  BUF_X2 BUFF1_34( .Z(N1197), .A(N574) );
  BUF_X1 BUFF1_35( .Z(N1209), .A(N137) );
  BUF_X1 BUFF1_36( .Z(N1213), .A(N137) );
  BUF_X1 BUFF1_37( .Z(N1216), .A(N141) );
  INV_X1 NOT1_38( .ZN(N1219), .A(N583) );
  BUF_X1 BUFF1_39( .Z(N1223), .A(N577) );
  BUF_X1 BUFF1_40( .Z(N1235), .A(N580) );
  BUF_X1 BUFF1_41( .Z(N1247), .A(N577) );
  BUF_X1 BUFF1_42( .Z(N1259), .A(N580) );
  BUF_X1 BUFF1_43( .Z(N1271), .A(N254) );
  BUF_X1 BUFF1_44( .Z(N1280), .A(N251) );
  BUF_X1 BUFF1_45( .Z(N1292), .A(N251) );
  BUF_X1 BUFF1_46( .Z(N1303), .A(N248) );
  BUF_X1 BUFF1_47( .Z(N1315), .A(N248) );
  BUF_X1 BUFF1_48( .Z(N1327), .A(N610) );
  BUF_X4 BUFF1_49( .Z(N1339), .A(N607) );
  BUF_X1 BUFF1_50( .Z(N1351), .A(N613) );
  BUF_X1 BUFF1_51( .Z(N1363), .A(N616) );
  BUF_X1 BUFF1_52( .Z(N1375), .A(N210) );
  BUF_X1 BUFF1_53( .Z(N1378), .A(N210) );
  BUF_X1 BUFF1_54( .Z(N1381), .A(N218) );
  BUF_X1 BUFF1_55( .Z(N1384), .A(N218) );
  BUF_X1 BUFF1_56( .Z(N1387), .A(N226) );
  BUF_X1 BUFF1_57( .Z(N1390), .A(N226) );
  BUF_X1 BUFF1_58( .Z(N1393), .A(N234) );
  BUF_X1 BUFF1_59( .Z(N1396), .A(N234) );
  BUF_X1 BUFF1_60( .Z(N1415), .A(N257) );
  BUF_X1 BUFF1_61( .Z(N1418), .A(N257) );
  BUF_X1 BUFF1_62( .Z(N1421), .A(N265) );
  BUF_X1 BUFF1_63( .Z(N1424), .A(N265) );
  BUF_X1 BUFF1_64( .Z(N1427), .A(N273) );
  BUF_X1 BUFF1_65( .Z(N1430), .A(N273) );
  BUF_X1 BUFF1_66( .Z(N1433), .A(N281) );
  BUF_X1 BUFF1_67( .Z(N1436), .A(N281) );
  BUF_X1 BUFF1_68( .Z(N1455), .A(N335) );
  BUF_X1 BUFF1_69( .Z(N1462), .A(N335) );
  BUF_X1 BUFF1_70( .Z(N1469), .A(N206) );
  AND2_X1 AND2_71( .ZN(N1475), .A1(N27), .A2(N31) );
  BUF_X1 BUFF1_72( .Z(N1479), .A(N1) );
  BUF_X4 BUFF1_73( .Z(N1482), .A(N588) );
  BUF_X1 BUFF1_74( .Z(N1492), .A(N293) );
  BUF_X1 BUFF1_75( .Z(N1495), .A(N302) );
  BUF_X1 BUFF1_76( .Z(N1498), .A(N308) );
  BUF_X1 BUFF1_77( .Z(N1501), .A(N308) );
  BUF_X1 BUFF1_78( .Z(N1504), .A(N316) );
  BUF_X1 BUFF1_79( .Z(N1507), .A(N316) );
  BUF_X1 BUFF1_80( .Z(N1510), .A(N324) );
  BUF_X1 BUFF1_81( .Z(N1513), .A(N324) );
  BUF_X1 BUFF1_82( .Z(N1516), .A(N341) );
  BUF_X4 BUFF1_83( .Z(N1519), .A(N341) );
  BUF_X1 BUFF1_84( .Z(N1522), .A(N351) );
  BUF_X8 BUFF1_85( .Z(N1525), .A(N351) );
  BUF_X1 BUFF1_86( .Z(N1542), .A(N257) );
  BUF_X1 BUFF1_87( .Z(N1545), .A(N257) );
  BUF_X1 BUFF1_88( .Z(N1548), .A(N265) );
  BUF_X1 BUFF1_89( .Z(N1551), .A(N265) );
  BUF_X1 BUFF1_90( .Z(N1554), .A(N273) );
  BUF_X1 BUFF1_91( .Z(N1557), .A(N273) );
  BUF_X1 BUFF1_92( .Z(N1560), .A(N281) );
  BUF_X1 BUFF1_93( .Z(N1563), .A(N281) );
  BUF_X1 BUFF1_94( .Z(N1566), .A(N332) );
  BUF_X1 BUFF1_95( .Z(N1573), .A(N332) );
  BUF_X1 BUFF1_96( .Z(N1580), .A(N549) );
  AND2_X1 AND2_97( .ZN(N1583), .A1(N31), .A2(N27) );
  INV_X1 NOT1_98( .ZN(N1588), .A(N588) );
  BUF_X1 BUFF1_99( .Z(N1594), .A(N324) );
  BUF_X1 BUFF1_100( .Z(N1597), .A(N324) );
  BUF_X1 BUFF1_101( .Z(N1600), .A(N341) );
  BUF_X1 BUFF1_102( .Z(N1603), .A(N341) );
  BUF_X8 BUFF1_103( .Z(N1606), .A(N351) );
  BUF_X1 BUFF1_104( .Z(N1609), .A(N351) );
  BUF_X1 BUFF1_105( .Z(N1612), .A(N293) );
  BUF_X1 BUFF1_106( .Z(N1615), .A(N302) );
  BUF_X1 BUFF1_107( .Z(N1618), .A(N308) );
  BUF_X1 BUFF1_108( .Z(N1621), .A(N308) );
  BUF_X8 BUFF1_109( .Z(N1624), .A(N316) );
  BUF_X1 BUFF1_110( .Z(N1627), .A(N316) );
  BUF_X1 BUFF1_111( .Z(N1630), .A(N361) );
  BUF_X1 BUFF1_112( .Z(N1633), .A(N361) );
  BUF_X1 BUFF1_113( .Z(N1636), .A(N210) );
  BUF_X1 BUFF1_114( .Z(N1639), .A(N210) );
  BUF_X1 BUFF1_115( .Z(N1642), .A(N218) );
  BUF_X1 BUFF1_116( .Z(N1645), .A(N218) );
  BUF_X1 BUFF1_117( .Z(N1648), .A(N226) );
  BUF_X1 BUFF1_118( .Z(N1651), .A(N226) );
  BUF_X1 BUFF1_119( .Z(N1654), .A(N234) );
  BUF_X1 BUFF1_120( .Z(N1657), .A(N234) );
  INV_X1 NOT1_121( .ZN(N1660), .A(N324) );
  BUF_X1 BUFF1_122( .Z(N1663), .A(N242) );
  BUF_X1 BUFF1_123( .Z(N1675), .A(N242) );
  BUF_X1 BUFF1_124( .Z(N1685), .A(N254) );
  BUF_X1 BUFF1_125( .Z(N1697), .A(N610) );
  BUF_X1 BUFF1_126( .Z(N1709), .A(N607) );
  BUF_X1 BUFF1_127( .Z(N1721), .A(N625) );
  BUF_X1 BUFF1_128( .Z(N1727), .A(N619) );
  BUF_X1 BUFF1_129( .Z(N1731), .A(N613) );
  BUF_X1 BUFF1_130( .Z(N1743), .A(N616) );
  INV_X1 NOT1_131( .ZN(N1755), .A(N599) );
  INV_X1 NOT1_132( .ZN(N1758), .A(N603) );
  BUF_X1 BUFF1_133( .Z(N1761), .A(N619) );
  BUF_X1 BUFF1_134( .Z(N1769), .A(N625) );
  BUF_X1 BUFF1_135( .Z(N1777), .A(N619) );
  BUF_X1 BUFF1_136( .Z(N1785), .A(N625) );
  BUF_X1 BUFF1_137( .Z(N1793), .A(N619) );
  BUF_X1 BUFF1_138( .Z(N1800), .A(N625) );
  BUF_X1 BUFF1_139( .Z(N1807), .A(N619) );
  BUF_X8 BUFF1_140( .Z(N1814), .A(N625) );
  BUF_X1 BUFF1_141( .Z(N1821), .A(N299) );
  BUF_X1 BUFF1_142( .Z(N1824), .A(N446) );
  BUF_X1 BUFF1_143( .Z(N1827), .A(N457) );
  BUF_X1 BUFF1_144( .Z(N1830), .A(N468) );
  BUF_X1 BUFF1_145( .Z(N1833), .A(N422) );
  BUF_X1 BUFF1_146( .Z(N1836), .A(N435) );
  BUF_X1 BUFF1_147( .Z(N1839), .A(N389) );
  BUF_X1 BUFF1_148( .Z(N1842), .A(N400) );
  BUF_X1 BUFF1_149( .Z(N1845), .A(N411) );
  BUF_X1 BUFF1_150( .Z(N1848), .A(N374) );
  BUF_X1 BUFF1_151( .Z(N1851), .A(N4) );
  BUF_X1 BUFF1_152( .Z(N1854), .A(N446) );
  BUF_X1 BUFF1_153( .Z(N1857), .A(N457) );
  BUF_X1 BUFF1_154( .Z(N1860), .A(N468) );
  BUF_X1 BUFF1_155( .Z(N1863), .A(N435) );
  BUF_X1 BUFF1_156( .Z(N1866), .A(N389) );
  BUF_X1 BUFF1_157( .Z(N1869), .A(N400) );
  BUF_X1 BUFF1_158( .Z(N1872), .A(N411) );
  BUF_X1 BUFF1_159( .Z(N1875), .A(N422) );
  BUF_X1 BUFF1_160( .Z(N1878), .A(N374) );
  BUF_X1 BUFF1_161( .Z(N1881), .A(N479) );
  BUF_X1 BUFF1_162( .Z(N1884), .A(N490) );
  BUF_X1 BUFF1_163( .Z(N1887), .A(N503) );
  BUF_X1 BUFF1_164( .Z(N1890), .A(N514) );
  BUF_X1 BUFF1_165( .Z(N1893), .A(N523) );
  BUF_X1 BUFF1_166( .Z(N1896), .A(N534) );
  BUF_X1 BUFF1_167( .Z(N1899), .A(N54) );
  BUF_X1 BUFF1_168( .Z(N1902), .A(N479) );
  BUF_X1 BUFF1_169( .Z(N1905), .A(N503) );
  BUF_X1 BUFF1_170( .Z(N1908), .A(N514) );
  BUF_X1 BUFF1_171( .Z(N1911), .A(N523) );
  BUF_X4 BUFF1_172( .Z(N1914), .A(N534) );
  BUF_X1 BUFF1_173( .Z(N1917), .A(N490) );
  BUF_X1 BUFF1_174( .Z(N1920), .A(N361) );
  BUF_X1 BUFF1_175( .Z(N1923), .A(N369) );
  BUF_X1 BUFF1_176( .Z(N1926), .A(N341) );
  BUF_X1 BUFF1_177( .Z(N1929), .A(N351) );
  BUF_X1 BUFF1_178( .Z(N1932), .A(N308) );
  BUF_X1 BUFF1_179( .Z(N1935), .A(N316) );
  BUF_X1 BUFF1_180( .Z(N1938), .A(N293) );
  BUF_X1 BUFF1_181( .Z(N1941), .A(N302) );
  BUF_X1 BUFF1_182( .Z(N1944), .A(N281) );
  BUF_X1 BUFF1_183( .Z(N1947), .A(N289) );
  BUF_X1 BUFF1_184( .Z(N1950), .A(N265) );
  BUF_X1 BUFF1_185( .Z(N1953), .A(N273) );
  BUF_X1 BUFF1_186( .Z(N1956), .A(N234) );
  BUF_X1 BUFF1_187( .Z(N1959), .A(N257) );
  BUF_X1 BUFF1_188( .Z(N1962), .A(N218) );
  BUF_X1 BUFF1_189( .Z(N1965), .A(N226) );
  BUF_X1 BUFF1_190( .Z(N1968), .A(N210) );
  INV_X1 NOT1_191( .ZN(N1972), .A(N1146) );
  AND2_X1 AND2_192( .ZN(N2054), .A1(N136), .A2(N1148) );
  INV_X1 NOT1_193( .ZN(N2060), .A(N1150) );
  INV_X1 NOT1_194( .ZN(N2061), .A(N1151) );
  BUF_X1 BUFF1_195( .Z(N2139), .A(N1209) );
  BUF_X1 BUFF1_196( .Z(N2142), .A(N1216) );
  BUF_X1 BUFF1_197( .Z(N2309), .A(N1479) );
  AND2_X1 AND2_198( .ZN(N2349), .A1(N1104), .A2(N514) );
  OR2_X1 OR2_199( .ZN(N2350), .A1(N1067), .A2(N514) );
  BUF_X1 BUFF1_200( .Z(N2387), .A(N1580) );
  BUF_X1 BUFF1_201( .Z(N2527), .A(N1821) );
  INV_X1 NOT1_202( .ZN(N2584), .A(N1580) );
  AND3_X1 AND3_203( .ZN(N2585), .A1(N170), .A2(N1161), .A3(N1173) );
  AND3_X1 AND3_204( .ZN(N2586), .A1(N173), .A2(N1161), .A3(N1173) );
  AND3_X1 AND3_205( .ZN(N2587), .A1(N167), .A2(N1161), .A3(N1173) );
  AND3_X1 AND3_206( .ZN(N2588), .A1(N164), .A2(N1161), .A3(N1173) );
  AND3_X1 AND3_207( .ZN(N2589), .A1(N161), .A2(N1161), .A3(N1173) );
  NAND2_X1 NAND2_208( .ZN(N2590), .A1(N1475), .A2(N140) );
  AND3_X1 AND3_209( .ZN(N2591), .A1(N185), .A2(N1185), .A3(N1197) );
  AND3_X1 AND3_210( .ZN(N2592), .A1(N158), .A2(N1185), .A3(N1197) );
  AND3_X2 AND3_211( .ZN(N2593), .A1(N152), .A2(N1185), .A3(N1197) );
  AND3_X2 AND3_212( .ZN(N2594), .A1(N146), .A2(N1185), .A3(N1197) );
  AND3_X2 AND3_213( .ZN(N2595), .A1(N170), .A2(N1223), .A3(N1235) );
  AND3_X1 AND3_214( .ZN(N2596), .A1(N173), .A2(N1223), .A3(N1235) );
  AND3_X1 AND3_215( .ZN(N2597), .A1(N167), .A2(N1223), .A3(N1235) );
  AND3_X1 AND3_216( .ZN(N2598), .A1(N164), .A2(N1223), .A3(N1235) );
  AND3_X1 AND3_217( .ZN(N2599), .A1(N161), .A2(N1223), .A3(N1235) );
  AND3_X1 AND3_218( .ZN(N2600), .A1(N185), .A2(N1247), .A3(N1259) );
  AND3_X1 AND3_219( .ZN(N2601), .A1(N158), .A2(N1247), .A3(N1259) );
  AND3_X1 AND3_220( .ZN(N2602), .A1(N152), .A2(N1247), .A3(N1259) );
  AND3_X1 AND3_221( .ZN(N2603), .A1(N146), .A2(N1247), .A3(N1259) );
  AND3_X1 AND3_222( .ZN(N2604), .A1(N106), .A2(N1731), .A3(N1743) );
  AND3_X1 AND3_223( .ZN(N2605), .A1(N61), .A2(N1327), .A3(N1339) );
  AND3_X1 AND3_224( .ZN(N2606), .A1(N106), .A2(N1697), .A3(N1709) );
  AND3_X1 AND3_225( .ZN(N2607), .A1(N49), .A2(N1697), .A3(N1709) );
  AND3_X1 AND3_226( .ZN(N2608), .A1(N103), .A2(N1697), .A3(N1709) );
  AND3_X1 AND3_227( .ZN(N2609), .A1(N40), .A2(N1697), .A3(N1709) );
  AND3_X1 AND3_228( .ZN(N2610), .A1(N37), .A2(N1697), .A3(N1709) );
  AND3_X1 AND3_229( .ZN(N2611), .A1(N20), .A2(N1327), .A3(N1339) );
  AND3_X1 AND3_230( .ZN(N2612), .A1(N17), .A2(N1327), .A3(N1339) );
  AND3_X1 AND3_231( .ZN(N2613), .A1(N70), .A2(N1327), .A3(N1339) );
  AND3_X1 AND3_232( .ZN(N2614), .A1(N64), .A2(N1327), .A3(N1339) );
  AND3_X1 AND3_233( .ZN(N2615), .A1(N49), .A2(N1731), .A3(N1743) );
  AND3_X1 AND3_234( .ZN(N2616), .A1(N103), .A2(N1731), .A3(N1743) );
  AND3_X1 AND3_235( .ZN(N2617), .A1(N40), .A2(N1731), .A3(N1743) );
  AND3_X1 AND3_236( .ZN(N2618), .A1(N37), .A2(N1731), .A3(N1743) );
  AND3_X1 AND3_237( .ZN(N2619), .A1(N20), .A2(N1351), .A3(N1363) );
  AND3_X1 AND3_238( .ZN(N2620), .A1(N17), .A2(N1351), .A3(N1363) );
  AND3_X1 AND3_239( .ZN(N2621), .A1(N70), .A2(N1351), .A3(N1363) );
  AND3_X1 AND3_240( .ZN(N2622), .A1(N64), .A2(N1351), .A3(N1363) );
  INV_X1 NOT1_241( .ZN(N2623), .A(N1475) );
  AND3_X1 AND3_242( .ZN(N2624), .A1(N123), .A2(N1758), .A3(N599) );
  AND2_X1 AND2_243( .ZN(N2625), .A1(N1777), .A2(N1785) );
  AND3_X1 AND3_244( .ZN(N2626), .A1(N61), .A2(N1351), .A3(N1363) );
  AND2_X1 AND2_245( .ZN(N2627), .A1(N1761), .A2(N1769) );
  INV_X1 NOT1_246( .ZN(N2628), .A(N1824) );
  INV_X1 NOT1_247( .ZN(N2629), .A(N1827) );
  INV_X1 NOT1_248( .ZN(N2630), .A(N1830) );
  INV_X1 NOT1_249( .ZN(N2631), .A(N1833) );
  INV_X1 NOT1_250( .ZN(N2632), .A(N1836) );
  INV_X1 NOT1_251( .ZN(N2633), .A(N1839) );
  INV_X2 NOT1_252( .ZN(N2634), .A(N1842) );
  INV_X2 NOT1_253( .ZN(N2635), .A(N1845) );
  INV_X1 NOT1_254( .ZN(N2636), .A(N1848) );
  INV_X1 NOT1_255( .ZN(N2637), .A(N1851) );
  INV_X1 NOT1_256( .ZN(N2638), .A(N1854) );
  INV_X1 NOT1_257( .ZN(N2639), .A(N1857) );
  INV_X1 NOT1_258( .ZN(N2640), .A(N1860) );
  INV_X1 NOT1_259( .ZN(N2641), .A(N1863) );
  INV_X1 NOT1_260( .ZN(N2642), .A(N1866) );
  INV_X1 NOT1_261( .ZN(N2643), .A(N1869) );
  INV_X1 NOT1_262( .ZN(N2644), .A(N1872) );
  INV_X1 NOT1_263( .ZN(N2645), .A(N1875) );
  INV_X1 NOT1_264( .ZN(N2646), .A(N1878) );
  BUF_X1 BUFF1_265( .Z(N2647), .A(N1209) );
  INV_X1 NOT1_266( .ZN(N2653), .A(N1161) );
  INV_X1 NOT1_267( .ZN(N2664), .A(N1173) );
  BUF_X1 BUFF1_268( .Z(N2675), .A(N1209) );
  INV_X1 NOT1_269( .ZN(N2681), .A(N1185) );
  INV_X1 NOT1_270( .ZN(N2692), .A(N1197) );
  AND3_X1 AND3_271( .ZN(N2703), .A1(N179), .A2(N1185), .A3(N1197) );
  BUF_X1 BUFF1_272( .Z(N2704), .A(N1479) );
  INV_X1 NOT1_273( .ZN(N2709), .A(N1881) );
  INV_X1 NOT1_274( .ZN(N2710), .A(N1884) );
  INV_X1 NOT1_275( .ZN(N2711), .A(N1887) );
  INV_X1 NOT1_276( .ZN(N2712), .A(N1890) );
  INV_X1 NOT1_277( .ZN(N2713), .A(N1893) );
  INV_X1 NOT1_278( .ZN(N2714), .A(N1896) );
  INV_X1 NOT1_279( .ZN(N2715), .A(N1899) );
  INV_X1 NOT1_280( .ZN(N2716), .A(N1902) );
  INV_X1 NOT1_281( .ZN(N2717), .A(N1905) );
  INV_X1 NOT1_282( .ZN(N2718), .A(N1908) );
  INV_X1 NOT1_283( .ZN(N2719), .A(N1911) );
  INV_X1 NOT1_284( .ZN(N2720), .A(N1914) );
  INV_X1 NOT1_285( .ZN(N2721), .A(N1917) );
  BUF_X1 BUFF1_286( .Z(N2722), .A(N1213) );
  INV_X1 NOT1_287( .ZN(N2728), .A(N1223) );
  INV_X1 NOT1_288( .ZN(N2739), .A(N1235) );
  BUF_X1 BUFF1_289( .Z(N2750), .A(N1213) );
  INV_X1 NOT1_290( .ZN(N2756), .A(N1247) );
  INV_X1 NOT1_291( .ZN(N2767), .A(N1259) );
  AND3_X1 AND3_292( .ZN(N2778), .A1(N179), .A2(N1247), .A3(N1259) );
  INV_X1 NOT1_293( .ZN(N2779), .A(N1327) );
  INV_X1 NOT1_294( .ZN(N2790), .A(N1339) );
  INV_X1 NOT1_295( .ZN(N2801), .A(N1351) );
  INV_X1 NOT1_296( .ZN(N2812), .A(N1363) );
  INV_X1 NOT1_297( .ZN(N2823), .A(N1375) );
  INV_X1 NOT1_298( .ZN(N2824), .A(N1378) );
  INV_X1 NOT1_299( .ZN(N2825), .A(N1381) );
  INV_X1 NOT1_300( .ZN(N2826), .A(N1384) );
  INV_X1 NOT1_301( .ZN(N2827), .A(N1387) );
  INV_X1 NOT1_302( .ZN(N2828), .A(N1390) );
  INV_X1 NOT1_303( .ZN(N2829), .A(N1393) );
  INV_X1 NOT1_304( .ZN(N2830), .A(N1396) );
  AND3_X1 AND3_305( .ZN(N2831), .A1(N1104), .A2(N457), .A3(N1378) );
  AND3_X2 AND3_306( .ZN(N2832), .A1(N1104), .A2(N468), .A3(N1384) );
  AND3_X2 AND3_307( .ZN(N2833), .A1(N1104), .A2(N422), .A3(N1390) );
  AND3_X1 AND3_308( .ZN(N2834), .A1(N1104), .A2(N435), .A3(N1396) );
  AND2_X1 AND2_309( .ZN(N2835), .A1(N1067), .A2(N1375) );
  AND2_X1 AND2_310( .ZN(N2836), .A1(N1067), .A2(N1381) );
  AND2_X1 AND2_311( .ZN(N2837), .A1(N1067), .A2(N1387) );
  AND2_X1 AND2_312( .ZN(N2838), .A1(N1067), .A2(N1393) );
  INV_X1 NOT1_313( .ZN(N2839), .A(N1415) );
  INV_X1 NOT1_314( .ZN(N2840), .A(N1418) );
  INV_X1 NOT1_315( .ZN(N2841), .A(N1421) );
  INV_X1 NOT1_316( .ZN(N2842), .A(N1424) );
  INV_X1 NOT1_317( .ZN(N2843), .A(N1427) );
  INV_X1 NOT1_318( .ZN(N2844), .A(N1430) );
  INV_X1 NOT1_319( .ZN(N2845), .A(N1433) );
  INV_X1 NOT1_320( .ZN(N2846), .A(N1436) );
  AND3_X1 AND3_321( .ZN(N2847), .A1(N1104), .A2(N389), .A3(N1418) );
  AND3_X1 AND3_322( .ZN(N2848), .A1(N1104), .A2(N400), .A3(N1424) );
  AND3_X1 AND3_323( .ZN(N2849), .A1(N1104), .A2(N411), .A3(N1430) );
  AND3_X1 AND3_324( .ZN(N2850), .A1(N1104), .A2(N374), .A3(N1436) );
  AND2_X1 AND2_325( .ZN(N2851), .A1(N1067), .A2(N1415) );
  AND2_X1 AND2_326( .ZN(N2852), .A1(N1067), .A2(N1421) );
  AND2_X1 AND2_327( .ZN(N2853), .A1(N1067), .A2(N1427) );
  AND2_X1 AND2_328( .ZN(N2854), .A1(N1067), .A2(N1433) );
  INV_X1 NOT1_329( .ZN(N2855), .A(N1455) );
  INV_X1 NOT1_330( .ZN(N2861), .A(N1462) );
  AND2_X1 AND2_331( .ZN(N2867), .A1(N292), .A2(N1455) );
  AND2_X1 AND2_332( .ZN(N2868), .A1(N288), .A2(N1455) );
  AND2_X1 AND2_333( .ZN(N2869), .A1(N280), .A2(N1455) );
  AND2_X1 AND2_334( .ZN(N2870), .A1(N272), .A2(N1455) );
  AND2_X1 AND2_335( .ZN(N2871), .A1(N264), .A2(N1455) );
  AND2_X4 AND2_336( .ZN(N2872), .A1(N241), .A2(N1462) );
  AND2_X1 AND2_337( .ZN(N2873), .A1(N233), .A2(N1462) );
  AND2_X1 AND2_338( .ZN(N2874), .A1(N225), .A2(N1462) );
  AND2_X1 AND2_339( .ZN(N2875), .A1(N217), .A2(N1462) );
  AND2_X1 AND2_340( .ZN(N2876), .A1(N209), .A2(N1462) );
  BUF_X1 BUFF1_341( .Z(N2877), .A(N1216) );
  INV_X1 NOT1_342( .ZN(N2882), .A(N1482) );
  INV_X1 NOT1_343( .ZN(N2891), .A(N1475) );
  INV_X1 NOT1_344( .ZN(N2901), .A(N1492) );
  INV_X1 NOT1_345( .ZN(N2902), .A(N1495) );
  INV_X1 NOT1_346( .ZN(N2903), .A(N1498) );
  INV_X1 NOT1_347( .ZN(N2904), .A(N1501) );
  INV_X1 NOT1_348( .ZN(N2905), .A(N1504) );
  INV_X1 NOT1_349( .ZN(N2906), .A(N1507) );
  AND2_X1 AND2_350( .ZN(N2907), .A1(N1303), .A2(N1495) );
  AND3_X1 AND3_351( .ZN(N2908), .A1(N1303), .A2(N479), .A3(N1501) );
  AND3_X1 AND3_352( .ZN(N2909), .A1(N1303), .A2(N490), .A3(N1507) );
  AND2_X1 AND2_353( .ZN(N2910), .A1(N1663), .A2(N1492) );
  AND2_X1 AND2_354( .ZN(N2911), .A1(N1663), .A2(N1498) );
  AND2_X1 AND2_355( .ZN(N2912), .A1(N1663), .A2(N1504) );
  INV_X1 NOT1_356( .ZN(N2913), .A(N1510) );
  INV_X8 NOT1_357( .ZN(N2914), .A(N1513) );
  INV_X1 NOT1_358( .ZN(N2915), .A(N1516) );
  INV_X1 NOT1_359( .ZN(N2916), .A(N1519) );
  INV_X1 NOT1_360( .ZN(N2917), .A(N1522) );
  INV_X1 NOT1_361( .ZN(N2918), .A(N1525) );
  AND3_X1 AND3_362( .ZN(N2919), .A1(N1104), .A2(N503), .A3(N1513) );
  INV_X1 NOT1_363( .ZN(N2920), .A(N2349) );
  AND3_X1 AND3_364( .ZN(N2921), .A1(N1104), .A2(N523), .A3(N1519) );
  AND3_X1 AND3_365( .ZN(N2922), .A1(N1104), .A2(N534), .A3(N1525) );
  AND2_X1 AND2_366( .ZN(N2923), .A1(N1067), .A2(N1510) );
  AND2_X1 AND2_367( .ZN(N2924), .A1(N1067), .A2(N1516) );
  AND2_X1 AND2_368( .ZN(N2925), .A1(N1067), .A2(N1522) );
  INV_X1 NOT1_369( .ZN(N2926), .A(N1542) );
  INV_X4 NOT1_370( .ZN(N2927), .A(N1545) );
  INV_X1 NOT1_371( .ZN(N2928), .A(N1548) );
  INV_X1 NOT1_372( .ZN(N2929), .A(N1551) );
  INV_X1 NOT1_373( .ZN(N2930), .A(N1554) );
  INV_X1 NOT1_374( .ZN(N2931), .A(N1557) );
  INV_X1 NOT1_375( .ZN(N2932), .A(N1560) );
  INV_X1 NOT1_376( .ZN(N2933), .A(N1563) );
  AND3_X1 AND3_377( .ZN(N2934), .A1(N1303), .A2(N389), .A3(N1545) );
  AND3_X1 AND3_378( .ZN(N2935), .A1(N1303), .A2(N400), .A3(N1551) );
  AND3_X1 AND3_379( .ZN(N2936), .A1(N1303), .A2(N411), .A3(N1557) );
  AND3_X1 AND3_380( .ZN(N2937), .A1(N1303), .A2(N374), .A3(N1563) );
  AND2_X1 AND2_381( .ZN(N2938), .A1(N1663), .A2(N1542) );
  AND2_X2 AND2_382( .ZN(N2939), .A1(N1663), .A2(N1548) );
  AND2_X1 AND2_383( .ZN(N2940), .A1(N1663), .A2(N1554) );
  AND2_X1 AND2_384( .ZN(N2941), .A1(N1663), .A2(N1560) );
  INV_X1 NOT1_385( .ZN(N2942), .A(N1566) );
  INV_X1 NOT1_386( .ZN(N2948), .A(N1573) );
  AND2_X1 AND2_387( .ZN(N2954), .A1(N372), .A2(N1566) );
  AND2_X1 AND2_388( .ZN(N2955), .A1(N366), .A2(N1566) );
  AND2_X1 AND2_389( .ZN(N2956), .A1(N358), .A2(N1566) );
  AND2_X1 AND2_390( .ZN(N2957), .A1(N348), .A2(N1566) );
  AND2_X1 AND2_391( .ZN(N2958), .A1(N338), .A2(N1566) );
  AND2_X1 AND2_392( .ZN(N2959), .A1(N331), .A2(N1573) );
  AND2_X1 AND2_393( .ZN(N2960), .A1(N323), .A2(N1573) );
  AND2_X1 AND2_394( .ZN(N2961), .A1(N315), .A2(N1573) );
  AND2_X1 AND2_395( .ZN(N2962), .A1(N307), .A2(N1573) );
  AND2_X1 AND2_396( .ZN(N2963), .A1(N299), .A2(N1573) );
  INV_X1 NOT1_397( .ZN(N2964), .A(N1588) );
  AND2_X1 AND2_398( .ZN(N2969), .A1(N83), .A2(N1588) );
  AND2_X1 AND2_399( .ZN(N2970), .A1(N86), .A2(N1588) );
  AND2_X1 AND2_400( .ZN(N2971), .A1(N88), .A2(N1588) );
  AND2_X1 AND2_401( .ZN(N2972), .A1(N88), .A2(N1588) );
  INV_X1 NOT1_402( .ZN(N2973), .A(N1594) );
  INV_X1 NOT1_403( .ZN(N2974), .A(N1597) );
  INV_X1 NOT1_404( .ZN(N2975), .A(N1600) );
  INV_X1 NOT1_405( .ZN(N2976), .A(N1603) );
  INV_X1 NOT1_406( .ZN(N2977), .A(N1606) );
  INV_X1 NOT1_407( .ZN(N2978), .A(N1609) );
  AND3_X1 AND3_408( .ZN(N2979), .A1(N1315), .A2(N503), .A3(N1597) );
  AND2_X1 AND2_409( .ZN(N2980), .A1(N1315), .A2(N514) );
  AND3_X1 AND3_410( .ZN(N2981), .A1(N1315), .A2(N523), .A3(N1603) );
  AND3_X1 AND3_411( .ZN(N2982), .A1(N1315), .A2(N534), .A3(N1609) );
  AND2_X1 AND2_412( .ZN(N2983), .A1(N1675), .A2(N1594) );
  OR2_X1 OR2_413( .ZN(N2984), .A1(N1675), .A2(N514) );
  AND2_X1 AND2_414( .ZN(N2985), .A1(N1675), .A2(N1600) );
  AND2_X1 AND2_415( .ZN(N2986), .A1(N1675), .A2(N1606) );
  INV_X1 NOT1_416( .ZN(N2987), .A(N1612) );
  INV_X1 NOT1_417( .ZN(N2988), .A(N1615) );
  INV_X1 NOT1_418( .ZN(N2989), .A(N1618) );
  INV_X1 NOT1_419( .ZN(N2990), .A(N1621) );
  INV_X1 NOT1_420( .ZN(N2991), .A(N1624) );
  INV_X1 NOT1_421( .ZN(N2992), .A(N1627) );
  AND2_X1 AND2_422( .ZN(N2993), .A1(N1315), .A2(N1615) );
  AND3_X2 AND3_423( .ZN(N2994), .A1(N1315), .A2(N479), .A3(N1621) );
  AND3_X1 AND3_424( .ZN(N2995), .A1(N1315), .A2(N490), .A3(N1627) );
  AND2_X1 AND2_425( .ZN(N2996), .A1(N1675), .A2(N1612) );
  AND2_X1 AND2_426( .ZN(N2997), .A1(N1675), .A2(N1618) );
  AND2_X1 AND2_427( .ZN(N2998), .A1(N1675), .A2(N1624) );
  INV_X1 NOT1_428( .ZN(N2999), .A(N1630) );
  BUF_X1 BUFF1_429( .Z(N3000), .A(N1469) );
  BUF_X1 BUFF1_430( .Z(N3003), .A(N1469) );
  INV_X1 NOT1_431( .ZN(N3006), .A(N1633) );
  BUF_X1 BUFF1_432( .Z(N3007), .A(N1469) );
  BUF_X1 BUFF1_433( .Z(N3010), .A(N1469) );
  AND2_X1 AND2_434( .ZN(N3013), .A1(N1315), .A2(N1630) );
  AND2_X1 AND2_435( .ZN(N3014), .A1(N1315), .A2(N1633) );
  INV_X1 NOT1_436( .ZN(N3015), .A(N1636) );
  INV_X1 NOT1_437( .ZN(N3016), .A(N1639) );
  INV_X1 NOT1_438( .ZN(N3017), .A(N1642) );
  INV_X1 NOT1_439( .ZN(N3018), .A(N1645) );
  INV_X1 NOT1_440( .ZN(N3019), .A(N1648) );
  INV_X1 NOT1_441( .ZN(N3020), .A(N1651) );
  INV_X1 NOT1_442( .ZN(N3021), .A(N1654) );
  INV_X1 NOT1_443( .ZN(N3022), .A(N1657) );
  AND3_X2 AND3_444( .ZN(N3023), .A1(N1303), .A2(N457), .A3(N1639) );
  AND3_X2 AND3_445( .ZN(N3024), .A1(N1303), .A2(N468), .A3(N1645) );
  AND3_X1 AND3_446( .ZN(N3025), .A1(N1303), .A2(N422), .A3(N1651) );
  AND3_X1 AND3_447( .ZN(N3026), .A1(N1303), .A2(N435), .A3(N1657) );
  AND2_X1 AND2_448( .ZN(N3027), .A1(N1663), .A2(N1636) );
  AND2_X1 AND2_449( .ZN(N3028), .A1(N1663), .A2(N1642) );
  AND2_X1 AND2_450( .ZN(N3029), .A1(N1663), .A2(N1648) );
  AND2_X1 AND2_451( .ZN(N3030), .A1(N1663), .A2(N1654) );
  INV_X1 NOT1_452( .ZN(N3031), .A(N1920) );
  INV_X1 NOT1_453( .ZN(N3032), .A(N1923) );
  INV_X1 NOT1_454( .ZN(N3033), .A(N1926) );
  INV_X1 NOT1_455( .ZN(N3034), .A(N1929) );
  BUF_X1 BUFF1_456( .Z(N3035), .A(N1660) );
  BUF_X1 BUFF1_457( .Z(N3038), .A(N1660) );
  INV_X1 NOT1_458( .ZN(N3041), .A(N1697) );
  INV_X1 NOT1_459( .ZN(N3052), .A(N1709) );
  INV_X1 NOT1_460( .ZN(N3063), .A(N1721) );
  INV_X1 NOT1_461( .ZN(N3068), .A(N1727) );
  AND2_X1 AND2_462( .ZN(N3071), .A1(N97), .A2(N1721) );
  AND2_X1 AND2_463( .ZN(N3072), .A1(N94), .A2(N1721) );
  AND2_X1 AND2_464( .ZN(N3073), .A1(N97), .A2(N1721) );
  AND2_X1 AND2_465( .ZN(N3074), .A1(N94), .A2(N1721) );
  INV_X1 NOT1_466( .ZN(N3075), .A(N1731) );
  INV_X1 NOT1_467( .ZN(N3086), .A(N1743) );
  INV_X1 NOT1_468( .ZN(N3097), .A(N1761) );
  INV_X1 NOT1_469( .ZN(N3108), .A(N1769) );
  INV_X1 NOT1_470( .ZN(N3119), .A(N1777) );
  INV_X1 NOT1_471( .ZN(N3130), .A(N1785) );
  INV_X1 NOT1_472( .ZN(N3141), .A(N1944) );
  INV_X1 NOT1_473( .ZN(N3142), .A(N1947) );
  INV_X1 NOT1_474( .ZN(N3143), .A(N1950) );
  INV_X1 NOT1_475( .ZN(N3144), .A(N1953) );
  INV_X1 NOT1_476( .ZN(N3145), .A(N1956) );
  INV_X1 NOT1_477( .ZN(N3146), .A(N1959) );
  INV_X1 NOT1_478( .ZN(N3147), .A(N1793) );
  INV_X1 NOT1_479( .ZN(N3158), .A(N1800) );
  INV_X1 NOT1_480( .ZN(N3169), .A(N1807) );
  INV_X1 NOT1_481( .ZN(N3180), .A(N1814) );
  BUF_X1 BUFF1_482( .Z(N3191), .A(N1821) );
  INV_X1 NOT1_483( .ZN(N3194), .A(N1932) );
  INV_X1 NOT1_484( .ZN(N3195), .A(N1935) );
  INV_X1 NOT1_485( .ZN(N3196), .A(N1938) );
  INV_X1 NOT1_486( .ZN(N3197), .A(N1941) );
  INV_X1 NOT1_487( .ZN(N3198), .A(N1962) );
  INV_X1 NOT1_488( .ZN(N3199), .A(N1965) );
  BUF_X1 BUFF1_489( .Z(N3200), .A(N1469) );
  INV_X1 NOT1_490( .ZN(N3203), .A(N1968) );
  BUF_X1 BUFF1_491( .Z(N3357), .A(N2704) );
  BUF_X1 BUFF1_492( .Z(N3358), .A(N2704) );
  BUF_X1 BUFF1_493( .Z(N3359), .A(N2704) );
  BUF_X1 BUFF1_494( .Z(N3360), .A(N2704) );
  AND3_X1 AND3_495( .ZN(N3401), .A1(N457), .A2(N1092), .A3(N2824) );
  AND3_X1 AND3_496( .ZN(N3402), .A1(N468), .A2(N1092), .A3(N2826) );
  AND3_X1 AND3_497( .ZN(N3403), .A1(N422), .A2(N1092), .A3(N2828) );
  AND3_X1 AND3_498( .ZN(N3404), .A1(N435), .A2(N1092), .A3(N2830) );
  AND2_X1 AND2_499( .ZN(N3405), .A1(N1080), .A2(N2823) );
  AND2_X1 AND2_500( .ZN(N3406), .A1(N1080), .A2(N2825) );
  AND2_X1 AND2_501( .ZN(N3407), .A1(N1080), .A2(N2827) );
  AND2_X1 AND2_502( .ZN(N3408), .A1(N1080), .A2(N2829) );
  AND3_X1 AND3_503( .ZN(N3409), .A1(N389), .A2(N1092), .A3(N2840) );
  AND3_X1 AND3_504( .ZN(N3410), .A1(N400), .A2(N1092), .A3(N2842) );
  AND3_X1 AND3_505( .ZN(N3411), .A1(N411), .A2(N1092), .A3(N2844) );
  AND3_X1 AND3_506( .ZN(N3412), .A1(N374), .A2(N1092), .A3(N2846) );
  AND2_X1 AND2_507( .ZN(N3413), .A1(N1080), .A2(N2839) );
  AND2_X1 AND2_508( .ZN(N3414), .A1(N1080), .A2(N2841) );
  AND2_X1 AND2_509( .ZN(N3415), .A1(N1080), .A2(N2843) );
  AND2_X1 AND2_510( .ZN(N3416), .A1(N1080), .A2(N2845) );
  AND2_X1 AND2_511( .ZN(N3444), .A1(N1280), .A2(N2902) );
  AND3_X1 AND3_512( .ZN(N3445), .A1(N479), .A2(N1280), .A3(N2904) );
  AND3_X1 AND3_513( .ZN(N3446), .A1(N490), .A2(N1280), .A3(N2906) );
  AND2_X1 AND2_514( .ZN(N3447), .A1(N1685), .A2(N2901) );
  AND2_X1 AND2_515( .ZN(N3448), .A1(N1685), .A2(N2903) );
  AND2_X1 AND2_516( .ZN(N3449), .A1(N1685), .A2(N2905) );
  AND3_X1 AND3_517( .ZN(N3450), .A1(N503), .A2(N1092), .A3(N2914) );
  AND3_X1 AND3_518( .ZN(N3451), .A1(N523), .A2(N1092), .A3(N2916) );
  AND3_X1 AND3_519( .ZN(N3452), .A1(N534), .A2(N1092), .A3(N2918) );
  AND2_X2 AND2_520( .ZN(N3453), .A1(N1080), .A2(N2913) );
  AND2_X2 AND2_521( .ZN(N3454), .A1(N1080), .A2(N2915) );
  AND2_X1 AND2_522( .ZN(N3455), .A1(N1080), .A2(N2917) );
  AND2_X1 AND2_523( .ZN(N3456), .A1(N2920), .A2(N2350) );
  AND3_X1 AND3_524( .ZN(N3459), .A1(N389), .A2(N1280), .A3(N2927) );
  AND3_X1 AND3_525( .ZN(N3460), .A1(N400), .A2(N1280), .A3(N2929) );
  AND3_X1 AND3_526( .ZN(N3461), .A1(N411), .A2(N1280), .A3(N2931) );
  AND3_X1 AND3_527( .ZN(N3462), .A1(N374), .A2(N1280), .A3(N2933) );
  AND2_X1 AND2_528( .ZN(N3463), .A1(N1685), .A2(N2926) );
  AND2_X1 AND2_529( .ZN(N3464), .A1(N1685), .A2(N2928) );
  AND2_X1 AND2_530( .ZN(N3465), .A1(N1685), .A2(N2930) );
  AND2_X1 AND2_531( .ZN(N3466), .A1(N1685), .A2(N2932) );
  AND3_X1 AND3_532( .ZN(N3481), .A1(N503), .A2(N1292), .A3(N2974) );
  INV_X1 NOT1_533( .ZN(N3482), .A(N2980) );
  AND3_X1 AND3_534( .ZN(N3483), .A1(N523), .A2(N1292), .A3(N2976) );
  AND3_X1 AND3_535( .ZN(N3484), .A1(N534), .A2(N1292), .A3(N2978) );
  AND2_X1 AND2_536( .ZN(N3485), .A1(N1271), .A2(N2973) );
  AND2_X1 AND2_537( .ZN(N3486), .A1(N1271), .A2(N2975) );
  AND2_X1 AND2_538( .ZN(N3487), .A1(N1271), .A2(N2977) );
  AND2_X1 AND2_539( .ZN(N3488), .A1(N1292), .A2(N2988) );
  AND3_X1 AND3_540( .ZN(N3489), .A1(N479), .A2(N1292), .A3(N2990) );
  AND3_X2 AND3_541( .ZN(N3490), .A1(N490), .A2(N1292), .A3(N2992) );
  AND2_X2 AND2_542( .ZN(N3491), .A1(N1271), .A2(N2987) );
  AND2_X1 AND2_543( .ZN(N3492), .A1(N1271), .A2(N2989) );
  AND2_X1 AND2_544( .ZN(N3493), .A1(N1271), .A2(N2991) );
  AND2_X1 AND2_545( .ZN(N3502), .A1(N1292), .A2(N2999) );
  AND2_X1 AND2_546( .ZN(N3503), .A1(N1292), .A2(N3006) );
  AND3_X1 AND3_547( .ZN(N3504), .A1(N457), .A2(N1280), .A3(N3016) );
  AND3_X1 AND3_548( .ZN(N3505), .A1(N468), .A2(N1280), .A3(N3018) );
  AND3_X1 AND3_549( .ZN(N3506), .A1(N422), .A2(N1280), .A3(N3020) );
  AND3_X1 AND3_550( .ZN(N3507), .A1(N435), .A2(N1280), .A3(N3022) );
  AND2_X1 AND2_551( .ZN(N3508), .A1(N1685), .A2(N3015) );
  AND2_X1 AND2_552( .ZN(N3509), .A1(N1685), .A2(N3017) );
  AND2_X1 AND2_553( .ZN(N3510), .A1(N1685), .A2(N3019) );
  AND2_X1 AND2_554( .ZN(N3511), .A1(N1685), .A2(N3021) );
  NAND2_X1 NAND2_555( .ZN(N3512), .A1(N1923), .A2(N3031) );
  NAND2_X1 NAND2_556( .ZN(N3513), .A1(N1920), .A2(N3032) );
  NAND2_X1 NAND2_557( .ZN(N3514), .A1(N1929), .A2(N3033) );
  NAND2_X1 NAND2_558( .ZN(N3515), .A1(N1926), .A2(N3034) );
  NAND2_X1 NAND2_559( .ZN(N3558), .A1(N1947), .A2(N3141) );
  NAND2_X1 NAND2_560( .ZN(N3559), .A1(N1944), .A2(N3142) );
  NAND2_X1 NAND2_561( .ZN(N3560), .A1(N1953), .A2(N3143) );
  NAND2_X1 NAND2_562( .ZN(N3561), .A1(N1950), .A2(N3144) );
  NAND2_X1 NAND2_563( .ZN(N3562), .A1(N1959), .A2(N3145) );
  NAND2_X1 NAND2_564( .ZN(N3563), .A1(N1956), .A2(N3146) );
  BUF_X1 BUFF1_565( .Z(N3604), .A(N3191) );
  NAND2_X1 NAND2_566( .ZN(N3605), .A1(N1935), .A2(N3194) );
  NAND2_X1 NAND2_567( .ZN(N3606), .A1(N1932), .A2(N3195) );
  NAND2_X1 NAND2_568( .ZN(N3607), .A1(N1941), .A2(N3196) );
  NAND2_X1 NAND2_569( .ZN(N3608), .A1(N1938), .A2(N3197) );
  NAND2_X1 NAND2_570( .ZN(N3609), .A1(N1965), .A2(N3198) );
  NAND2_X1 NAND2_571( .ZN(N3610), .A1(N1962), .A2(N3199) );
  INV_X1 NOT1_572( .ZN(N3613), .A(N3191) );
  AND2_X1 AND2_573( .ZN(N3614), .A1(N2882), .A2(N2891) );
  AND2_X1 AND2_574( .ZN(N3615), .A1(N1482), .A2(N2891) );
  AND3_X1 AND3_575( .ZN(N3616), .A1(N200), .A2(N2653), .A3(N1173) );
  AND3_X1 AND3_576( .ZN(N3617), .A1(N203), .A2(N2653), .A3(N1173) );
  AND3_X1 AND3_577( .ZN(N3618), .A1(N197), .A2(N2653), .A3(N1173) );
  AND3_X1 AND3_578( .ZN(N3619), .A1(N194), .A2(N2653), .A3(N1173) );
  AND3_X1 AND3_579( .ZN(N3620), .A1(N191), .A2(N2653), .A3(N1173) );
  AND3_X1 AND3_580( .ZN(N3621), .A1(N182), .A2(N2681), .A3(N1197) );
  AND3_X1 AND3_581( .ZN(N3622), .A1(N188), .A2(N2681), .A3(N1197) );
  AND3_X1 AND3_582( .ZN(N3623), .A1(N155), .A2(N2681), .A3(N1197) );
  AND3_X1 AND3_583( .ZN(N3624), .A1(N149), .A2(N2681), .A3(N1197) );
  AND2_X1 AND2_584( .ZN(N3625), .A1(N2882), .A2(N2891) );
  AND2_X1 AND2_585( .ZN(N3626), .A1(N1482), .A2(N2891) );
  AND3_X1 AND3_586( .ZN(N3627), .A1(N200), .A2(N2728), .A3(N1235) );
  AND3_X1 AND3_587( .ZN(N3628), .A1(N203), .A2(N2728), .A3(N1235) );
  AND3_X1 AND3_588( .ZN(N3629), .A1(N197), .A2(N2728), .A3(N1235) );
  AND3_X1 AND3_589( .ZN(N3630), .A1(N194), .A2(N2728), .A3(N1235) );
  AND3_X1 AND3_590( .ZN(N3631), .A1(N191), .A2(N2728), .A3(N1235) );
  AND3_X1 AND3_591( .ZN(N3632), .A1(N182), .A2(N2756), .A3(N1259) );
  AND3_X1 AND3_592( .ZN(N3633), .A1(N188), .A2(N2756), .A3(N1259) );
  AND3_X1 AND3_593( .ZN(N3634), .A1(N155), .A2(N2756), .A3(N1259) );
  AND3_X1 AND3_594( .ZN(N3635), .A1(N149), .A2(N2756), .A3(N1259) );
  AND2_X1 AND2_595( .ZN(N3636), .A1(N2882), .A2(N2891) );
  AND2_X1 AND2_596( .ZN(N3637), .A1(N1482), .A2(N2891) );
  AND3_X1 AND3_597( .ZN(N3638), .A1(N109), .A2(N3075), .A3(N1743) );
  AND2_X1 AND2_598( .ZN(N3639), .A1(N2882), .A2(N2891) );
  AND2_X1 AND2_599( .ZN(N3640), .A1(N1482), .A2(N2891) );
  AND3_X1 AND3_600( .ZN(N3641), .A1(N11), .A2(N2779), .A3(N1339) );
  AND3_X1 AND3_601( .ZN(N3642), .A1(N109), .A2(N3041), .A3(N1709) );
  AND3_X1 AND3_602( .ZN(N3643), .A1(N46), .A2(N3041), .A3(N1709) );
  AND3_X1 AND3_603( .ZN(N3644), .A1(N100), .A2(N3041), .A3(N1709) );
  AND3_X1 AND3_604( .ZN(N3645), .A1(N91), .A2(N3041), .A3(N1709) );
  AND3_X1 AND3_605( .ZN(N3646), .A1(N43), .A2(N3041), .A3(N1709) );
  AND3_X2 AND3_606( .ZN(N3647), .A1(N76), .A2(N2779), .A3(N1339) );
  AND3_X2 AND3_607( .ZN(N3648), .A1(N73), .A2(N2779), .A3(N1339) );
  AND3_X1 AND3_608( .ZN(N3649), .A1(N67), .A2(N2779), .A3(N1339) );
  AND3_X1 AND3_609( .ZN(N3650), .A1(N14), .A2(N2779), .A3(N1339) );
  AND3_X1 AND3_610( .ZN(N3651), .A1(N46), .A2(N3075), .A3(N1743) );
  AND3_X1 AND3_611( .ZN(N3652), .A1(N100), .A2(N3075), .A3(N1743) );
  AND3_X1 AND3_612( .ZN(N3653), .A1(N91), .A2(N3075), .A3(N1743) );
  AND3_X1 AND3_613( .ZN(N3654), .A1(N43), .A2(N3075), .A3(N1743) );
  AND3_X1 AND3_614( .ZN(N3655), .A1(N76), .A2(N2801), .A3(N1363) );
  AND3_X1 AND3_615( .ZN(N3656), .A1(N73), .A2(N2801), .A3(N1363) );
  AND3_X1 AND3_616( .ZN(N3657), .A1(N67), .A2(N2801), .A3(N1363) );
  AND3_X1 AND3_617( .ZN(N3658), .A1(N14), .A2(N2801), .A3(N1363) );
  AND3_X1 AND3_618( .ZN(N3659), .A1(N120), .A2(N3119), .A3(N1785) );
  AND3_X1 AND3_619( .ZN(N3660), .A1(N11), .A2(N2801), .A3(N1363) );
  AND3_X1 AND3_620( .ZN(N3661), .A1(N118), .A2(N3097), .A3(N1769) );
  AND3_X1 AND3_621( .ZN(N3662), .A1(N176), .A2(N2681), .A3(N1197) );
  AND3_X1 AND3_622( .ZN(N3663), .A1(N176), .A2(N2756), .A3(N1259) );
  OR2_X2 OR2_623( .ZN(N3664), .A1(N2831), .A2(N3401) );
  OR2_X1 OR2_624( .ZN(N3665), .A1(N2832), .A2(N3402) );
  OR2_X1 OR2_625( .ZN(N3666), .A1(N2833), .A2(N3403) );
  OR2_X1 OR2_626( .ZN(N3667), .A1(N2834), .A2(N3404) );
  OR3_X1 OR3_627( .ZN(N3668), .A1(N2835), .A2(N3405), .A3(N457) );
  OR3_X1 OR3_628( .ZN(N3669), .A1(N2836), .A2(N3406), .A3(N468) );
  OR3_X1 OR3_629( .ZN(N3670), .A1(N2837), .A2(N3407), .A3(N422) );
  OR3_X1 OR3_630( .ZN(N3671), .A1(N2838), .A2(N3408), .A3(N435) );
  OR2_X1 OR2_631( .ZN(N3672), .A1(N2847), .A2(N3409) );
  OR2_X1 OR2_632( .ZN(N3673), .A1(N2848), .A2(N3410) );
  OR2_X1 OR2_633( .ZN(N3674), .A1(N2849), .A2(N3411) );
  OR2_X1 OR2_634( .ZN(N3675), .A1(N2850), .A2(N3412) );
  OR3_X4 OR3_635( .ZN(N3676), .A1(N2851), .A2(N3413), .A3(N389) );
  OR3_X1 OR3_636( .ZN(N3677), .A1(N2852), .A2(N3414), .A3(N400) );
  OR3_X1 OR3_637( .ZN(N3678), .A1(N2853), .A2(N3415), .A3(N411) );
  OR3_X1 OR3_638( .ZN(N3679), .A1(N2854), .A2(N3416), .A3(N374) );
  AND2_X1 AND2_639( .ZN(N3680), .A1(N289), .A2(N2855) );
  AND2_X1 AND2_640( .ZN(N3681), .A1(N281), .A2(N2855) );
  AND2_X1 AND2_641( .ZN(N3682), .A1(N273), .A2(N2855) );
  AND2_X1 AND2_642( .ZN(N3683), .A1(N265), .A2(N2855) );
  AND2_X1 AND2_643( .ZN(N3684), .A1(N257), .A2(N2855) );
  AND2_X1 AND2_644( .ZN(N3685), .A1(N234), .A2(N2861) );
  AND2_X1 AND2_645( .ZN(N3686), .A1(N226), .A2(N2861) );
  AND2_X1 AND2_646( .ZN(N3687), .A1(N218), .A2(N2861) );
  AND2_X1 AND2_647( .ZN(N3688), .A1(N210), .A2(N2861) );
  AND2_X1 AND2_648( .ZN(N3689), .A1(N206), .A2(N2861) );
  INV_X1 NOT1_649( .ZN(N3691), .A(N2891) );
  OR2_X1 OR2_650( .ZN(N3700), .A1(N2907), .A2(N3444) );
  OR2_X1 OR2_651( .ZN(N3701), .A1(N2908), .A2(N3445) );
  OR2_X1 OR2_652( .ZN(N3702), .A1(N2909), .A2(N3446) );
  OR3_X1 OR3_653( .ZN(N3703), .A1(N2911), .A2(N3448), .A3(N479) );
  OR3_X1 OR3_654( .ZN(N3704), .A1(N2912), .A2(N3449), .A3(N490) );
  OR2_X1 OR2_655( .ZN(N3705), .A1(N2910), .A2(N3447) );
  OR2_X1 OR2_656( .ZN(N3708), .A1(N2919), .A2(N3450) );
  OR2_X1 OR2_657( .ZN(N3709), .A1(N2921), .A2(N3451) );
  OR2_X1 OR2_658( .ZN(N3710), .A1(N2922), .A2(N3452) );
  OR3_X1 OR3_659( .ZN(N3711), .A1(N2923), .A2(N3453), .A3(N503) );
  OR3_X1 OR3_660( .ZN(N3712), .A1(N2924), .A2(N3454), .A3(N523) );
  OR3_X1 OR3_661( .ZN(N3713), .A1(N2925), .A2(N3455), .A3(N534) );
  OR2_X1 OR2_662( .ZN(N3715), .A1(N2934), .A2(N3459) );
  OR2_X1 OR2_663( .ZN(N3716), .A1(N2935), .A2(N3460) );
  OR2_X1 OR2_664( .ZN(N3717), .A1(N2936), .A2(N3461) );
  OR2_X1 OR2_665( .ZN(N3718), .A1(N2937), .A2(N3462) );
  OR3_X1 OR3_666( .ZN(N3719), .A1(N2938), .A2(N3463), .A3(N389) );
  OR3_X1 OR3_667( .ZN(N3720), .A1(N2939), .A2(N3464), .A3(N400) );
  OR3_X1 OR3_668( .ZN(N3721), .A1(N2940), .A2(N3465), .A3(N411) );
  OR3_X1 OR3_669( .ZN(N3722), .A1(N2941), .A2(N3466), .A3(N374) );
  AND2_X1 AND2_670( .ZN(N3723), .A1(N369), .A2(N2942) );
  AND2_X1 AND2_671( .ZN(N3724), .A1(N361), .A2(N2942) );
  AND2_X1 AND2_672( .ZN(N3725), .A1(N351), .A2(N2942) );
  AND2_X1 AND2_673( .ZN(N3726), .A1(N341), .A2(N2942) );
  AND2_X1 AND2_674( .ZN(N3727), .A1(N324), .A2(N2948) );
  AND2_X1 AND2_675( .ZN(N3728), .A1(N316), .A2(N2948) );
  AND2_X1 AND2_676( .ZN(N3729), .A1(N308), .A2(N2948) );
  AND2_X1 AND2_677( .ZN(N3730), .A1(N302), .A2(N2948) );
  AND2_X1 AND2_678( .ZN(N3731), .A1(N293), .A2(N2948) );
  OR2_X1 OR2_679( .ZN(N3732), .A1(N2942), .A2(N2958) );
  AND2_X1 AND2_680( .ZN(N3738), .A1(N83), .A2(N2964) );
  AND2_X1 AND2_681( .ZN(N3739), .A1(N87), .A2(N2964) );
  AND2_X1 AND2_682( .ZN(N3740), .A1(N34), .A2(N2964) );
  AND2_X1 AND2_683( .ZN(N3741), .A1(N34), .A2(N2964) );
  OR2_X1 OR2_684( .ZN(N3742), .A1(N2979), .A2(N3481) );
  OR2_X1 OR2_685( .ZN(N3743), .A1(N2981), .A2(N3483) );
  OR2_X1 OR2_686( .ZN(N3744), .A1(N2982), .A2(N3484) );
  OR3_X1 OR3_687( .ZN(N3745), .A1(N2983), .A2(N3485), .A3(N503) );
  OR3_X1 OR3_688( .ZN(N3746), .A1(N2985), .A2(N3486), .A3(N523) );
  OR3_X1 OR3_689( .ZN(N3747), .A1(N2986), .A2(N3487), .A3(N534) );
  OR2_X1 OR2_690( .ZN(N3748), .A1(N2993), .A2(N3488) );
  OR2_X1 OR2_691( .ZN(N3749), .A1(N2994), .A2(N3489) );
  OR2_X1 OR2_692( .ZN(N3750), .A1(N2995), .A2(N3490) );
  OR3_X1 OR3_693( .ZN(N3751), .A1(N2997), .A2(N3492), .A3(N479) );
  OR3_X1 OR3_694( .ZN(N3752), .A1(N2998), .A2(N3493), .A3(N490) );
  INV_X1 NOT1_695( .ZN(N3753), .A(N3000) );
  INV_X1 NOT1_696( .ZN(N3754), .A(N3003) );
  INV_X1 NOT1_697( .ZN(N3755), .A(N3007) );
  INV_X1 NOT1_698( .ZN(N3756), .A(N3010) );
  OR2_X1 OR2_699( .ZN(N3757), .A1(N3013), .A2(N3502) );
  AND3_X1 AND3_700( .ZN(N3758), .A1(N1315), .A2(N446), .A3(N3003) );
  OR2_X1 OR2_701( .ZN(N3759), .A1(N3014), .A2(N3503) );
  AND3_X1 AND3_702( .ZN(N3760), .A1(N1315), .A2(N446), .A3(N3010) );
  AND2_X1 AND2_703( .ZN(N3761), .A1(N1675), .A2(N3000) );
  AND2_X1 AND2_704( .ZN(N3762), .A1(N1675), .A2(N3007) );
  OR2_X1 OR2_705( .ZN(N3763), .A1(N3023), .A2(N3504) );
  OR2_X1 OR2_706( .ZN(N3764), .A1(N3024), .A2(N3505) );
  OR2_X1 OR2_707( .ZN(N3765), .A1(N3025), .A2(N3506) );
  OR2_X1 OR2_708( .ZN(N3766), .A1(N3026), .A2(N3507) );
  OR3_X1 OR3_709( .ZN(N3767), .A1(N3027), .A2(N3508), .A3(N457) );
  OR3_X2 OR3_710( .ZN(N3768), .A1(N3028), .A2(N3509), .A3(N468) );
  OR3_X1 OR3_711( .ZN(N3769), .A1(N3029), .A2(N3510), .A3(N422) );
  OR3_X1 OR3_712( .ZN(N3770), .A1(N3030), .A2(N3511), .A3(N435) );
  NAND2_X1 NAND2_713( .ZN(N3771), .A1(N3512), .A2(N3513) );
  NAND2_X1 NAND2_714( .ZN(N3775), .A1(N3514), .A2(N3515) );
  INV_X1 NOT1_715( .ZN(N3779), .A(N3035) );
  INV_X1 NOT1_716( .ZN(N3780), .A(N3038) );
  AND3_X1 AND3_717( .ZN(N3781), .A1(N117), .A2(N3097), .A3(N1769) );
  AND3_X1 AND3_718( .ZN(N3782), .A1(N126), .A2(N3097), .A3(N1769) );
  AND3_X1 AND3_719( .ZN(N3783), .A1(N127), .A2(N3097), .A3(N1769) );
  AND3_X1 AND3_720( .ZN(N3784), .A1(N128), .A2(N3097), .A3(N1769) );
  AND3_X2 AND3_721( .ZN(N3785), .A1(N131), .A2(N3119), .A3(N1785) );
  AND3_X2 AND3_722( .ZN(N3786), .A1(N129), .A2(N3119), .A3(N1785) );
  AND3_X1 AND3_723( .ZN(N3787), .A1(N119), .A2(N3119), .A3(N1785) );
  AND3_X1 AND3_724( .ZN(N3788), .A1(N130), .A2(N3119), .A3(N1785) );
  NAND2_X1 NAND2_725( .ZN(N3789), .A1(N3558), .A2(N3559) );
  NAND2_X1 NAND2_726( .ZN(N3793), .A1(N3560), .A2(N3561) );
  NAND2_X1 NAND2_727( .ZN(N3797), .A1(N3562), .A2(N3563) );
  AND3_X1 AND3_728( .ZN(N3800), .A1(N122), .A2(N3147), .A3(N1800) );
  AND3_X1 AND3_729( .ZN(N3801), .A1(N113), .A2(N3147), .A3(N1800) );
  AND3_X1 AND3_730( .ZN(N3802), .A1(N53), .A2(N3147), .A3(N1800) );
  AND3_X1 AND3_731( .ZN(N3803), .A1(N114), .A2(N3147), .A3(N1800) );
  AND3_X1 AND3_732( .ZN(N3804), .A1(N115), .A2(N3147), .A3(N1800) );
  AND3_X1 AND3_733( .ZN(N3805), .A1(N52), .A2(N3169), .A3(N1814) );
  AND3_X1 AND3_734( .ZN(N3806), .A1(N112), .A2(N3169), .A3(N1814) );
  AND3_X1 AND3_735( .ZN(N3807), .A1(N116), .A2(N3169), .A3(N1814) );
  AND3_X1 AND3_736( .ZN(N3808), .A1(N121), .A2(N3169), .A3(N1814) );
  AND3_X1 AND3_737( .ZN(N3809), .A1(N123), .A2(N3169), .A3(N1814) );
  NAND2_X1 NAND2_738( .ZN(N3810), .A1(N3607), .A2(N3608) );
  NAND2_X1 NAND2_739( .ZN(N3813), .A1(N3605), .A2(N3606) );
  AND2_X1 AND2_740( .ZN(N3816), .A1(N3482), .A2(N2984) );
  OR2_X1 OR2_741( .ZN(N3819), .A1(N2996), .A2(N3491) );
  INV_X1 NOT1_742( .ZN(N3822), .A(N3200) );
  NAND2_X1 NAND2_743( .ZN(N3823), .A1(N3200), .A2(N3203) );
  NAND2_X1 NAND2_744( .ZN(N3824), .A1(N3609), .A2(N3610) );
  INV_X1 NOT1_745( .ZN(N3827), .A(N3456) );
  OR2_X1 OR2_746( .ZN(N3828), .A1(N3739), .A2(N2970) );
  OR2_X1 OR2_747( .ZN(N3829), .A1(N3740), .A2(N2971) );
  OR2_X1 OR2_748( .ZN(N3830), .A1(N3741), .A2(N2972) );
  OR2_X1 OR2_749( .ZN(N3831), .A1(N3738), .A2(N2969) );
  INV_X1 NOT1_750( .ZN(N3834), .A(N3664) );
  INV_X1 NOT1_751( .ZN(N3835), .A(N3665) );
  INV_X1 NOT1_752( .ZN(N3836), .A(N3666) );
  INV_X1 NOT1_753( .ZN(N3837), .A(N3667) );
  INV_X1 NOT1_754( .ZN(N3838), .A(N3672) );
  INV_X1 NOT1_755( .ZN(N3839), .A(N3673) );
  INV_X1 NOT1_756( .ZN(N3840), .A(N3674) );
  INV_X1 NOT1_757( .ZN(N3841), .A(N3675) );
  OR2_X1 OR2_758( .ZN(N3842), .A1(N3681), .A2(N2868) );
  OR2_X1 OR2_759( .ZN(N3849), .A1(N3682), .A2(N2869) );
  OR2_X1 OR2_760( .ZN(N3855), .A1(N3683), .A2(N2870) );
  OR2_X1 OR2_761( .ZN(N3861), .A1(N3684), .A2(N2871) );
  OR2_X1 OR2_762( .ZN(N3867), .A1(N3685), .A2(N2872) );
  OR2_X1 OR2_763( .ZN(N3873), .A1(N3686), .A2(N2873) );
  OR2_X1 OR2_764( .ZN(N3881), .A1(N3687), .A2(N2874) );
  OR2_X1 OR2_765( .ZN(N3887), .A1(N3688), .A2(N2875) );
  OR2_X1 OR2_766( .ZN(N3893), .A1(N3689), .A2(N2876) );
  INV_X1 NOT1_767( .ZN(N3908), .A(N3701) );
  INV_X1 NOT1_768( .ZN(N3909), .A(N3702) );
  INV_X1 NOT1_769( .ZN(N3911), .A(N3700) );
  INV_X1 NOT1_770( .ZN(N3914), .A(N3708) );
  INV_X1 NOT1_771( .ZN(N3915), .A(N3709) );
  INV_X1 NOT1_772( .ZN(N3916), .A(N3710) );
  INV_X1 NOT1_773( .ZN(N3917), .A(N3715) );
  INV_X1 NOT1_774( .ZN(N3918), .A(N3716) );
  INV_X1 NOT1_775( .ZN(N3919), .A(N3717) );
  INV_X1 NOT1_776( .ZN(N3920), .A(N3718) );
  OR2_X1 OR2_777( .ZN(N3921), .A1(N3724), .A2(N2955) );
  OR2_X1 OR2_778( .ZN(N3927), .A1(N3725), .A2(N2956) );
  OR2_X1 OR2_779( .ZN(N3933), .A1(N3726), .A2(N2957) );
  OR2_X1 OR2_780( .ZN(N3942), .A1(N3727), .A2(N2959) );
  OR2_X1 OR2_781( .ZN(N3948), .A1(N3728), .A2(N2960) );
  OR2_X1 OR2_782( .ZN(N3956), .A1(N3729), .A2(N2961) );
  OR2_X1 OR2_783( .ZN(N3962), .A1(N3730), .A2(N2962) );
  OR2_X1 OR2_784( .ZN(N3968), .A1(N3731), .A2(N2963) );
  INV_X1 NOT1_785( .ZN(N3975), .A(N3742) );
  INV_X1 NOT1_786( .ZN(N3976), .A(N3743) );
  INV_X1 NOT1_787( .ZN(N3977), .A(N3744) );
  INV_X1 NOT1_788( .ZN(N3978), .A(N3749) );
  INV_X1 NOT1_789( .ZN(N3979), .A(N3750) );
  AND3_X1 AND3_790( .ZN(N3980), .A1(N446), .A2(N1292), .A3(N3754) );
  AND3_X1 AND3_791( .ZN(N3981), .A1(N446), .A2(N1292), .A3(N3756) );
  AND2_X1 AND2_792( .ZN(N3982), .A1(N1271), .A2(N3753) );
  AND2_X1 AND2_793( .ZN(N3983), .A1(N1271), .A2(N3755) );
  INV_X1 NOT1_794( .ZN(N3984), .A(N3757) );
  INV_X1 NOT1_795( .ZN(N3987), .A(N3759) );
  INV_X1 NOT1_796( .ZN(N3988), .A(N3763) );
  INV_X1 NOT1_797( .ZN(N3989), .A(N3764) );
  INV_X1 NOT1_798( .ZN(N3990), .A(N3765) );
  INV_X1 NOT1_799( .ZN(N3991), .A(N3766) );
  AND3_X1 AND3_800( .ZN(N3998), .A1(N3456), .A2(N3119), .A3(N3130) );
  OR2_X1 OR2_801( .ZN(N4008), .A1(N3723), .A2(N2954) );
  OR2_X1 OR2_802( .ZN(N4011), .A1(N3680), .A2(N2867) );
  INV_X1 NOT1_803( .ZN(N4021), .A(N3748) );
  NAND2_X1 NAND2_804( .ZN(N4024), .A1(N1968), .A2(N3822) );
  INV_X1 NOT1_805( .ZN(N4027), .A(N3705) );
  AND2_X1 AND2_806( .ZN(N4031), .A1(N3828), .A2(N1583) );
  AND3_X1 AND3_807( .ZN(N4032), .A1(N24), .A2(N2882), .A3(N3691) );
  AND3_X1 AND3_808( .ZN(N4033), .A1(N25), .A2(N1482), .A3(N3691) );
  AND3_X1 AND3_809( .ZN(N4034), .A1(N26), .A2(N2882), .A3(N3691) );
  AND3_X1 AND3_810( .ZN(N4035), .A1(N81), .A2(N1482), .A3(N3691) );
  AND2_X1 AND2_811( .ZN(N4036), .A1(N3829), .A2(N1583) );
  AND3_X1 AND3_812( .ZN(N4037), .A1(N79), .A2(N2882), .A3(N3691) );
  AND3_X1 AND3_813( .ZN(N4038), .A1(N23), .A2(N1482), .A3(N3691) );
  AND3_X2 AND3_814( .ZN(N4039), .A1(N82), .A2(N2882), .A3(N3691) );
  AND3_X2 AND3_815( .ZN(N4040), .A1(N80), .A2(N1482), .A3(N3691) );
  AND2_X1 AND2_816( .ZN(N4041), .A1(N3830), .A2(N1583) );
  AND2_X1 AND2_817( .ZN(N4042), .A1(N3831), .A2(N1583) );
  AND2_X1 AND2_818( .ZN(N4067), .A1(N3732), .A2(N514) );
  AND2_X1 AND2_819( .ZN(N4080), .A1(N514), .A2(N3732) );
  AND2_X1 AND2_820( .ZN(N4088), .A1(N3834), .A2(N3668) );
  AND2_X1 AND2_821( .ZN(N4091), .A1(N3835), .A2(N3669) );
  AND2_X1 AND2_822( .ZN(N4094), .A1(N3836), .A2(N3670) );
  AND2_X1 AND2_823( .ZN(N4097), .A1(N3837), .A2(N3671) );
  AND2_X1 AND2_824( .ZN(N4100), .A1(N3838), .A2(N3676) );
  AND2_X1 AND2_825( .ZN(N4103), .A1(N3839), .A2(N3677) );
  AND2_X1 AND2_826( .ZN(N4106), .A1(N3840), .A2(N3678) );
  AND2_X1 AND2_827( .ZN(N4109), .A1(N3841), .A2(N3679) );
  AND2_X1 AND2_828( .ZN(N4144), .A1(N3908), .A2(N3703) );
  AND2_X1 AND2_829( .ZN(N4147), .A1(N3909), .A2(N3704) );
  BUF_X1 BUFF1_830( .Z(N4150), .A(N3705) );
  AND2_X1 AND2_831( .ZN(N4153), .A1(N3914), .A2(N3711) );
  AND2_X1 AND2_832( .ZN(N4156), .A1(N3915), .A2(N3712) );
  AND2_X1 AND2_833( .ZN(N4159), .A1(N3916), .A2(N3713) );
  OR2_X1 OR2_834( .ZN(N4183), .A1(N3758), .A2(N3980) );
  OR2_X1 OR2_835( .ZN(N4184), .A1(N3760), .A2(N3981) );
  OR3_X1 OR3_836( .ZN(N4185), .A1(N3761), .A2(N3982), .A3(N446) );
  OR3_X1 OR3_837( .ZN(N4186), .A1(N3762), .A2(N3983), .A3(N446) );
  INV_X1 NOT1_838( .ZN(N4188), .A(N3771) );
  INV_X1 NOT1_839( .ZN(N4191), .A(N3775) );
  AND3_X1 AND3_840( .ZN(N4196), .A1(N3775), .A2(N3771), .A3(N3035) );
  AND3_X1 AND3_841( .ZN(N4197), .A1(N3987), .A2(N3119), .A3(N3130) );
  AND2_X1 AND2_842( .ZN(N4198), .A1(N3920), .A2(N3722) );
  INV_X1 NOT1_843( .ZN(N4199), .A(N3816) );
  INV_X1 NOT1_844( .ZN(N4200), .A(N3789) );
  INV_X1 NOT1_845( .ZN(N4203), .A(N3793) );
  BUF_X1 BUFF1_846( .Z(N4206), .A(N3797) );
  BUF_X1 BUFF1_847( .Z(N4209), .A(N3797) );
  BUF_X1 BUFF1_848( .Z(N4212), .A(N3732) );
  BUF_X1 BUFF1_849( .Z(N4215), .A(N3732) );
  BUF_X1 BUFF1_850( .Z(N4219), .A(N3732) );
  INV_X1 NOT1_851( .ZN(N4223), .A(N3810) );
  INV_X1 NOT1_852( .ZN(N4224), .A(N3813) );
  AND2_X1 AND2_853( .ZN(N4225), .A1(N3918), .A2(N3720) );
  AND2_X1 AND2_854( .ZN(N4228), .A1(N3919), .A2(N3721) );
  AND2_X1 AND2_855( .ZN(N4231), .A1(N3991), .A2(N3770) );
  AND2_X1 AND2_856( .ZN(N4234), .A1(N3917), .A2(N3719) );
  AND2_X1 AND2_857( .ZN(N4237), .A1(N3989), .A2(N3768) );
  AND2_X1 AND2_858( .ZN(N4240), .A1(N3990), .A2(N3769) );
  AND2_X1 AND2_859( .ZN(N4243), .A1(N3988), .A2(N3767) );
  AND2_X1 AND2_860( .ZN(N4246), .A1(N3976), .A2(N3746) );
  AND2_X1 AND2_861( .ZN(N4249), .A1(N3977), .A2(N3747) );
  AND2_X1 AND2_862( .ZN(N4252), .A1(N3975), .A2(N3745) );
  AND2_X1 AND2_863( .ZN(N4255), .A1(N3978), .A2(N3751) );
  AND2_X1 AND2_864( .ZN(N4258), .A1(N3979), .A2(N3752) );
  INV_X1 NOT1_865( .ZN(N4263), .A(N3819) );
  NAND2_X1 NAND2_866( .ZN(N4264), .A1(N4024), .A2(N3823) );
  INV_X1 NOT1_867( .ZN(N4267), .A(N3824) );
  AND2_X1 AND2_868( .ZN(N4268), .A1(N446), .A2(N3893) );
  INV_X1 NOT1_869( .ZN(N4269), .A(N3911) );
  INV_X1 NOT1_870( .ZN(N4270), .A(N3984) );
  AND2_X1 AND2_871( .ZN(N4271), .A1(N3893), .A2(N446) );
  INV_X1 NOT1_872( .ZN(N4272), .A(N4031) );
  OR4_X1 OR4_873( .ZN(N4273), .A1(N4032), .A2(N4033), .A3(N3614), .A4(N3615) );
  OR4_X1 OR4_874( .ZN(N4274), .A1(N4034), .A2(N4035), .A3(N3625), .A4(N3626) );
  INV_X1 NOT1_875( .ZN(N4275), .A(N4036) );
  OR4_X1 OR4_876( .ZN(N4276), .A1(N4037), .A2(N4038), .A3(N3636), .A4(N3637) );
  OR4_X1 OR4_877( .ZN(N4277), .A1(N4039), .A2(N4040), .A3(N3639), .A4(N3640) );
  INV_X1 NOT1_878( .ZN(N4278), .A(N4041) );
  INV_X1 NOT1_879( .ZN(N4279), .A(N4042) );
  AND2_X1 AND2_880( .ZN(N4280), .A1(N3887), .A2(N457) );
  AND2_X1 AND2_881( .ZN(N4284), .A1(N3881), .A2(N468) );
  AND2_X1 AND2_882( .ZN(N4290), .A1(N422), .A2(N3873) );
  AND2_X1 AND2_883( .ZN(N4297), .A1(N3867), .A2(N435) );
  AND2_X1 AND2_884( .ZN(N4298), .A1(N3861), .A2(N389) );
  AND2_X2 AND2_885( .ZN(N4301), .A1(N3855), .A2(N400) );
  AND2_X2 AND2_886( .ZN(N4305), .A1(N3849), .A2(N411) );
  AND2_X1 AND2_887( .ZN(N4310), .A1(N3842), .A2(N374) );
  AND2_X1 AND2_888( .ZN(N4316), .A1(N457), .A2(N3887) );
  AND2_X1 AND2_889( .ZN(N4320), .A1(N468), .A2(N3881) );
  AND2_X1 AND2_890( .ZN(N4325), .A1(N422), .A2(N3873) );
  AND2_X1 AND2_891( .ZN(N4331), .A1(N435), .A2(N3867) );
  AND2_X1 AND2_892( .ZN(N4332), .A1(N389), .A2(N3861) );
  AND2_X1 AND2_893( .ZN(N4336), .A1(N400), .A2(N3855) );
  AND2_X1 AND2_894( .ZN(N4342), .A1(N411), .A2(N3849) );
  AND2_X1 AND2_895( .ZN(N4349), .A1(N374), .A2(N3842) );
  INV_X1 NOT1_896( .ZN(N4357), .A(N3968) );
  INV_X1 NOT1_897( .ZN(N4364), .A(N3962) );
  BUF_X4 BUFF1_898( .Z(N4375), .A(N3962) );
  AND2_X1 AND2_899( .ZN(N4379), .A1(N3956), .A2(N479) );
  AND2_X1 AND2_900( .ZN(N4385), .A1(N490), .A2(N3948) );
  AND2_X1 AND2_901( .ZN(N4392), .A1(N3942), .A2(N503) );
  AND2_X1 AND2_902( .ZN(N4396), .A1(N3933), .A2(N523) );
  AND2_X1 AND2_903( .ZN(N4400), .A1(N3927), .A2(N534) );
  INV_X1 NOT1_904( .ZN(N4405), .A(N3921) );
  BUF_X1 BUFF1_905( .Z(N4412), .A(N3921) );
  INV_X1 NOT1_906( .ZN(N4418), .A(N3968) );
  INV_X1 NOT1_907( .ZN(N4425), .A(N3962) );
  BUF_X1 BUFF1_908( .Z(N4436), .A(N3962) );
  AND2_X1 AND2_909( .ZN(N4440), .A1(N479), .A2(N3956) );
  AND2_X1 AND2_910( .ZN(N4445), .A1(N490), .A2(N3948) );
  AND2_X1 AND2_911( .ZN(N4451), .A1(N503), .A2(N3942) );
  AND2_X1 AND2_912( .ZN(N4456), .A1(N523), .A2(N3933) );
  AND2_X1 AND2_913( .ZN(N4462), .A1(N534), .A2(N3927) );
  BUF_X1 BUFF1_914( .Z(N4469), .A(N3921) );
  INV_X1 NOT1_915( .ZN(N4477), .A(N3921) );
  BUF_X1 BUFF1_916( .Z(N4512), .A(N3968) );
  INV_X1 NOT1_917( .ZN(N4515), .A(N4183) );
  INV_X1 NOT1_918( .ZN(N4516), .A(N4184) );
  INV_X1 NOT1_919( .ZN(N4521), .A(N4008) );
  INV_X4 NOT1_920( .ZN(N4523), .A(N4011) );
  INV_X1 NOT1_921( .ZN(N4524), .A(N4198) );
  INV_X1 NOT1_922( .ZN(N4532), .A(N3984) );
  AND3_X1 AND3_923( .ZN(N4547), .A1(N3911), .A2(N3169), .A3(N3180) );
  BUF_X1 BUFF1_924( .Z(N4548), .A(N3893) );
  BUF_X1 BUFF1_925( .Z(N4551), .A(N3887) );
  BUF_X1 BUFF1_926( .Z(N4554), .A(N3881) );
  BUF_X4 BUFF1_927( .Z(N4557), .A(N3873) );
  BUF_X1 BUFF1_928( .Z(N4560), .A(N3867) );
  BUF_X1 BUFF1_929( .Z(N4563), .A(N3861) );
  BUF_X1 BUFF1_930( .Z(N4566), .A(N3855) );
  BUF_X1 BUFF1_931( .Z(N4569), .A(N3849) );
  BUF_X1 BUFF1_932( .Z(N4572), .A(N3842) );
  NOR2_X1 NOR2_933( .ZN(N4575), .A1(N422), .A2(N3873) );
  BUF_X1 BUFF1_934( .Z(N4578), .A(N3893) );
  BUF_X1 BUFF1_935( .Z(N4581), .A(N3887) );
  BUF_X1 BUFF1_936( .Z(N4584), .A(N3881) );
  BUF_X1 BUFF1_937( .Z(N4587), .A(N3867) );
  BUF_X1 BUFF1_938( .Z(N4590), .A(N3861) );
  BUF_X1 BUFF1_939( .Z(N4593), .A(N3855) );
  BUF_X1 BUFF1_940( .Z(N4596), .A(N3849) );
  BUF_X1 BUFF1_941( .Z(N4599), .A(N3873) );
  BUF_X1 BUFF1_942( .Z(N4602), .A(N3842) );
  NOR2_X1 NOR2_943( .ZN(N4605), .A1(N422), .A2(N3873) );
  NOR2_X1 NOR2_944( .ZN(N4608), .A1(N374), .A2(N3842) );
  BUF_X1 BUFF1_945( .Z(N4611), .A(N3956) );
  BUF_X1 BUFF1_946( .Z(N4614), .A(N3948) );
  BUF_X1 BUFF1_947( .Z(N4617), .A(N3942) );
  BUF_X1 BUFF1_948( .Z(N4621), .A(N3933) );
  BUF_X1 BUFF1_949( .Z(N4624), .A(N3927) );
  NOR2_X1 NOR2_950( .ZN(N4627), .A1(N490), .A2(N3948) );
  BUF_X1 BUFF1_951( .Z(N4630), .A(N3956) );
  BUF_X1 BUFF1_952( .Z(N4633), .A(N3942) );
  BUF_X1 BUFF1_953( .Z(N4637), .A(N3933) );
  BUF_X1 BUFF1_954( .Z(N4640), .A(N3927) );
  BUF_X1 BUFF1_955( .Z(N4643), .A(N3948) );
  NOR2_X1 NOR2_956( .ZN(N4646), .A1(N490), .A2(N3948) );
  BUF_X1 BUFF1_957( .Z(N4649), .A(N3927) );
  BUF_X1 BUFF1_958( .Z(N4652), .A(N3933) );
  BUF_X1 BUFF1_959( .Z(N4655), .A(N3921) );
  BUF_X1 BUFF1_960( .Z(N4658), .A(N3942) );
  BUF_X1 BUFF1_961( .Z(N4662), .A(N3956) );
  BUF_X1 BUFF1_962( .Z(N4665), .A(N3948) );
  BUF_X1 BUFF1_963( .Z(N4668), .A(N3968) );
  BUF_X1 BUFF1_964( .Z(N4671), .A(N3962) );
  BUF_X1 BUFF1_965( .Z(N4674), .A(N3873) );
  BUF_X1 BUFF1_966( .Z(N4677), .A(N3867) );
  BUF_X1 BUFF1_967( .Z(N4680), .A(N3887) );
  BUF_X1 BUFF1_968( .Z(N4683), .A(N3881) );
  BUF_X1 BUFF1_969( .Z(N4686), .A(N3893) );
  BUF_X1 BUFF1_970( .Z(N4689), .A(N3849) );
  BUF_X1 BUFF1_971( .Z(N4692), .A(N3842) );
  BUF_X1 BUFF1_972( .Z(N4695), .A(N3861) );
  BUF_X1 BUFF1_973( .Z(N4698), .A(N3855) );
  NAND2_X1 NAND2_974( .ZN(N4701), .A1(N3813), .A2(N4223) );
  NAND2_X1 NAND2_975( .ZN(N4702), .A1(N3810), .A2(N4224) );
  INV_X1 NOT1_976( .ZN(N4720), .A(N4021) );
  NAND2_X1 NAND2_977( .ZN(N4721), .A1(N4021), .A2(N4263) );
  INV_X1 NOT1_978( .ZN(N4724), .A(N4147) );
  INV_X1 NOT1_979( .ZN(N4725), .A(N4144) );
  INV_X1 NOT1_980( .ZN(N4726), .A(N4159) );
  INV_X1 NOT1_981( .ZN(N4727), .A(N4156) );
  INV_X1 NOT1_982( .ZN(N4728), .A(N4153) );
  INV_X1 NOT1_983( .ZN(N4729), .A(N4097) );
  INV_X4 NOT1_984( .ZN(N4730), .A(N4094) );
  INV_X1 NOT1_985( .ZN(N4731), .A(N4091) );
  INV_X1 NOT1_986( .ZN(N4732), .A(N4088) );
  INV_X1 NOT1_987( .ZN(N4733), .A(N4109) );
  INV_X1 NOT1_988( .ZN(N4734), .A(N4106) );
  INV_X1 NOT1_989( .ZN(N4735), .A(N4103) );
  INV_X1 NOT1_990( .ZN(N4736), .A(N4100) );
  AND2_X1 AND2_991( .ZN(N4737), .A1(N4273), .A2(N2877) );
  AND2_X1 AND2_992( .ZN(N4738), .A1(N4274), .A2(N2877) );
  AND2_X1 AND2_993( .ZN(N4739), .A1(N4276), .A2(N2877) );
  AND2_X1 AND2_994( .ZN(N4740), .A1(N4277), .A2(N2877) );
  AND3_X1 AND3_995( .ZN(N4741), .A1(N4150), .A2(N1758), .A3(N1755) );
  INV_X1 NOT1_996( .ZN(N4855), .A(N4212) );
  NAND2_X1 NAND2_997( .ZN(N4856), .A1(N4212), .A2(N2712) );
  NAND2_X1 NAND2_998( .ZN(N4908), .A1(N4215), .A2(N2718) );
  INV_X1 NOT1_999( .ZN(N4909), .A(N4215) );
  AND2_X1 AND2_1000( .ZN(N4939), .A1(N4515), .A2(N4185) );
  AND2_X1 AND2_1001( .ZN(N4942), .A1(N4516), .A2(N4186) );
  INV_X1 NOT1_1002( .ZN(N4947), .A(N4219) );
  AND3_X1 AND3_1003( .ZN(N4953), .A1(N4188), .A2(N3775), .A3(N3779) );
  AND3_X1 AND3_1004( .ZN(N4954), .A1(N3771), .A2(N4191), .A3(N3780) );
  AND3_X1 AND3_1005( .ZN(N4955), .A1(N4191), .A2(N4188), .A3(N3038) );
  AND3_X2 AND3_1006( .ZN(N4956), .A1(N4109), .A2(N3097), .A3(N3108) );
  AND3_X1 AND3_1007( .ZN(N4957), .A1(N4106), .A2(N3097), .A3(N3108) );
  AND3_X1 AND3_1008( .ZN(N4958), .A1(N4103), .A2(N3097), .A3(N3108) );
  AND3_X1 AND3_1009( .ZN(N4959), .A1(N4100), .A2(N3097), .A3(N3108) );
  AND3_X1 AND3_1010( .ZN(N4960), .A1(N4159), .A2(N3119), .A3(N3130) );
  AND3_X1 AND3_1011( .ZN(N4961), .A1(N4156), .A2(N3119), .A3(N3130) );
  INV_X1 NOT1_1012( .ZN(N4965), .A(N4225) );
  INV_X1 NOT1_1013( .ZN(N4966), .A(N4228) );
  INV_X1 NOT1_1014( .ZN(N4967), .A(N4231) );
  INV_X1 NOT1_1015( .ZN(N4968), .A(N4234) );
  INV_X1 NOT1_1016( .ZN(N4972), .A(N4246) );
  INV_X1 NOT1_1017( .ZN(N4973), .A(N4249) );
  INV_X1 NOT1_1018( .ZN(N4974), .A(N4252) );
  NAND2_X1 NAND2_1019( .ZN(N4975), .A1(N4252), .A2(N4199) );
  INV_X1 NOT1_1020( .ZN(N4976), .A(N4206) );
  INV_X4 NOT1_1021( .ZN(N4977), .A(N4209) );
  AND3_X1 AND3_1022( .ZN(N4978), .A1(N3793), .A2(N3789), .A3(N4206) );
  AND3_X1 AND3_1023( .ZN(N4979), .A1(N4203), .A2(N4200), .A3(N4209) );
  AND3_X1 AND3_1024( .ZN(N4980), .A1(N4097), .A2(N3147), .A3(N3158) );
  AND3_X1 AND3_1025( .ZN(N4981), .A1(N4094), .A2(N3147), .A3(N3158) );
  AND3_X1 AND3_1026( .ZN(N4982), .A1(N4091), .A2(N3147), .A3(N3158) );
  AND3_X1 AND3_1027( .ZN(N4983), .A1(N4088), .A2(N3147), .A3(N3158) );
  AND3_X1 AND3_1028( .ZN(N4984), .A1(N4153), .A2(N3169), .A3(N3180) );
  AND3_X1 AND3_1029( .ZN(N4985), .A1(N4147), .A2(N3169), .A3(N3180) );
  AND3_X1 AND3_1030( .ZN(N4986), .A1(N4144), .A2(N3169), .A3(N3180) );
  AND3_X1 AND3_1031( .ZN(N4987), .A1(N4150), .A2(N3169), .A3(N3180) );
  NAND2_X1 NAND2_1032( .ZN(N5049), .A1(N4701), .A2(N4702) );
  INV_X1 NOT1_1033( .ZN(N5052), .A(N4237) );
  INV_X1 NOT1_1034( .ZN(N5053), .A(N4240) );
  INV_X1 NOT1_1035( .ZN(N5054), .A(N4243) );
  INV_X1 NOT1_1036( .ZN(N5055), .A(N4255) );
  INV_X1 NOT1_1037( .ZN(N5056), .A(N4258) );
  NAND2_X1 NAND2_1038( .ZN(N5057), .A1(N3819), .A2(N4720) );
  INV_X1 NOT1_1039( .ZN(N5058), .A(N4264) );
  NAND2_X1 NAND2_1040( .ZN(N5059), .A1(N4264), .A2(N4267) );
  AND4_X1 AND4_1041( .ZN(N5060), .A1(N4724), .A2(N4725), .A3(N4269), .A4(N4027) );
  AND4_X1 AND4_1042( .ZN(N5061), .A1(N4726), .A2(N4727), .A3(N3827), .A4(N4728) );
  AND4_X1 AND4_1043( .ZN(N5062), .A1(N4729), .A2(N4730), .A3(N4731), .A4(N4732) );
  AND4_X1 AND4_1044( .ZN(N5063), .A1(N4733), .A2(N4734), .A3(N4735), .A4(N4736) );
  AND2_X1 AND2_1045( .ZN(N5065), .A1(N4357), .A2(N4375) );
  AND3_X1 AND3_1046( .ZN(N5066), .A1(N4364), .A2(N4357), .A3(N4379) );
  AND2_X1 AND2_1047( .ZN(N5067), .A1(N4418), .A2(N4436) );
  AND3_X1 AND3_1048( .ZN(N5068), .A1(N4425), .A2(N4418), .A3(N4440) );
  INV_X1 NOT1_1049( .ZN(N5069), .A(N4548) );
  NAND2_X1 NAND2_1050( .ZN(N5070), .A1(N4548), .A2(N2628) );
  INV_X1 NOT1_1051( .ZN(N5071), .A(N4551) );
  NAND2_X1 NAND2_1052( .ZN(N5072), .A1(N4551), .A2(N2629) );
  INV_X1 NOT1_1053( .ZN(N5073), .A(N4554) );
  NAND2_X1 NAND2_1054( .ZN(N5074), .A1(N4554), .A2(N2630) );
  INV_X1 NOT1_1055( .ZN(N5075), .A(N4557) );
  NAND2_X1 NAND2_1056( .ZN(N5076), .A1(N4557), .A2(N2631) );
  INV_X1 NOT1_1057( .ZN(N5077), .A(N4560) );
  NAND2_X1 NAND2_1058( .ZN(N5078), .A1(N4560), .A2(N2632) );
  INV_X1 NOT1_1059( .ZN(N5079), .A(N4563) );
  NAND2_X1 NAND2_1060( .ZN(N5080), .A1(N4563), .A2(N2633) );
  INV_X1 NOT1_1061( .ZN(N5081), .A(N4566) );
  NAND2_X1 NAND2_1062( .ZN(N5082), .A1(N4566), .A2(N2634) );
  INV_X1 NOT1_1063( .ZN(N5083), .A(N4569) );
  NAND2_X1 NAND2_1064( .ZN(N5084), .A1(N4569), .A2(N2635) );
  INV_X1 NOT1_1065( .ZN(N5085), .A(N4572) );
  NAND2_X1 NAND2_1066( .ZN(N5086), .A1(N4572), .A2(N2636) );
  INV_X1 NOT1_1067( .ZN(N5087), .A(N4575) );
  NAND2_X1 NAND2_1068( .ZN(N5088), .A1(N4578), .A2(N2638) );
  INV_X1 NOT1_1069( .ZN(N5089), .A(N4578) );
  NAND2_X1 NAND2_1070( .ZN(N5090), .A1(N4581), .A2(N2639) );
  INV_X1 NOT1_1071( .ZN(N5091), .A(N4581) );
  NAND2_X1 NAND2_1072( .ZN(N5092), .A1(N4584), .A2(N2640) );
  INV_X1 NOT1_1073( .ZN(N5093), .A(N4584) );
  NAND2_X1 NAND2_1074( .ZN(N5094), .A1(N4587), .A2(N2641) );
  INV_X1 NOT1_1075( .ZN(N5095), .A(N4587) );
  NAND2_X1 NAND2_1076( .ZN(N5096), .A1(N4590), .A2(N2642) );
  INV_X1 NOT1_1077( .ZN(N5097), .A(N4590) );
  NAND2_X1 NAND2_1078( .ZN(N5098), .A1(N4593), .A2(N2643) );
  INV_X1 NOT1_1079( .ZN(N5099), .A(N4593) );
  NAND2_X1 NAND2_1080( .ZN(N5100), .A1(N4596), .A2(N2644) );
  INV_X1 NOT1_1081( .ZN(N5101), .A(N4596) );
  NAND2_X1 NAND2_1082( .ZN(N5102), .A1(N4599), .A2(N2645) );
  INV_X1 NOT1_1083( .ZN(N5103), .A(N4599) );
  NAND2_X1 NAND2_1084( .ZN(N5104), .A1(N4602), .A2(N2646) );
  INV_X2 NOT1_1085( .ZN(N5105), .A(N4602) );
  INV_X1 NOT1_1086( .ZN(N5106), .A(N4611) );
  NAND2_X1 NAND2_1087( .ZN(N5107), .A1(N4611), .A2(N2709) );
  INV_X1 NOT1_1088( .ZN(N5108), .A(N4614) );
  NAND2_X1 NAND2_1089( .ZN(N5109), .A1(N4614), .A2(N2710) );
  INV_X1 NOT1_1090( .ZN(N5110), .A(N4617) );
  NAND2_X1 NAND2_1091( .ZN(N5111), .A1(N4617), .A2(N2711) );
  NAND2_X1 NAND2_1092( .ZN(N5112), .A1(N1890), .A2(N4855) );
  INV_X1 NOT1_1093( .ZN(N5113), .A(N4621) );
  NAND2_X1 NAND2_1094( .ZN(N5114), .A1(N4621), .A2(N2713) );
  INV_X1 NOT1_1095( .ZN(N5115), .A(N4624) );
  NAND2_X1 NAND2_1096( .ZN(N5116), .A1(N4624), .A2(N2714) );
  AND2_X1 AND2_1097( .ZN(N5117), .A1(N4364), .A2(N4379) );
  AND2_X1 AND2_1098( .ZN(N5118), .A1(N4364), .A2(N4379) );
  AND2_X1 AND2_1099( .ZN(N5119), .A1(N54), .A2(N4405) );
  INV_X1 NOT1_1100( .ZN(N5120), .A(N4627) );
  NAND2_X1 NAND2_1101( .ZN(N5121), .A1(N4630), .A2(N2716) );
  INV_X1 NOT1_1102( .ZN(N5122), .A(N4630) );
  NAND2_X1 NAND2_1103( .ZN(N5123), .A1(N4633), .A2(N2717) );
  INV_X1 NOT1_1104( .ZN(N5124), .A(N4633) );
  NAND2_X1 NAND2_1105( .ZN(N5125), .A1(N1908), .A2(N4909) );
  NAND2_X1 NAND2_1106( .ZN(N5126), .A1(N4637), .A2(N2719) );
  INV_X1 NOT1_1107( .ZN(N5127), .A(N4637) );
  NAND2_X2 NAND2_1108( .ZN(N5128), .A1(N4640), .A2(N2720) );
  INV_X1 NOT1_1109( .ZN(N5129), .A(N4640) );
  NAND2_X1 NAND2_1110( .ZN(N5130), .A1(N4643), .A2(N2721) );
  INV_X1 NOT1_1111( .ZN(N5131), .A(N4643) );
  AND2_X1 AND2_1112( .ZN(N5132), .A1(N4425), .A2(N4440) );
  AND2_X1 AND2_1113( .ZN(N5133), .A1(N4425), .A2(N4440) );
  INV_X1 NOT1_1114( .ZN(N5135), .A(N4649) );
  INV_X1 NOT1_1115( .ZN(N5136), .A(N4652) );
  NAND2_X1 NAND2_1116( .ZN(N5137), .A1(N4655), .A2(N4521) );
  INV_X1 NOT1_1117( .ZN(N5138), .A(N4655) );
  INV_X1 NOT1_1118( .ZN(N5139), .A(N4658) );
  NAND2_X2 NAND2_1119( .ZN(N5140), .A1(N4658), .A2(N4947) );
  INV_X1 NOT1_1120( .ZN(N5141), .A(N4674) );
  INV_X1 NOT1_1121( .ZN(N5142), .A(N4677) );
  INV_X1 NOT1_1122( .ZN(N5143), .A(N4680) );
  INV_X1 NOT1_1123( .ZN(N5144), .A(N4683) );
  NAND2_X1 NAND2_1124( .ZN(N5145), .A1(N4686), .A2(N4523) );
  INV_X1 NOT1_1125( .ZN(N5146), .A(N4686) );
  NOR2_X1 NOR2_1126( .ZN(N5147), .A1(N4953), .A2(N4196) );
  NOR2_X1 NOR2_1127( .ZN(N5148), .A1(N4954), .A2(N4955) );
  INV_X1 NOT1_1128( .ZN(N5150), .A(N4524) );
  NAND2_X1 NAND2_1129( .ZN(N5153), .A1(N4228), .A2(N4965) );
  NAND2_X1 NAND2_1130( .ZN(N5154), .A1(N4225), .A2(N4966) );
  NAND2_X1 NAND2_1131( .ZN(N5155), .A1(N4234), .A2(N4967) );
  NAND2_X1 NAND2_1132( .ZN(N5156), .A1(N4231), .A2(N4968) );
  INV_X1 NOT1_1133( .ZN(N5157), .A(N4532) );
  NAND2_X1 NAND2_1134( .ZN(N5160), .A1(N4249), .A2(N4972) );
  NAND2_X1 NAND2_1135( .ZN(N5161), .A1(N4246), .A2(N4973) );
  NAND2_X1 NAND2_1136( .ZN(N5162), .A1(N3816), .A2(N4974) );
  AND3_X1 AND3_1137( .ZN(N5163), .A1(N4200), .A2(N3793), .A3(N4976) );
  AND3_X1 AND3_1138( .ZN(N5164), .A1(N3789), .A2(N4203), .A3(N4977) );
  AND3_X1 AND3_1139( .ZN(N5165), .A1(N4942), .A2(N3147), .A3(N3158) );
  INV_X1 NOT1_1140( .ZN(N5166), .A(N4512) );
  BUF_X1 BUFF1_1141( .Z(N5169), .A(N4290) );
  INV_X1 NOT1_1142( .ZN(N5172), .A(N4605) );
  BUF_X1 BUFF1_1143( .Z(N5173), .A(N4325) );
  INV_X1 NOT1_1144( .ZN(N5176), .A(N4608) );
  BUF_X1 BUFF1_1145( .Z(N5177), .A(N4349) );
  BUF_X1 BUFF1_1146( .Z(N5180), .A(N4405) );
  BUF_X1 BUFF1_1147( .Z(N5183), .A(N4357) );
  BUF_X1 BUFF1_1148( .Z(N5186), .A(N4357) );
  BUF_X1 BUFF1_1149( .Z(N5189), .A(N4364) );
  BUF_X1 BUFF1_1150( .Z(N5192), .A(N4364) );
  BUF_X1 BUFF1_1151( .Z(N5195), .A(N4385) );
  INV_X1 NOT1_1152( .ZN(N5198), .A(N4646) );
  BUF_X1 BUFF1_1153( .Z(N5199), .A(N4418) );
  BUF_X1 BUFF1_1154( .Z(N5202), .A(N4425) );
  BUF_X1 BUFF1_1155( .Z(N5205), .A(N4445) );
  BUF_X1 BUFF1_1156( .Z(N5208), .A(N4418) );
  BUF_X1 BUFF1_1157( .Z(N5211), .A(N4425) );
  BUF_X1 BUFF1_1158( .Z(N5214), .A(N4477) );
  BUF_X1 BUFF1_1159( .Z(N5217), .A(N4469) );
  BUF_X1 BUFF1_1160( .Z(N5220), .A(N4477) );
  INV_X1 NOT1_1161( .ZN(N5223), .A(N4662) );
  INV_X1 NOT1_1162( .ZN(N5224), .A(N4665) );
  INV_X1 NOT1_1163( .ZN(N5225), .A(N4668) );
  INV_X1 NOT1_1164( .ZN(N5226), .A(N4671) );
  INV_X1 NOT1_1165( .ZN(N5227), .A(N4689) );
  INV_X1 NOT1_1166( .ZN(N5228), .A(N4692) );
  INV_X1 NOT1_1167( .ZN(N5229), .A(N4695) );
  INV_X1 NOT1_1168( .ZN(N5230), .A(N4698) );
  NAND2_X1 NAND2_1169( .ZN(N5232), .A1(N4240), .A2(N5052) );
  NAND2_X1 NAND2_1170( .ZN(N5233), .A1(N4237), .A2(N5053) );
  NAND2_X1 NAND2_1171( .ZN(N5234), .A1(N4258), .A2(N5055) );
  NAND2_X1 NAND2_1172( .ZN(N5235), .A1(N4255), .A2(N5056) );
  NAND2_X1 NAND2_1173( .ZN(N5236), .A1(N4721), .A2(N5057) );
  NAND2_X1 NAND2_1174( .ZN(N5239), .A1(N3824), .A2(N5058) );
  AND3_X1 AND3_1175( .ZN(N5240), .A1(N5060), .A2(N5061), .A3(N4270) );
  INV_X1 NOT1_1176( .ZN(N5241), .A(N4939) );
  NAND2_X1 NAND2_1177( .ZN(N5242), .A1(N1824), .A2(N5069) );
  NAND2_X1 NAND2_1178( .ZN(N5243), .A1(N1827), .A2(N5071) );
  NAND2_X1 NAND2_1179( .ZN(N5244), .A1(N1830), .A2(N5073) );
  NAND2_X1 NAND2_1180( .ZN(N5245), .A1(N1833), .A2(N5075) );
  NAND2_X1 NAND2_1181( .ZN(N5246), .A1(N1836), .A2(N5077) );
  NAND2_X1 NAND2_1182( .ZN(N5247), .A1(N1839), .A2(N5079) );
  NAND2_X1 NAND2_1183( .ZN(N5248), .A1(N1842), .A2(N5081) );
  NAND2_X1 NAND2_1184( .ZN(N5249), .A1(N1845), .A2(N5083) );
  NAND2_X1 NAND2_1185( .ZN(N5250), .A1(N1848), .A2(N5085) );
  NAND2_X2 NAND2_1186( .ZN(N5252), .A1(N1854), .A2(N5089) );
  NAND2_X2 NAND2_1187( .ZN(N5253), .A1(N1857), .A2(N5091) );
  NAND2_X2 NAND2_1188( .ZN(N5254), .A1(N1860), .A2(N5093) );
  NAND2_X2 NAND2_1189( .ZN(N5255), .A1(N1863), .A2(N5095) );
  NAND2_X2 NAND2_1190( .ZN(N5256), .A1(N1866), .A2(N5097) );
  NAND2_X2 NAND2_1191( .ZN(N5257), .A1(N1869), .A2(N5099) );
  NAND2_X2 NAND2_1192( .ZN(N5258), .A1(N1872), .A2(N5101) );
  NAND2_X1 NAND2_1193( .ZN(N5259), .A1(N1875), .A2(N5103) );
  NAND2_X1 NAND2_1194( .ZN(N5260), .A1(N1878), .A2(N5105) );
  NAND2_X1 NAND2_1195( .ZN(N5261), .A1(N1881), .A2(N5106) );
  NAND2_X1 NAND2_1196( .ZN(N5262), .A1(N1884), .A2(N5108) );
  NAND2_X1 NAND2_1197( .ZN(N5263), .A1(N1887), .A2(N5110) );
  NAND2_X1 NAND2_1198( .ZN(N5264), .A1(N5112), .A2(N4856) );
  NAND2_X1 NAND2_1199( .ZN(N5274), .A1(N1893), .A2(N5113) );
  NAND2_X1 NAND2_1200( .ZN(N5275), .A1(N1896), .A2(N5115) );
  NAND2_X1 NAND2_1201( .ZN(N5282), .A1(N1902), .A2(N5122) );
  NAND2_X1 NAND2_1202( .ZN(N5283), .A1(N1905), .A2(N5124) );
  NAND2_X1 NAND2_1203( .ZN(N5284), .A1(N4908), .A2(N5125) );
  NAND2_X1 NAND2_1204( .ZN(N5298), .A1(N1911), .A2(N5127) );
  NAND2_X1 NAND2_1205( .ZN(N5299), .A1(N1914), .A2(N5129) );
  NAND2_X1 NAND2_1206( .ZN(N5300), .A1(N1917), .A2(N5131) );
  NAND2_X1 NAND2_1207( .ZN(N5303), .A1(N4652), .A2(N5135) );
  NAND2_X1 NAND2_1208( .ZN(N5304), .A1(N4649), .A2(N5136) );
  NAND2_X1 NAND2_1209( .ZN(N5305), .A1(N4008), .A2(N5138) );
  NAND2_X1 NAND2_1210( .ZN(N5306), .A1(N4219), .A2(N5139) );
  NAND2_X1 NAND2_1211( .ZN(N5307), .A1(N4677), .A2(N5141) );
  NAND2_X1 NAND2_1212( .ZN(N5308), .A1(N4674), .A2(N5142) );
  NAND2_X1 NAND2_1213( .ZN(N5309), .A1(N4683), .A2(N5143) );
  NAND2_X1 NAND2_1214( .ZN(N5310), .A1(N4680), .A2(N5144) );
  NAND2_X1 NAND2_1215( .ZN(N5311), .A1(N4011), .A2(N5146) );
  INV_X1 NOT1_1216( .ZN(N5312), .A(N5049) );
  NAND2_X1 NAND2_1217( .ZN(N5315), .A1(N5153), .A2(N5154) );
  NAND2_X1 NAND2_1218( .ZN(N5319), .A1(N5155), .A2(N5156) );
  NAND2_X1 NAND2_1219( .ZN(N5324), .A1(N5160), .A2(N5161) );
  NAND2_X1 NAND2_1220( .ZN(N5328), .A1(N5162), .A2(N4975) );
  NOR2_X1 NOR2_1221( .ZN(N5331), .A1(N5163), .A2(N4978) );
  NOR2_X1 NOR2_1222( .ZN(N5332), .A1(N5164), .A2(N4979) );
  OR2_X1 OR2_1223( .ZN(N5346), .A1(N4412), .A2(N5119) );
  NAND2_X1 NAND2_1224( .ZN(N5363), .A1(N4665), .A2(N5223) );
  NAND2_X1 NAND2_1225( .ZN(N5364), .A1(N4662), .A2(N5224) );
  NAND2_X1 NAND2_1226( .ZN(N5365), .A1(N4671), .A2(N5225) );
  NAND2_X1 NAND2_1227( .ZN(N5366), .A1(N4668), .A2(N5226) );
  NAND2_X1 NAND2_1228( .ZN(N5367), .A1(N4692), .A2(N5227) );
  NAND2_X1 NAND2_1229( .ZN(N5368), .A1(N4689), .A2(N5228) );
  NAND2_X1 NAND2_1230( .ZN(N5369), .A1(N4698), .A2(N5229) );
  NAND2_X1 NAND2_1231( .ZN(N5370), .A1(N4695), .A2(N5230) );
  NAND2_X1 NAND2_1232( .ZN(N5371), .A1(N5148), .A2(N5147) );
  BUF_X1 BUFF1_1233( .Z(N5374), .A(N4939) );
  NAND2_X1 NAND2_1234( .ZN(N5377), .A1(N5232), .A2(N5233) );
  NAND2_X1 NAND2_1235( .ZN(N5382), .A1(N5234), .A2(N5235) );
  NAND2_X1 NAND2_1236( .ZN(N5385), .A1(N5239), .A2(N5059) );
  AND3_X1 AND3_1237( .ZN(N5388), .A1(N5062), .A2(N5063), .A3(N5241) );
  NAND2_X1 NAND2_1238( .ZN(N5389), .A1(N5242), .A2(N5070) );
  NAND2_X1 NAND2_1239( .ZN(N5396), .A1(N5243), .A2(N5072) );
  NAND2_X1 NAND2_1240( .ZN(N5407), .A1(N5244), .A2(N5074) );
  NAND2_X1 NAND2_1241( .ZN(N5418), .A1(N5245), .A2(N5076) );
  NAND2_X1 NAND2_1242( .ZN(N5424), .A1(N5246), .A2(N5078) );
  NAND2_X1 NAND2_1243( .ZN(N5431), .A1(N5247), .A2(N5080) );
  NAND2_X1 NAND2_1244( .ZN(N5441), .A1(N5248), .A2(N5082) );
  NAND2_X1 NAND2_1245( .ZN(N5452), .A1(N5249), .A2(N5084) );
  NAND2_X1 NAND2_1246( .ZN(N5462), .A1(N5250), .A2(N5086) );
  INV_X4 NOT1_1247( .ZN(N5469), .A(N5169) );
  NAND2_X1 NAND2_1248( .ZN(N5470), .A1(N5088), .A2(N5252) );
  NAND2_X1 NAND2_1249( .ZN(N5477), .A1(N5090), .A2(N5253) );
  NAND2_X1 NAND2_1250( .ZN(N5488), .A1(N5092), .A2(N5254) );
  NAND2_X1 NAND2_1251( .ZN(N5498), .A1(N5094), .A2(N5255) );
  NAND2_X1 NAND2_1252( .ZN(N5506), .A1(N5096), .A2(N5256) );
  NAND2_X1 NAND2_1253( .ZN(N5520), .A1(N5098), .A2(N5257) );
  NAND2_X1 NAND2_1254( .ZN(N5536), .A1(N5100), .A2(N5258) );
  NAND2_X1 NAND2_1255( .ZN(N5549), .A1(N5102), .A2(N5259) );
  NAND2_X1 NAND2_1256( .ZN(N5555), .A1(N5104), .A2(N5260) );
  NAND2_X1 NAND2_1257( .ZN(N5562), .A1(N5261), .A2(N5107) );
  NAND2_X1 NAND2_1258( .ZN(N5573), .A1(N5262), .A2(N5109) );
  NAND2_X1 NAND2_1259( .ZN(N5579), .A1(N5263), .A2(N5111) );
  NAND2_X1 NAND2_1260( .ZN(N5595), .A1(N5274), .A2(N5114) );
  NAND2_X1 NAND2_1261( .ZN(N5606), .A1(N5275), .A2(N5116) );
  NAND2_X1 NAND2_1262( .ZN(N5616), .A1(N5180), .A2(N2715) );
  INV_X1 NOT1_1263( .ZN(N5617), .A(N5180) );
  INV_X1 NOT1_1264( .ZN(N5618), .A(N5183) );
  INV_X1 NOT1_1265( .ZN(N5619), .A(N5186) );
  INV_X1 NOT1_1266( .ZN(N5620), .A(N5189) );
  INV_X1 NOT1_1267( .ZN(N5621), .A(N5192) );
  INV_X1 NOT1_1268( .ZN(N5622), .A(N5195) );
  NAND2_X1 NAND2_1269( .ZN(N5624), .A1(N5121), .A2(N5282) );
  NAND2_X1 NAND2_1270( .ZN(N5634), .A1(N5123), .A2(N5283) );
  NAND2_X1 NAND2_1271( .ZN(N5655), .A1(N5126), .A2(N5298) );
  NAND2_X1 NAND2_1272( .ZN(N5671), .A1(N5128), .A2(N5299) );
  NAND2_X1 NAND2_1273( .ZN(N5684), .A1(N5130), .A2(N5300) );
  INV_X1 NOT1_1274( .ZN(N5690), .A(N5202) );
  INV_X1 NOT1_1275( .ZN(N5691), .A(N5211) );
  NAND2_X1 NAND2_1276( .ZN(N5692), .A1(N5303), .A2(N5304) );
  NAND2_X1 NAND2_1277( .ZN(N5696), .A1(N5137), .A2(N5305) );
  NAND2_X1 NAND2_1278( .ZN(N5700), .A1(N5306), .A2(N5140) );
  NAND2_X1 NAND2_1279( .ZN(N5703), .A1(N5307), .A2(N5308) );
  NAND2_X1 NAND2_1280( .ZN(N5707), .A1(N5309), .A2(N5310) );
  NAND2_X1 NAND2_1281( .ZN(N5711), .A1(N5145), .A2(N5311) );
  AND2_X1 AND2_1282( .ZN(N5726), .A1(N5166), .A2(N4512) );
  INV_X1 NOT1_1283( .ZN(N5727), .A(N5173) );
  INV_X1 NOT1_1284( .ZN(N5728), .A(N5177) );
  INV_X1 NOT1_1285( .ZN(N5730), .A(N5199) );
  INV_X1 NOT1_1286( .ZN(N5731), .A(N5205) );
  INV_X1 NOT1_1287( .ZN(N5732), .A(N5208) );
  INV_X1 NOT1_1288( .ZN(N5733), .A(N5214) );
  INV_X1 NOT1_1289( .ZN(N5734), .A(N5217) );
  INV_X1 NOT1_1290( .ZN(N5735), .A(N5220) );
  NAND2_X1 NAND2_1291( .ZN(N5736), .A1(N5365), .A2(N5366) );
  NAND2_X1 NAND2_1292( .ZN(N5739), .A1(N5363), .A2(N5364) );
  NAND2_X1 NAND2_1293( .ZN(N5742), .A1(N5369), .A2(N5370) );
  NAND2_X1 NAND2_1294( .ZN(N5745), .A1(N5367), .A2(N5368) );
  INV_X1 NOT1_1295( .ZN(N5755), .A(N5236) );
  NAND2_X1 NAND2_1296( .ZN(N5756), .A1(N5332), .A2(N5331) );
  AND2_X1 AND2_1297( .ZN(N5954), .A1(N5264), .A2(N4396) );
  NAND2_X1 NAND2_1298( .ZN(N5955), .A1(N1899), .A2(N5617) );
  INV_X1 NOT1_1299( .ZN(N5956), .A(N5346) );
  AND2_X1 AND2_1300( .ZN(N6005), .A1(N5284), .A2(N4456) );
  AND2_X1 AND2_1301( .ZN(N6006), .A1(N5284), .A2(N4456) );
  INV_X1 NOT1_1302( .ZN(N6023), .A(N5371) );
  NAND2_X1 NAND2_1303( .ZN(N6024), .A1(N5371), .A2(N5312) );
  INV_X1 NOT1_1304( .ZN(N6025), .A(N5315) );
  INV_X1 NOT1_1305( .ZN(N6028), .A(N5324) );
  BUF_X1 BUFF1_1306( .Z(N6031), .A(N5319) );
  BUF_X2 BUFF1_1307( .Z(N6034), .A(N5319) );
  BUF_X2 BUFF1_1308( .Z(N6037), .A(N5328) );
  BUF_X2 BUFF1_1309( .Z(N6040), .A(N5328) );
  INV_X1 NOT1_1310( .ZN(N6044), .A(N5385) );
  OR2_X1 OR2_1311( .ZN(N6045), .A1(N5166), .A2(N5726) );
  BUF_X1 BUFF1_1312( .Z(N6048), .A(N5264) );
  BUF_X1 BUFF1_1313( .Z(N6051), .A(N5284) );
  BUF_X1 BUFF1_1314( .Z(N6054), .A(N5284) );
  INV_X1 NOT1_1315( .ZN(N6065), .A(N5374) );
  NAND2_X1 NAND2_1316( .ZN(N6066), .A1(N5374), .A2(N5054) );
  INV_X1 NOT1_1317( .ZN(N6067), .A(N5377) );
  INV_X1 NOT1_1318( .ZN(N6068), .A(N5382) );
  NAND2_X1 NAND2_1319( .ZN(N6069), .A1(N5382), .A2(N5755) );
  AND2_X1 AND2_1320( .ZN(N6071), .A1(N5470), .A2(N4316) );
  AND3_X1 AND3_1321( .ZN(N6072), .A1(N5477), .A2(N5470), .A3(N4320) );
  AND4_X1 AND4_1322( .ZN(N6073), .A1(N5488), .A2(N5470), .A3(N4325), .A4(N5477) );
  AND4_X1 AND4_1323( .ZN(N6074), .A1(N5562), .A2(N4357), .A3(N4385), .A4(N4364) );
  AND2_X1 AND2_1324( .ZN(N6075), .A1(N5389), .A2(N4280) );
  AND3_X1 AND3_1325( .ZN(N6076), .A1(N5396), .A2(N5389), .A3(N4284) );
  AND4_X1 AND4_1326( .ZN(N6077), .A1(N5407), .A2(N5389), .A3(N4290), .A4(N5396) );
  AND4_X1 AND4_1327( .ZN(N6078), .A1(N5624), .A2(N4418), .A3(N4445), .A4(N4425) );
  INV_X1 NOT1_1328( .ZN(N6079), .A(N5418) );
  AND4_X1 AND4_1329( .ZN(N6080), .A1(N5396), .A2(N5418), .A3(N5407), .A4(N5389) );
  AND2_X1 AND2_1330( .ZN(N6083), .A1(N5396), .A2(N4284) );
  AND3_X1 AND3_1331( .ZN(N6084), .A1(N5407), .A2(N4290), .A3(N5396) );
  AND3_X1 AND3_1332( .ZN(N6085), .A1(N5418), .A2(N5407), .A3(N5396) );
  AND2_X1 AND2_1333( .ZN(N6086), .A1(N5396), .A2(N4284) );
  AND3_X1 AND3_1334( .ZN(N6087), .A1(N4290), .A2(N5407), .A3(N5396) );
  AND2_X1 AND2_1335( .ZN(N6088), .A1(N5407), .A2(N4290) );
  AND2_X1 AND2_1336( .ZN(N6089), .A1(N5418), .A2(N5407) );
  AND2_X1 AND2_1337( .ZN(N6090), .A1(N5407), .A2(N4290) );
  AND4_X1 AND5_1338_A( .ZN(extra0), .A1(N5431), .A2(N5462), .A3(N5441), .A4(N5424) );
  AND2_X1 AND5_1338( .ZN(N6091), .A1(extra0), .A2(N5452) );
  AND2_X1 AND2_1339( .ZN(N6094), .A1(N5424), .A2(N4298) );
  AND3_X1 AND3_1340( .ZN(N6095), .A1(N5431), .A2(N5424), .A3(N4301) );
  AND4_X1 AND4_1341( .ZN(N6096), .A1(N5441), .A2(N5424), .A3(N4305), .A4(N5431) );
  AND4_X1 AND5_1342_A( .ZN(extra1), .A1(N5452), .A2(N5441), .A3(N5424), .A4(N4310) );
  AND2_X1 AND5_1342( .ZN(N6097), .A1(extra1), .A2(N5431) );
  AND2_X1 AND2_1343( .ZN(N6098), .A1(N5431), .A2(N4301) );
  AND3_X1 AND3_1344( .ZN(N6099), .A1(N5441), .A2(N4305), .A3(N5431) );
  AND4_X1 AND4_1345( .ZN(N6100), .A1(N5452), .A2(N5441), .A3(N4310), .A4(N5431) );
  AND4_X1 AND5_1346_A( .ZN(extra2), .A1(N4), .A2(N5462), .A3(N5441), .A4(N5452) );
  AND2_X1 AND5_1346( .ZN(N6101), .A1(extra2), .A2(N5431) );
  AND2_X1 AND2_1347( .ZN(N6102), .A1(N4305), .A2(N5441) );
  AND3_X1 AND3_1348( .ZN(N6103), .A1(N5452), .A2(N5441), .A3(N4310) );
  AND4_X1 AND4_1349( .ZN(N6104), .A1(N4), .A2(N5462), .A3(N5441), .A4(N5452) );
  AND2_X1 AND2_1350( .ZN(N6105), .A1(N5452), .A2(N4310) );
  AND3_X1 AND3_1351( .ZN(N6106), .A1(N4), .A2(N5462), .A3(N5452) );
  AND2_X1 AND2_1352( .ZN(N6107), .A1(N4), .A2(N5462) );
  AND4_X1 AND4_1353( .ZN(N6108), .A1(N5549), .A2(N5488), .A3(N5477), .A4(N5470) );
  AND2_X1 AND2_1354( .ZN(N6111), .A1(N5477), .A2(N4320) );
  AND3_X1 AND3_1355( .ZN(N6112), .A1(N5488), .A2(N4325), .A3(N5477) );
  AND3_X1 AND3_1356( .ZN(N6113), .A1(N5549), .A2(N5488), .A3(N5477) );
  AND2_X1 AND2_1357( .ZN(N6114), .A1(N5477), .A2(N4320) );
  AND3_X1 AND3_1358( .ZN(N6115), .A1(N5488), .A2(N4325), .A3(N5477) );
  AND2_X1 AND2_1359( .ZN(N6116), .A1(N5488), .A2(N4325) );
  AND4_X1 AND5_1360_A( .ZN(extra3), .A1(N5555), .A2(N5536), .A3(N5520), .A4(N5506) );
  AND2_X1 AND5_1360( .ZN(N6117), .A1(extra3), .A2(N5498) );
  AND2_X1 AND2_1361( .ZN(N6120), .A1(N5498), .A2(N4332) );
  AND3_X1 AND3_1362( .ZN(N6121), .A1(N5506), .A2(N5498), .A3(N4336) );
  AND4_X1 AND4_1363( .ZN(N6122), .A1(N5520), .A2(N5498), .A3(N4342), .A4(N5506) );
  AND4_X1 AND5_1364_A( .ZN(extra4), .A1(N5536), .A2(N5520), .A3(N5498), .A4(N4349) );
  AND2_X1 AND5_1364( .ZN(N6123), .A1(extra4), .A2(N5506) );
  AND2_X1 AND2_1365( .ZN(N6124), .A1(N5506), .A2(N4336) );
  AND3_X1 AND3_1366( .ZN(N6125), .A1(N5520), .A2(N4342), .A3(N5506) );
  AND4_X1 AND4_1367( .ZN(N6126), .A1(N5536), .A2(N5520), .A3(N4349), .A4(N5506) );
  AND4_X1 AND4_1368( .ZN(N6127), .A1(N5555), .A2(N5520), .A3(N5506), .A4(N5536) );
  AND2_X1 AND2_1369( .ZN(N6128), .A1(N5506), .A2(N4336) );
  AND3_X1 AND3_1370( .ZN(N6129), .A1(N5520), .A2(N4342), .A3(N5506) );
  AND4_X1 AND4_1371( .ZN(N6130), .A1(N5536), .A2(N5520), .A3(N4349), .A4(N5506) );
  AND2_X1 AND2_1372( .ZN(N6131), .A1(N5520), .A2(N4342) );
  AND3_X1 AND3_1373( .ZN(N6132), .A1(N5536), .A2(N5520), .A3(N4349) );
  AND3_X1 AND3_1374( .ZN(N6133), .A1(N5555), .A2(N5520), .A3(N5536) );
  AND2_X1 AND2_1375( .ZN(N6134), .A1(N5520), .A2(N4342) );
  AND3_X1 AND3_1376( .ZN(N6135), .A1(N5536), .A2(N5520), .A3(N4349) );
  AND2_X1 AND2_1377( .ZN(N6136), .A1(N5536), .A2(N4349) );
  AND2_X1 AND2_1378( .ZN(N6137), .A1(N5549), .A2(N5488) );
  AND2_X1 AND2_1379( .ZN(N6138), .A1(N5555), .A2(N5536) );
  INV_X1 NOT1_1380( .ZN(N6139), .A(N5573) );
  AND4_X1 AND4_1381( .ZN(N6140), .A1(N4364), .A2(N5573), .A3(N5562), .A4(N4357) );
  AND3_X1 AND3_1382( .ZN(N6143), .A1(N5562), .A2(N4385), .A3(N4364) );
  AND3_X1 AND3_1383( .ZN(N6144), .A1(N5573), .A2(N5562), .A3(N4364) );
  AND3_X1 AND3_1384( .ZN(N6145), .A1(N4385), .A2(N5562), .A3(N4364) );
  AND2_X1 AND2_1385( .ZN(N6146), .A1(N5562), .A2(N4385) );
  AND2_X1 AND2_1386( .ZN(N6147), .A1(N5573), .A2(N5562) );
  AND2_X1 AND2_1387( .ZN(N6148), .A1(N5562), .A2(N4385) );
  AND4_X1 AND5_1388_A( .ZN(extra5), .A1(N5264), .A2(N4405), .A3(N5595), .A4(N5579) );
  AND2_X2 AND5_1388( .ZN(N6149), .A1(extra5), .A2(N5606) );
  AND2_X2 AND2_1389( .ZN(N6152), .A1(N5579), .A2(N4067) );
  AND3_X2 AND3_1390( .ZN(N6153), .A1(N5264), .A2(N5579), .A3(N4396) );
  AND4_X1 AND4_1391( .ZN(N6154), .A1(N5595), .A2(N5579), .A3(N4400), .A4(N5264) );
  AND4_X1 AND5_1392_A( .ZN(extra6), .A1(N5606), .A2(N5595), .A3(N5579), .A4(N4412) );
  AND2_X1 AND5_1392( .ZN(N6155), .A1(extra6), .A2(N5264) );
  AND3_X1 AND3_1393( .ZN(N6156), .A1(N5595), .A2(N4400), .A3(N5264) );
  AND4_X1 AND4_1394( .ZN(N6157), .A1(N5606), .A2(N5595), .A3(N4412), .A4(N5264) );
  AND4_X1 AND5_1395_A( .ZN(extra7), .A1(N54), .A2(N4405), .A3(N5595), .A4(N5606) );
  AND2_X1 AND5_1395( .ZN(N6158), .A1(extra7), .A2(N5264) );
  AND2_X1 AND2_1396( .ZN(N6159), .A1(N4400), .A2(N5595) );
  AND3_X1 AND3_1397( .ZN(N6160), .A1(N5606), .A2(N5595), .A3(N4412) );
  AND4_X1 AND4_1398( .ZN(N6161), .A1(N54), .A2(N4405), .A3(N5595), .A4(N5606) );
  AND2_X1 AND2_1399( .ZN(N6162), .A1(N5606), .A2(N4412) );
  AND3_X1 AND3_1400( .ZN(N6163), .A1(N54), .A2(N4405), .A3(N5606) );
  NAND2_X1 NAND2_1401( .ZN(N6164), .A1(N5616), .A2(N5955) );
  AND4_X1 AND4_1402( .ZN(N6168), .A1(N5684), .A2(N5624), .A3(N4425), .A4(N4418) );
  AND3_X1 AND3_1403( .ZN(N6171), .A1(N5624), .A2(N4445), .A3(N4425) );
  AND3_X1 AND3_1404( .ZN(N6172), .A1(N5684), .A2(N5624), .A3(N4425) );
  AND3_X1 AND3_1405( .ZN(N6173), .A1(N5624), .A2(N4445), .A3(N4425) );
  AND2_X1 AND2_1406( .ZN(N6174), .A1(N5624), .A2(N4445) );
  AND4_X1 AND5_1407_A( .ZN(extra8), .A1(N4477), .A2(N5671), .A3(N5655), .A4(N5284) );
  AND2_X1 AND5_1407( .ZN(N6175), .A1(extra8), .A2(N5634) );
  AND2_X1 AND2_1408( .ZN(N6178), .A1(N5634), .A2(N4080) );
  AND3_X1 AND3_1409( .ZN(N6179), .A1(N5284), .A2(N5634), .A3(N4456) );
  AND4_X1 AND4_1410( .ZN(N6180), .A1(N5655), .A2(N5634), .A3(N4462), .A4(N5284) );
  AND4_X1 AND5_1411_A( .ZN(extra9), .A1(N5671), .A2(N5655), .A3(N5634), .A4(N4469) );
  AND2_X1 AND5_1411( .ZN(N6181), .A1(extra9), .A2(N5284) );
  AND3_X1 AND3_1412( .ZN(N6182), .A1(N5655), .A2(N4462), .A3(N5284) );
  AND4_X1 AND4_1413( .ZN(N6183), .A1(N5671), .A2(N5655), .A3(N4469), .A4(N5284) );
  AND4_X1 AND4_1414( .ZN(N6184), .A1(N4477), .A2(N5655), .A3(N5284), .A4(N5671) );
  AND3_X1 AND3_1415( .ZN(N6185), .A1(N5655), .A2(N4462), .A3(N5284) );
  AND4_X1 AND4_1416( .ZN(N6186), .A1(N5671), .A2(N5655), .A3(N4469), .A4(N5284) );
  AND2_X1 AND2_1417( .ZN(N6187), .A1(N5655), .A2(N4462) );
  AND3_X1 AND3_1418( .ZN(N6188), .A1(N5671), .A2(N5655), .A3(N4469) );
  AND3_X1 AND3_1419( .ZN(N6189), .A1(N4477), .A2(N5655), .A3(N5671) );
  AND2_X1 AND2_1420( .ZN(N6190), .A1(N5655), .A2(N4462) );
  AND3_X1 AND3_1421( .ZN(N6191), .A1(N5671), .A2(N5655), .A3(N4469) );
  AND2_X1 AND2_1422( .ZN(N6192), .A1(N5671), .A2(N4469) );
  AND2_X1 AND2_1423( .ZN(N6193), .A1(N5684), .A2(N5624) );
  AND2_X1 AND2_1424( .ZN(N6194), .A1(N4477), .A2(N5671) );
  INV_X1 NOT1_1425( .ZN(N6197), .A(N5692) );
  INV_X1 NOT1_1426( .ZN(N6200), .A(N5696) );
  INV_X1 NOT1_1427( .ZN(N6203), .A(N5703) );
  INV_X1 NOT1_1428( .ZN(N6206), .A(N5707) );
  BUF_X1 BUFF1_1429( .Z(N6209), .A(N5700) );
  BUF_X1 BUFF1_1430( .Z(N6212), .A(N5700) );
  BUF_X1 BUFF1_1431( .Z(N6215), .A(N5711) );
  BUF_X1 BUFF1_1432( .Z(N6218), .A(N5711) );
  NAND2_X1 NAND2_1433( .ZN(N6221), .A1(N5049), .A2(N6023) );
  INV_X1 NOT1_1434( .ZN(N6234), .A(N5756) );
  NAND2_X1 NAND2_1435( .ZN(N6235), .A1(N5756), .A2(N6044) );
  BUF_X1 BUFF1_1436( .Z(N6238), .A(N5462) );
  BUF_X1 BUFF1_1437( .Z(N6241), .A(N5389) );
  BUF_X1 BUFF1_1438( .Z(N6244), .A(N5389) );
  BUF_X1 BUFF1_1439( .Z(N6247), .A(N5396) );
  BUF_X1 BUFF1_1440( .Z(N6250), .A(N5396) );
  BUF_X1 BUFF1_1441( .Z(N6253), .A(N5407) );
  BUF_X1 BUFF1_1442( .Z(N6256), .A(N5407) );
  BUF_X1 BUFF1_1443( .Z(N6259), .A(N5424) );
  BUF_X1 BUFF1_1444( .Z(N6262), .A(N5431) );
  BUF_X1 BUFF1_1445( .Z(N6265), .A(N5441) );
  BUF_X1 BUFF1_1446( .Z(N6268), .A(N5452) );
  BUF_X1 BUFF1_1447( .Z(N6271), .A(N5549) );
  BUF_X1 BUFF1_1448( .Z(N6274), .A(N5488) );
  BUF_X1 BUFF1_1449( .Z(N6277), .A(N5470) );
  BUF_X1 BUFF1_1450( .Z(N6280), .A(N5477) );
  BUF_X4 BUFF1_1451( .Z(N6283), .A(N5549) );
  BUF_X4 BUFF1_1452( .Z(N6286), .A(N5488) );
  BUF_X4 BUFF1_1453( .Z(N6289), .A(N5470) );
  BUF_X4 BUFF1_1454( .Z(N6292), .A(N5477) );
  BUF_X1 BUFF1_1455( .Z(N6295), .A(N5555) );
  BUF_X1 BUFF1_1456( .Z(N6298), .A(N5536) );
  BUF_X1 BUFF1_1457( .Z(N6301), .A(N5498) );
  BUF_X1 BUFF1_1458( .Z(N6304), .A(N5520) );
  BUF_X1 BUFF1_1459( .Z(N6307), .A(N5506) );
  BUF_X1 BUFF1_1460( .Z(N6310), .A(N5506) );
  BUF_X1 BUFF1_1461( .Z(N6313), .A(N5555) );
  BUF_X1 BUFF1_1462( .Z(N6316), .A(N5536) );
  BUF_X1 BUFF1_1463( .Z(N6319), .A(N5498) );
  BUF_X1 BUFF1_1464( .Z(N6322), .A(N5520) );
  BUF_X1 BUFF1_1465( .Z(N6325), .A(N5562) );
  BUF_X1 BUFF1_1466( .Z(N6328), .A(N5562) );
  BUF_X1 BUFF1_1467( .Z(N6331), .A(N5579) );
  BUF_X1 BUFF1_1468( .Z(N6335), .A(N5595) );
  BUF_X1 BUFF1_1469( .Z(N6338), .A(N5606) );
  BUF_X1 BUFF1_1470( .Z(N6341), .A(N5684) );
  BUF_X1 BUFF1_1471( .Z(N6344), .A(N5624) );
  BUF_X1 BUFF1_1472( .Z(N6347), .A(N5684) );
  BUF_X1 BUFF1_1473( .Z(N6350), .A(N5624) );
  BUF_X1 BUFF1_1474( .Z(N6353), .A(N5671) );
  BUF_X8 BUFF1_1475( .Z(N6356), .A(N5634) );
  BUF_X8 BUFF1_1476( .Z(N6359), .A(N5655) );
  BUF_X1 BUFF1_1477( .Z(N6364), .A(N5671) );
  BUF_X1 BUFF1_1478( .Z(N6367), .A(N5634) );
  BUF_X1 BUFF1_1479( .Z(N6370), .A(N5655) );
  INV_X1 NOT1_1480( .ZN(N6373), .A(N5736) );
  INV_X1 NOT1_1481( .ZN(N6374), .A(N5739) );
  INV_X1 NOT1_1482( .ZN(N6375), .A(N5742) );
  INV_X1 NOT1_1483( .ZN(N6376), .A(N5745) );
  NAND2_X1 NAND2_1484( .ZN(N6377), .A1(N4243), .A2(N6065) );
  NAND2_X1 NAND2_1485( .ZN(N6378), .A1(N5236), .A2(N6068) );
  OR4_X1 OR4_1486( .ZN(N6382), .A1(N4268), .A2(N6071), .A3(N6072), .A4(N6073) );
  OR4_X1 OR4_1487( .ZN(N6386), .A1(N3968), .A2(N5065), .A3(N5066), .A4(N6074) );
  OR4_X1 OR4_1488( .ZN(N6388), .A1(N4271), .A2(N6075), .A3(N6076), .A4(N6077) );
  OR4_X1 OR4_1489( .ZN(N6392), .A1(N3968), .A2(N5067), .A3(N5068), .A4(N6078) );
  OR4_X1 OR5_1490_A( .ZN(extra10), .A1(N4297), .A2(N6094), .A3(N6095), .A4(N6096) );
  OR2_X1 OR5_1490( .ZN(N6397), .A1(extra10), .A2(N6097) );
  OR2_X1 OR2_1491( .ZN(N6411), .A1(N4320), .A2(N6116) );
  OR4_X2 OR5_1492_A( .ZN(extra11), .A1(N4331), .A2(N6120), .A3(N6121), .A4(N6122) );
  OR2_X2 OR5_1492( .ZN(N6415), .A1(extra11), .A2(N6123) );
  OR2_X1 OR2_1493( .ZN(N6419), .A1(N4342), .A2(N6136) );
  OR4_X1 OR5_1494_A( .ZN(extra12), .A1(N4392), .A2(N6152), .A3(N6153), .A4(N6154) );
  OR2_X1 OR5_1494( .ZN(N6427), .A1(extra12), .A2(N6155) );
  INV_X1 NOT1_1495( .ZN(N6434), .A(N6048) );
  OR2_X1 OR2_1496( .ZN(N6437), .A1(N4440), .A2(N6174) );
  OR4_X1 OR5_1497_A( .ZN(extra13), .A1(N4451), .A2(N6178), .A3(N6179), .A4(N6180) );
  OR2_X1 OR5_1497( .ZN(N6441), .A1(extra13), .A2(N6181) );
  OR2_X1 OR2_1498( .ZN(N6445), .A1(N4462), .A2(N6192) );
  INV_X1 NOT1_1499( .ZN(N6448), .A(N6051) );
  INV_X1 NOT1_1500( .ZN(N6449), .A(N6054) );
  NAND2_X1 NAND2_1501( .ZN(N6466), .A1(N6221), .A2(N6024) );
  INV_X1 NOT1_1502( .ZN(N6469), .A(N6031) );
  INV_X1 NOT1_1503( .ZN(N6470), .A(N6034) );
  INV_X1 NOT1_1504( .ZN(N6471), .A(N6037) );
  INV_X1 NOT1_1505( .ZN(N6472), .A(N6040) );
  AND3_X1 AND3_1506( .ZN(N6473), .A1(N5315), .A2(N4524), .A3(N6031) );
  AND3_X1 AND3_1507( .ZN(N6474), .A1(N6025), .A2(N5150), .A3(N6034) );
  AND3_X1 AND3_1508( .ZN(N6475), .A1(N5324), .A2(N4532), .A3(N6037) );
  AND3_X1 AND3_1509( .ZN(N6476), .A1(N6028), .A2(N5157), .A3(N6040) );
  NAND2_X1 NAND2_1510( .ZN(N6477), .A1(N5385), .A2(N6234) );
  NAND2_X1 NAND2_1511( .ZN(N6478), .A1(N6045), .A2(N132) );
  OR4_X1 OR4_1512( .ZN(N6482), .A1(N4280), .A2(N6083), .A3(N6084), .A4(N6085) );
  NOR3_X1 NOR3_1513( .ZN(N6486), .A1(N4280), .A2(N6086), .A3(N6087) );
  OR3_X1 OR3_1514( .ZN(N6490), .A1(N4284), .A2(N6088), .A3(N6089) );
  NOR2_X1 NOR2_1515( .ZN(N6494), .A1(N4284), .A2(N6090) );
  OR4_X1 OR5_1516_A( .ZN(extra14), .A1(N4298), .A2(N6098), .A3(N6099), .A4(N6100) );
  OR2_X1 OR5_1516( .ZN(N6500), .A1(extra14), .A2(N6101) );
  OR4_X1 OR4_1517( .ZN(N6504), .A1(N4301), .A2(N6102), .A3(N6103), .A4(N6104) );
  OR3_X1 OR3_1518( .ZN(N6508), .A1(N4305), .A2(N6105), .A3(N6106) );
  OR2_X1 OR2_1519( .ZN(N6512), .A1(N4310), .A2(N6107) );
  OR4_X1 OR4_1520( .ZN(N6516), .A1(N4316), .A2(N6111), .A3(N6112), .A4(N6113) );
  NOR3_X1 NOR3_1521( .ZN(N6526), .A1(N4316), .A2(N6114), .A3(N6115) );
  OR4_X1 OR4_1522( .ZN(N6536), .A1(N4336), .A2(N6131), .A3(N6132), .A4(N6133) );
  OR4_X1 OR5_1523_A( .ZN(extra15), .A1(N4332), .A2(N6124), .A3(N6125), .A4(N6126) );
  OR2_X1 OR5_1523( .ZN(N6539), .A1(extra15), .A2(N6127) );
  NOR3_X1 NOR3_1524( .ZN(N6553), .A1(N4336), .A2(N6134), .A3(N6135) );
  NOR3_X1 NOR4_1525_A( .ZN(extra16), .A1(N4332), .A2(N6128), .A3(N6129) );
  NOR2_X1 NOR4_1525( .ZN(N6556), .A1(extra16), .A2(N6130) );
  OR4_X1 OR4_1526( .ZN(N6566), .A1(N4375), .A2(N5117), .A3(N6143), .A4(N6144) );
  NOR3_X1 NOR3_1527( .ZN(N6569), .A1(N4375), .A2(N5118), .A3(N6145) );
  OR3_X1 OR3_1528( .ZN(N6572), .A1(N4379), .A2(N6146), .A3(N6147) );
  NOR2_X1 NOR2_1529( .ZN(N6575), .A1(N4379), .A2(N6148) );
  OR4_X1 OR5_1530_A( .ZN(extra17), .A1(N4067), .A2(N5954), .A3(N6156), .A4(N6157) );
  OR2_X1 OR5_1530( .ZN(N6580), .A1(extra17), .A2(N6158) );
  OR4_X1 OR4_1531( .ZN(N6584), .A1(N4396), .A2(N6159), .A3(N6160), .A4(N6161) );
  OR3_X1 OR3_1532( .ZN(N6587), .A1(N4400), .A2(N6162), .A3(N6163) );
  OR4_X1 OR4_1533( .ZN(N6592), .A1(N4436), .A2(N5132), .A3(N6171), .A4(N6172) );
  NOR3_X1 NOR3_1534( .ZN(N6599), .A1(N4436), .A2(N5133), .A3(N6173) );
  OR4_X1 OR4_1535( .ZN(N6606), .A1(N4456), .A2(N6187), .A3(N6188), .A4(N6189) );
  OR4_X1 OR5_1536_A( .ZN(extra18), .A1(N4080), .A2(N6005), .A3(N6182), .A4(N6183) );
  OR2_X1 OR5_1536( .ZN(N6609), .A1(extra18), .A2(N6184) );
  NOR3_X1 NOR3_1537( .ZN(N6619), .A1(N4456), .A2(N6190), .A3(N6191) );
  NOR3_X1 NOR4_1538_A( .ZN(extra19), .A1(N4080), .A2(N6006), .A3(N6185) );
  NOR2_X1 NOR4_1538( .ZN(N6622), .A1(extra19), .A2(N6186) );
  NAND2_X1 NAND2_1539( .ZN(N6630), .A1(N5739), .A2(N6373) );
  NAND2_X1 NAND2_1540( .ZN(N6631), .A1(N5736), .A2(N6374) );
  NAND2_X1 NAND2_1541( .ZN(N6632), .A1(N5745), .A2(N6375) );
  NAND2_X1 NAND2_1542( .ZN(N6633), .A1(N5742), .A2(N6376) );
  NAND2_X1 NAND2_1543( .ZN(N6634), .A1(N6377), .A2(N6066) );
  NAND2_X1 NAND2_1544( .ZN(N6637), .A1(N6069), .A2(N6378) );
  INV_X1 NOT1_1545( .ZN(N6640), .A(N6164) );
  AND2_X1 AND2_1546( .ZN(N6641), .A1(N6108), .A2(N6117) );
  AND2_X1 AND2_1547( .ZN(N6643), .A1(N6140), .A2(N6149) );
  AND2_X1 AND2_1548( .ZN(N6646), .A1(N6168), .A2(N6175) );
  AND2_X1 AND2_1549( .ZN(N6648), .A1(N6080), .A2(N6091) );
  NAND2_X1 NAND2_1550( .ZN(N6650), .A1(N6238), .A2(N2637) );
  INV_X1 NOT1_1551( .ZN(N6651), .A(N6238) );
  INV_X1 NOT1_1552( .ZN(N6653), .A(N6241) );
  INV_X1 NOT1_1553( .ZN(N6655), .A(N6244) );
  INV_X1 NOT1_1554( .ZN(N6657), .A(N6247) );
  INV_X1 NOT1_1555( .ZN(N6659), .A(N6250) );
  NAND2_X1 NAND2_1556( .ZN(N6660), .A1(N6253), .A2(N5087) );
  INV_X1 NOT1_1557( .ZN(N6661), .A(N6253) );
  NAND2_X1 NAND2_1558( .ZN(N6662), .A1(N6256), .A2(N5469) );
  INV_X1 NOT1_1559( .ZN(N6663), .A(N6256) );
  AND2_X1 AND2_1560( .ZN(N6664), .A1(N6091), .A2(N4) );
  INV_X1 NOT1_1561( .ZN(N6666), .A(N6259) );
  INV_X1 NOT1_1562( .ZN(N6668), .A(N6262) );
  INV_X1 NOT1_1563( .ZN(N6670), .A(N6265) );
  INV_X2 NOT1_1564( .ZN(N6672), .A(N6268) );
  INV_X2 NOT1_1565( .ZN(N6675), .A(N6117) );
  INV_X1 NOT1_1566( .ZN(N6680), .A(N6280) );
  INV_X1 NOT1_1567( .ZN(N6681), .A(N6292) );
  INV_X1 NOT1_1568( .ZN(N6682), .A(N6307) );
  INV_X1 NOT1_1569( .ZN(N6683), .A(N6310) );
  NAND2_X1 NAND2_1570( .ZN(N6689), .A1(N6325), .A2(N5120) );
  INV_X1 NOT1_1571( .ZN(N6690), .A(N6325) );
  NAND2_X1 NAND2_1572( .ZN(N6691), .A1(N6328), .A2(N5622) );
  INV_X1 NOT1_1573( .ZN(N6692), .A(N6328) );
  AND2_X1 AND2_1574( .ZN(N6693), .A1(N6149), .A2(N54) );
  INV_X1 NOT1_1575( .ZN(N6695), .A(N6331) );
  INV_X1 NOT1_1576( .ZN(N6698), .A(N6335) );
  NAND2_X1 NAND2_1577( .ZN(N6699), .A1(N6338), .A2(N5956) );
  INV_X1 NOT1_1578( .ZN(N6700), .A(N6338) );
  INV_X1 NOT1_1579( .ZN(N6703), .A(N6175) );
  INV_X1 NOT1_1580( .ZN(N6708), .A(N6209) );
  INV_X1 NOT1_1581( .ZN(N6709), .A(N6212) );
  INV_X1 NOT1_1582( .ZN(N6710), .A(N6215) );
  INV_X1 NOT1_1583( .ZN(N6711), .A(N6218) );
  AND3_X1 AND3_1584( .ZN(N6712), .A1(N5696), .A2(N5692), .A3(N6209) );
  AND3_X1 AND3_1585( .ZN(N6713), .A1(N6200), .A2(N6197), .A3(N6212) );
  AND3_X1 AND3_1586( .ZN(N6714), .A1(N5707), .A2(N5703), .A3(N6215) );
  AND3_X1 AND3_1587( .ZN(N6715), .A1(N6206), .A2(N6203), .A3(N6218) );
  BUF_X1 BUFF1_1588( .Z(N6716), .A(N6466) );
  AND3_X1 AND3_1589( .ZN(N6718), .A1(N6164), .A2(N1777), .A3(N3130) );
  AND3_X1 AND3_1590( .ZN(N6719), .A1(N5150), .A2(N5315), .A3(N6469) );
  AND3_X1 AND3_1591( .ZN(N6720), .A1(N4524), .A2(N6025), .A3(N6470) );
  AND3_X1 AND3_1592( .ZN(N6721), .A1(N5157), .A2(N5324), .A3(N6471) );
  AND3_X1 AND3_1593( .ZN(N6722), .A1(N4532), .A2(N6028), .A3(N6472) );
  NAND2_X1 NAND2_1594( .ZN(N6724), .A1(N6477), .A2(N6235) );
  INV_X1 NOT1_1595( .ZN(N6739), .A(N6271) );
  INV_X1 NOT1_1596( .ZN(N6740), .A(N6274) );
  INV_X1 NOT1_1597( .ZN(N6741), .A(N6277) );
  INV_X1 NOT1_1598( .ZN(N6744), .A(N6283) );
  INV_X1 NOT1_1599( .ZN(N6745), .A(N6286) );
  INV_X1 NOT1_1600( .ZN(N6746), .A(N6289) );
  INV_X1 NOT1_1601( .ZN(N6751), .A(N6295) );
  INV_X1 NOT1_1602( .ZN(N6752), .A(N6298) );
  INV_X1 NOT1_1603( .ZN(N6753), .A(N6301) );
  INV_X2 NOT1_1604( .ZN(N6754), .A(N6304) );
  INV_X2 NOT1_1605( .ZN(N6755), .A(N6322) );
  INV_X4 NOT1_1606( .ZN(N6760), .A(N6313) );
  INV_X4 NOT1_1607( .ZN(N6761), .A(N6316) );
  INV_X8 NOT1_1608( .ZN(N6762), .A(N6319) );
  INV_X1 NOT1_1609( .ZN(N6772), .A(N6341) );
  INV_X1 NOT1_1610( .ZN(N6773), .A(N6344) );
  INV_X1 NOT1_1611( .ZN(N6776), .A(N6347) );
  INV_X1 NOT1_1612( .ZN(N6777), .A(N6350) );
  INV_X1 NOT1_1613( .ZN(N6782), .A(N6353) );
  INV_X1 NOT1_1614( .ZN(N6783), .A(N6356) );
  INV_X1 NOT1_1615( .ZN(N6784), .A(N6359) );
  INV_X1 NOT1_1616( .ZN(N6785), .A(N6370) );
  INV_X1 NOT1_1617( .ZN(N6790), .A(N6364) );
  INV_X1 NOT1_1618( .ZN(N6791), .A(N6367) );
  NAND2_X1 NAND2_1619( .ZN(N6792), .A1(N6630), .A2(N6631) );
  NAND2_X1 NAND2_1620( .ZN(N6795), .A1(N6632), .A2(N6633) );
  AND2_X1 AND2_1621( .ZN(N6801), .A1(N6108), .A2(N6415) );
  AND2_X1 AND2_1622( .ZN(N6802), .A1(N6427), .A2(N6140) );
  AND2_X1 AND2_1623( .ZN(N6803), .A1(N6397), .A2(N6080) );
  AND2_X1 AND2_1624( .ZN(N6804), .A1(N6168), .A2(N6441) );
  INV_X1 NOT1_1625( .ZN(N6805), .A(N6466) );
  NAND2_X1 NAND2_1626( .ZN(N6806), .A1(N1851), .A2(N6651) );
  INV_X1 NOT1_1627( .ZN(N6807), .A(N6482) );
  NAND2_X1 NAND2_1628( .ZN(N6808), .A1(N6482), .A2(N6653) );
  INV_X1 NOT1_1629( .ZN(N6809), .A(N6486) );
  NAND2_X1 NAND2_1630( .ZN(N6810), .A1(N6486), .A2(N6655) );
  INV_X1 NOT1_1631( .ZN(N6811), .A(N6490) );
  NAND2_X1 NAND2_1632( .ZN(N6812), .A1(N6490), .A2(N6657) );
  INV_X1 NOT1_1633( .ZN(N6813), .A(N6494) );
  NAND2_X1 NAND2_1634( .ZN(N6814), .A1(N6494), .A2(N6659) );
  NAND2_X1 NAND2_1635( .ZN(N6815), .A1(N4575), .A2(N6661) );
  NAND2_X1 NAND2_1636( .ZN(N6816), .A1(N5169), .A2(N6663) );
  OR2_X1 OR2_1637( .ZN(N6817), .A1(N6397), .A2(N6664) );
  INV_X1 NOT1_1638( .ZN(N6823), .A(N6500) );
  NAND2_X1 NAND2_1639( .ZN(N6824), .A1(N6500), .A2(N6666) );
  INV_X1 NOT1_1640( .ZN(N6825), .A(N6504) );
  NAND2_X1 NAND2_1641( .ZN(N6826), .A1(N6504), .A2(N6668) );
  INV_X1 NOT1_1642( .ZN(N6827), .A(N6508) );
  NAND2_X1 NAND2_1643( .ZN(N6828), .A1(N6508), .A2(N6670) );
  INV_X1 NOT1_1644( .ZN(N6829), .A(N6512) );
  NAND2_X1 NAND2_1645( .ZN(N6830), .A1(N6512), .A2(N6672) );
  INV_X1 NOT1_1646( .ZN(N6831), .A(N6415) );
  INV_X1 NOT1_1647( .ZN(N6834), .A(N6566) );
  NAND2_X1 NAND2_1648( .ZN(N6835), .A1(N6566), .A2(N5618) );
  INV_X1 NOT1_1649( .ZN(N6836), .A(N6569) );
  NAND2_X1 NAND2_1650( .ZN(N6837), .A1(N6569), .A2(N5619) );
  INV_X1 NOT1_1651( .ZN(N6838), .A(N6572) );
  NAND2_X1 NAND2_1652( .ZN(N6839), .A1(N6572), .A2(N5620) );
  INV_X1 NOT1_1653( .ZN(N6840), .A(N6575) );
  NAND2_X1 NAND2_1654( .ZN(N6841), .A1(N6575), .A2(N5621) );
  NAND2_X1 NAND2_1655( .ZN(N6842), .A1(N4627), .A2(N6690) );
  NAND2_X1 NAND2_1656( .ZN(N6843), .A1(N5195), .A2(N6692) );
  OR2_X1 OR2_1657( .ZN(N6844), .A1(N6427), .A2(N6693) );
  INV_X1 NOT1_1658( .ZN(N6850), .A(N6580) );
  NAND2_X1 NAND2_1659( .ZN(N6851), .A1(N6580), .A2(N6695) );
  INV_X1 NOT1_1660( .ZN(N6852), .A(N6584) );
  NAND2_X1 NAND2_1661( .ZN(N6853), .A1(N6584), .A2(N6434) );
  INV_X1 NOT1_1662( .ZN(N6854), .A(N6587) );
  NAND2_X1 NAND2_1663( .ZN(N6855), .A1(N6587), .A2(N6698) );
  NAND2_X1 NAND2_1664( .ZN(N6856), .A1(N5346), .A2(N6700) );
  INV_X1 NOT1_1665( .ZN(N6857), .A(N6441) );
  AND3_X1 AND3_1666( .ZN(N6860), .A1(N6197), .A2(N5696), .A3(N6708) );
  AND3_X1 AND3_1667( .ZN(N6861), .A1(N5692), .A2(N6200), .A3(N6709) );
  AND3_X1 AND3_1668( .ZN(N6862), .A1(N6203), .A2(N5707), .A3(N6710) );
  AND3_X1 AND3_1669( .ZN(N6863), .A1(N5703), .A2(N6206), .A3(N6711) );
  OR3_X1 OR3_1670( .ZN(N6866), .A1(N4197), .A2(N6718), .A3(N3785) );
  NOR2_X1 NOR2_1671( .ZN(N6872), .A1(N6719), .A2(N6473) );
  NOR2_X1 NOR2_1672( .ZN(N6873), .A1(N6720), .A2(N6474) );
  NOR2_X1 NOR2_1673( .ZN(N6874), .A1(N6721), .A2(N6475) );
  NOR2_X1 NOR2_1674( .ZN(N6875), .A1(N6722), .A2(N6476) );
  INV_X1 NOT1_1675( .ZN(N6876), .A(N6637) );
  BUF_X1 BUFF1_1676( .Z(N6877), .A(N6724) );
  AND2_X1 AND2_1677( .ZN(N6879), .A1(N6045), .A2(N6478) );
  AND2_X1 AND2_1678( .ZN(N6880), .A1(N6478), .A2(N132) );
  OR2_X1 OR2_1679( .ZN(N6881), .A1(N6411), .A2(N6137) );
  INV_X1 NOT1_1680( .ZN(N6884), .A(N6516) );
  INV_X1 NOT1_1681( .ZN(N6885), .A(N6411) );
  INV_X1 NOT1_1682( .ZN(N6888), .A(N6526) );
  INV_X1 NOT1_1683( .ZN(N6889), .A(N6536) );
  NAND2_X1 NAND2_1684( .ZN(N6890), .A1(N6536), .A2(N5176) );
  OR2_X1 OR2_1685( .ZN(N6891), .A1(N6419), .A2(N6138) );
  INV_X1 NOT1_1686( .ZN(N6894), .A(N6539) );
  INV_X1 NOT1_1687( .ZN(N6895), .A(N6553) );
  NAND2_X1 NAND2_1688( .ZN(N6896), .A1(N6553), .A2(N5728) );
  INV_X1 NOT1_1689( .ZN(N6897), .A(N6419) );
  INV_X1 NOT1_1690( .ZN(N6900), .A(N6556) );
  OR2_X1 OR2_1691( .ZN(N6901), .A1(N6437), .A2(N6193) );
  INV_X1 NOT1_1692( .ZN(N6904), .A(N6592) );
  INV_X1 NOT1_1693( .ZN(N6905), .A(N6437) );
  INV_X1 NOT1_1694( .ZN(N6908), .A(N6599) );
  OR2_X1 OR2_1695( .ZN(N6909), .A1(N6445), .A2(N6194) );
  INV_X1 NOT1_1696( .ZN(N6912), .A(N6606) );
  INV_X1 NOT1_1697( .ZN(N6913), .A(N6609) );
  INV_X1 NOT1_1698( .ZN(N6914), .A(N6619) );
  NAND2_X1 NAND2_1699( .ZN(N6915), .A1(N6619), .A2(N5734) );
  INV_X1 NOT1_1700( .ZN(N6916), .A(N6445) );
  INV_X1 NOT1_1701( .ZN(N6919), .A(N6622) );
  INV_X1 NOT1_1702( .ZN(N6922), .A(N6634) );
  NAND2_X1 NAND2_1703( .ZN(N6923), .A1(N6634), .A2(N6067) );
  OR2_X1 OR2_1704( .ZN(N6924), .A1(N6382), .A2(N6801) );
  OR2_X1 OR2_1705( .ZN(N6925), .A1(N6386), .A2(N6802) );
  OR2_X1 OR2_1706( .ZN(N6926), .A1(N6388), .A2(N6803) );
  OR2_X1 OR2_1707( .ZN(N6927), .A1(N6392), .A2(N6804) );
  INV_X1 NOT1_1708( .ZN(N6930), .A(N6724) );
  NAND2_X1 NAND2_1709( .ZN(N6932), .A1(N6650), .A2(N6806) );
  NAND2_X1 NAND2_1710( .ZN(N6935), .A1(N6241), .A2(N6807) );
  NAND2_X1 NAND2_1711( .ZN(N6936), .A1(N6244), .A2(N6809) );
  NAND2_X1 NAND2_1712( .ZN(N6937), .A1(N6247), .A2(N6811) );
  NAND2_X1 NAND2_1713( .ZN(N6938), .A1(N6250), .A2(N6813) );
  NAND2_X1 NAND2_1714( .ZN(N6939), .A1(N6660), .A2(N6815) );
  NAND2_X1 NAND2_1715( .ZN(N6940), .A1(N6662), .A2(N6816) );
  NAND2_X1 NAND2_1716( .ZN(N6946), .A1(N6259), .A2(N6823) );
  NAND2_X1 NAND2_1717( .ZN(N6947), .A1(N6262), .A2(N6825) );
  NAND2_X1 NAND2_1718( .ZN(N6948), .A1(N6265), .A2(N6827) );
  NAND2_X2 NAND2_1719( .ZN(N6949), .A1(N6268), .A2(N6829) );
  NAND2_X2 NAND2_1720( .ZN(N6953), .A1(N5183), .A2(N6834) );
  NAND2_X2 NAND2_1721( .ZN(N6954), .A1(N5186), .A2(N6836) );
  NAND2_X2 NAND2_1722( .ZN(N6955), .A1(N5189), .A2(N6838) );
  NAND2_X2 NAND2_1723( .ZN(N6956), .A1(N5192), .A2(N6840) );
  NAND2_X1 NAND2_1724( .ZN(N6957), .A1(N6689), .A2(N6842) );
  NAND2_X1 NAND2_1725( .ZN(N6958), .A1(N6691), .A2(N6843) );
  NAND2_X1 NAND2_1726( .ZN(N6964), .A1(N6331), .A2(N6850) );
  NAND2_X1 NAND2_1727( .ZN(N6965), .A1(N6048), .A2(N6852) );
  NAND2_X1 NAND2_1728( .ZN(N6966), .A1(N6335), .A2(N6854) );
  NAND2_X1 NAND2_1729( .ZN(N6967), .A1(N6699), .A2(N6856) );
  NOR2_X1 NOR2_1730( .ZN(N6973), .A1(N6860), .A2(N6712) );
  NOR2_X1 NOR2_1731( .ZN(N6974), .A1(N6861), .A2(N6713) );
  NOR2_X1 NOR2_1732( .ZN(N6975), .A1(N6862), .A2(N6714) );
  NOR2_X1 NOR2_1733( .ZN(N6976), .A1(N6863), .A2(N6715) );
  INV_X1 NOT1_1734( .ZN(N6977), .A(N6792) );
  INV_X1 NOT1_1735( .ZN(N6978), .A(N6795) );
  OR2_X1 OR2_1736( .ZN(N6979), .A1(N6879), .A2(N6880) );
  NAND2_X1 NAND2_1737( .ZN(N6987), .A1(N4608), .A2(N6889) );
  NAND2_X1 NAND2_1738( .ZN(N6990), .A1(N5177), .A2(N6895) );
  NAND2_X1 NAND2_1739( .ZN(N6999), .A1(N5217), .A2(N6914) );
  NAND2_X1 NAND2_1740( .ZN(N7002), .A1(N5377), .A2(N6922) );
  NAND2_X1 NAND2_1741( .ZN(N7003), .A1(N6873), .A2(N6872) );
  NAND2_X1 NAND2_1742( .ZN(N7006), .A1(N6875), .A2(N6874) );
  AND3_X1 AND3_1743( .ZN(N7011), .A1(N6866), .A2(N2681), .A3(N2692) );
  AND3_X1 AND3_1744( .ZN(N7012), .A1(N6866), .A2(N2756), .A3(N2767) );
  AND3_X1 AND3_1745( .ZN(N7013), .A1(N6866), .A2(N2779), .A3(N2790) );
  INV_X1 NOT1_1746( .ZN(N7015), .A(N6866) );
  AND3_X1 AND3_1747( .ZN(N7016), .A1(N6866), .A2(N2801), .A3(N2812) );
  NAND2_X1 NAND2_1748( .ZN(N7018), .A1(N6935), .A2(N6808) );
  NAND2_X1 NAND2_1749( .ZN(N7019), .A1(N6936), .A2(N6810) );
  NAND2_X1 NAND2_1750( .ZN(N7020), .A1(N6937), .A2(N6812) );
  NAND2_X1 NAND2_1751( .ZN(N7021), .A1(N6938), .A2(N6814) );
  INV_X1 NOT1_1752( .ZN(N7022), .A(N6939) );
  INV_X1 NOT1_1753( .ZN(N7023), .A(N6817) );
  NAND2_X1 NAND2_1754( .ZN(N7028), .A1(N6946), .A2(N6824) );
  NAND2_X1 NAND2_1755( .ZN(N7031), .A1(N6947), .A2(N6826) );
  NAND2_X1 NAND2_1756( .ZN(N7034), .A1(N6948), .A2(N6828) );
  NAND2_X1 NAND2_1757( .ZN(N7037), .A1(N6949), .A2(N6830) );
  AND2_X1 AND2_1758( .ZN(N7040), .A1(N6817), .A2(N6079) );
  AND2_X1 AND2_1759( .ZN(N7041), .A1(N6831), .A2(N6675) );
  NAND2_X1 NAND2_1760( .ZN(N7044), .A1(N6953), .A2(N6835) );
  NAND2_X1 NAND2_1761( .ZN(N7045), .A1(N6954), .A2(N6837) );
  NAND2_X1 NAND2_1762( .ZN(N7046), .A1(N6955), .A2(N6839) );
  NAND2_X1 NAND2_1763( .ZN(N7047), .A1(N6956), .A2(N6841) );
  INV_X1 NOT1_1764( .ZN(N7048), .A(N6957) );
  INV_X1 NOT1_1765( .ZN(N7049), .A(N6844) );
  NAND2_X1 NAND2_1766( .ZN(N7054), .A1(N6964), .A2(N6851) );
  NAND2_X1 NAND2_1767( .ZN(N7057), .A1(N6965), .A2(N6853) );
  NAND2_X1 NAND2_1768( .ZN(N7060), .A1(N6966), .A2(N6855) );
  AND2_X1 AND2_1769( .ZN(N7064), .A1(N6844), .A2(N6139) );
  AND2_X1 AND2_1770( .ZN(N7065), .A1(N6857), .A2(N6703) );
  INV_X1 NOT1_1771( .ZN(N7072), .A(N6881) );
  NAND2_X1 NAND2_1772( .ZN(N7073), .A1(N6881), .A2(N5172) );
  INV_X1 NOT1_1773( .ZN(N7074), .A(N6885) );
  NAND2_X1 NAND2_1774( .ZN(N7075), .A1(N6885), .A2(N5727) );
  NAND2_X1 NAND2_1775( .ZN(N7076), .A1(N6890), .A2(N6987) );
  INV_X1 NOT1_1776( .ZN(N7079), .A(N6891) );
  NAND2_X1 NAND2_1777( .ZN(N7080), .A1(N6896), .A2(N6990) );
  INV_X1 NOT1_1778( .ZN(N7083), .A(N6897) );
  INV_X1 NOT1_1779( .ZN(N7084), .A(N6901) );
  NAND2_X1 NAND2_1780( .ZN(N7085), .A1(N6901), .A2(N5198) );
  INV_X1 NOT1_1781( .ZN(N7086), .A(N6905) );
  NAND2_X1 NAND2_1782( .ZN(N7087), .A1(N6905), .A2(N5731) );
  INV_X1 NOT1_1783( .ZN(N7088), .A(N6909) );
  NAND2_X1 NAND2_1784( .ZN(N7089), .A1(N6909), .A2(N6912) );
  NAND2_X1 NAND2_1785( .ZN(N7090), .A1(N6915), .A2(N6999) );
  INV_X1 NOT1_1786( .ZN(N7093), .A(N6916) );
  NAND2_X1 NAND2_1787( .ZN(N7094), .A1(N6974), .A2(N6973) );
  NAND2_X1 NAND2_1788( .ZN(N7097), .A1(N6976), .A2(N6975) );
  NAND2_X1 NAND2_1789( .ZN(N7101), .A1(N7002), .A2(N6923) );
  INV_X1 NOT1_1790( .ZN(N7105), .A(N6932) );
  INV_X1 NOT1_1791( .ZN(N7110), .A(N6967) );
  AND3_X1 AND3_1792( .ZN(N7114), .A1(N6979), .A2(N603), .A3(N1755) );
  INV_X1 NOT1_1793( .ZN(N7115), .A(N7019) );
  INV_X1 NOT1_1794( .ZN(N7116), .A(N7021) );
  AND2_X1 AND2_1795( .ZN(N7125), .A1(N6817), .A2(N7018) );
  AND2_X1 AND2_1796( .ZN(N7126), .A1(N6817), .A2(N7020) );
  AND2_X1 AND2_1797( .ZN(N7127), .A1(N6817), .A2(N7022) );
  INV_X1 NOT1_1798( .ZN(N7130), .A(N7045) );
  INV_X1 NOT1_1799( .ZN(N7131), .A(N7047) );
  AND2_X1 AND2_1800( .ZN(N7139), .A1(N6844), .A2(N7044) );
  AND2_X1 AND2_1801( .ZN(N7140), .A1(N6844), .A2(N7046) );
  AND2_X1 AND2_1802( .ZN(N7141), .A1(N6844), .A2(N7048) );
  AND3_X1 AND3_1803( .ZN(N7146), .A1(N6932), .A2(N1761), .A3(N3108) );
  AND3_X1 AND3_1804( .ZN(N7147), .A1(N6967), .A2(N1777), .A3(N3130) );
  INV_X1 NOT1_1805( .ZN(N7149), .A(N7003) );
  INV_X1 NOT1_1806( .ZN(N7150), .A(N7006) );
  NAND2_X1 NAND2_1807( .ZN(N7151), .A1(N7006), .A2(N6876) );
  NAND2_X1 NAND2_1808( .ZN(N7152), .A1(N4605), .A2(N7072) );
  NAND2_X1 NAND2_1809( .ZN(N7153), .A1(N5173), .A2(N7074) );
  NAND2_X1 NAND2_1810( .ZN(N7158), .A1(N4646), .A2(N7084) );
  NAND2_X1 NAND2_1811( .ZN(N7159), .A1(N5205), .A2(N7086) );
  NAND2_X1 NAND2_1812( .ZN(N7160), .A1(N6606), .A2(N7088) );
  INV_X1 NOT1_1813( .ZN(N7166), .A(N7037) );
  INV_X1 NOT1_1814( .ZN(N7167), .A(N7034) );
  INV_X1 NOT1_1815( .ZN(N7168), .A(N7031) );
  INV_X1 NOT1_1816( .ZN(N7169), .A(N7028) );
  INV_X1 NOT1_1817( .ZN(N7170), .A(N7060) );
  INV_X1 NOT1_1818( .ZN(N7171), .A(N7057) );
  INV_X1 NOT1_1819( .ZN(N7172), .A(N7054) );
  AND2_X1 AND2_1820( .ZN(N7173), .A1(N7115), .A2(N7023) );
  AND2_X2 AND2_1821( .ZN(N7174), .A1(N7116), .A2(N7023) );
  AND2_X1 AND2_1822( .ZN(N7175), .A1(N6940), .A2(N7023) );
  AND2_X1 AND2_1823( .ZN(N7176), .A1(N5418), .A2(N7023) );
  INV_X1 NOT1_1824( .ZN(N7177), .A(N7041) );
  AND2_X1 AND2_1825( .ZN(N7178), .A1(N7130), .A2(N7049) );
  AND2_X1 AND2_1826( .ZN(N7179), .A1(N7131), .A2(N7049) );
  AND2_X1 AND2_1827( .ZN(N7180), .A1(N6958), .A2(N7049) );
  AND2_X1 AND2_1828( .ZN(N7181), .A1(N5573), .A2(N7049) );
  INV_X2 NOT1_1829( .ZN(N7182), .A(N7065) );
  INV_X1 NOT1_1830( .ZN(N7183), .A(N7094) );
  NAND2_X1 NAND2_1831( .ZN(N7184), .A1(N7094), .A2(N6977) );
  INV_X1 NOT1_1832( .ZN(N7185), .A(N7097) );
  NAND2_X1 NAND2_1833( .ZN(N7186), .A1(N7097), .A2(N6978) );
  AND3_X1 AND3_1834( .ZN(N7187), .A1(N7037), .A2(N1761), .A3(N3108) );
  AND3_X1 AND3_1835( .ZN(N7188), .A1(N7034), .A2(N1761), .A3(N3108) );
  AND3_X1 AND3_1836( .ZN(N7189), .A1(N7031), .A2(N1761), .A3(N3108) );
  OR3_X1 OR3_1837( .ZN(N7190), .A1(N4956), .A2(N7146), .A3(N3781) );
  AND3_X1 AND3_1838( .ZN(N7196), .A1(N7060), .A2(N1777), .A3(N3130) );
  AND3_X1 AND3_1839( .ZN(N7197), .A1(N7057), .A2(N1777), .A3(N3130) );
  OR3_X1 OR3_1840( .ZN(N7198), .A1(N4960), .A2(N7147), .A3(N3786) );
  NAND2_X1 NAND2_1841( .ZN(N7204), .A1(N7101), .A2(N7149) );
  INV_X1 NOT1_1842( .ZN(N7205), .A(N7101) );
  NAND2_X1 NAND2_1843( .ZN(N7206), .A1(N6637), .A2(N7150) );
  AND3_X1 AND3_1844( .ZN(N7207), .A1(N7028), .A2(N1793), .A3(N3158) );
  AND3_X1 AND3_1845( .ZN(N7208), .A1(N7054), .A2(N1807), .A3(N3180) );
  NAND2_X2 NAND2_1846( .ZN(N7209), .A1(N7073), .A2(N7152) );
  NAND2_X1 NAND2_1847( .ZN(N7212), .A1(N7075), .A2(N7153) );
  INV_X1 NOT1_1848( .ZN(N7215), .A(N7076) );
  NAND2_X1 NAND2_1849( .ZN(N7216), .A1(N7076), .A2(N7079) );
  INV_X1 NOT1_1850( .ZN(N7217), .A(N7080) );
  NAND2_X1 NAND2_1851( .ZN(N7218), .A1(N7080), .A2(N7083) );
  NAND2_X1 NAND2_1852( .ZN(N7219), .A1(N7085), .A2(N7158) );
  NAND2_X1 NAND2_1853( .ZN(N7222), .A1(N7087), .A2(N7159) );
  NAND2_X1 NAND2_1854( .ZN(N7225), .A1(N7089), .A2(N7160) );
  INV_X1 NOT1_1855( .ZN(N7228), .A(N7090) );
  NAND2_X1 NAND2_1856( .ZN(N7229), .A1(N7090), .A2(N7093) );
  OR2_X1 OR2_1857( .ZN(N7236), .A1(N7173), .A2(N7125) );
  OR2_X1 OR2_1858( .ZN(N7239), .A1(N7174), .A2(N7126) );
  OR2_X1 OR2_1859( .ZN(N7242), .A1(N7175), .A2(N7127) );
  OR2_X1 OR2_1860( .ZN(N7245), .A1(N7176), .A2(N7040) );
  OR2_X1 OR2_1861( .ZN(N7250), .A1(N7178), .A2(N7139) );
  OR2_X1 OR2_1862( .ZN(N7257), .A1(N7179), .A2(N7140) );
  OR2_X1 OR2_1863( .ZN(N7260), .A1(N7180), .A2(N7141) );
  OR2_X1 OR2_1864( .ZN(N7263), .A1(N7181), .A2(N7064) );
  NAND2_X1 NAND2_1865( .ZN(N7268), .A1(N6792), .A2(N7183) );
  NAND2_X1 NAND2_1866( .ZN(N7269), .A1(N6795), .A2(N7185) );
  OR3_X1 OR3_1867( .ZN(N7270), .A1(N4957), .A2(N7187), .A3(N3782) );
  OR3_X1 OR3_1868( .ZN(N7276), .A1(N4958), .A2(N7188), .A3(N3783) );
  OR3_X1 OR3_1869( .ZN(N7282), .A1(N4959), .A2(N7189), .A3(N3784) );
  OR3_X1 OR3_1870( .ZN(N7288), .A1(N4961), .A2(N7196), .A3(N3787) );
  OR3_X1 OR3_1871( .ZN(N7294), .A1(N3998), .A2(N7197), .A3(N3788) );
  NAND2_X1 NAND2_1872( .ZN(N7300), .A1(N7003), .A2(N7205) );
  NAND2_X1 NAND2_1873( .ZN(N7301), .A1(N7206), .A2(N7151) );
  OR3_X1 OR3_1874( .ZN(N7304), .A1(N4980), .A2(N7207), .A3(N3800) );
  OR3_X1 OR3_1875( .ZN(N7310), .A1(N4984), .A2(N7208), .A3(N3805) );
  NAND2_X1 NAND2_1876( .ZN(N7320), .A1(N6891), .A2(N7215) );
  NAND2_X1 NAND2_1877( .ZN(N7321), .A1(N6897), .A2(N7217) );
  NAND2_X1 NAND2_1878( .ZN(N7328), .A1(N6916), .A2(N7228) );
  AND3_X1 AND3_1879( .ZN(N7338), .A1(N7190), .A2(N1185), .A3(N2692) );
  AND3_X1 AND3_1880( .ZN(N7339), .A1(N7198), .A2(N2681), .A3(N2692) );
  AND3_X1 AND3_1881( .ZN(N7340), .A1(N7190), .A2(N1247), .A3(N2767) );
  AND3_X1 AND3_1882( .ZN(N7341), .A1(N7198), .A2(N2756), .A3(N2767) );
  AND3_X1 AND3_1883( .ZN(N7342), .A1(N7190), .A2(N1327), .A3(N2790) );
  AND3_X1 AND3_1884( .ZN(N7349), .A1(N7198), .A2(N2779), .A3(N2790) );
  AND3_X1 AND3_1885( .ZN(N7357), .A1(N7198), .A2(N2801), .A3(N2812) );
  INV_X1 NOT1_1886( .ZN(N7363), .A(N7198) );
  AND3_X1 AND3_1887( .ZN(N7364), .A1(N7190), .A2(N1351), .A3(N2812) );
  INV_X1 NOT1_1888( .ZN(N7365), .A(N7190) );
  NAND2_X1 NAND2_1889( .ZN(N7394), .A1(N7268), .A2(N7184) );
  NAND2_X1 NAND2_1890( .ZN(N7397), .A1(N7269), .A2(N7186) );
  NAND2_X1 NAND2_1891( .ZN(N7402), .A1(N7204), .A2(N7300) );
  INV_X1 NOT1_1892( .ZN(N7405), .A(N7209) );
  NAND2_X1 NAND2_1893( .ZN(N7406), .A1(N7209), .A2(N6884) );
  INV_X1 NOT1_1894( .ZN(N7407), .A(N7212) );
  NAND2_X1 NAND2_1895( .ZN(N7408), .A1(N7212), .A2(N6888) );
  NAND2_X1 NAND2_1896( .ZN(N7409), .A1(N7320), .A2(N7216) );
  NAND2_X1 NAND2_1897( .ZN(N7412), .A1(N7321), .A2(N7218) );
  INV_X1 NOT1_1898( .ZN(N7415), .A(N7219) );
  NAND2_X1 NAND2_1899( .ZN(N7416), .A1(N7219), .A2(N6904) );
  INV_X1 NOT1_1900( .ZN(N7417), .A(N7222) );
  NAND2_X1 NAND2_1901( .ZN(N7418), .A1(N7222), .A2(N6908) );
  INV_X1 NOT1_1902( .ZN(N7419), .A(N7225) );
  NAND2_X1 NAND2_1903( .ZN(N7420), .A1(N7225), .A2(N6913) );
  NAND2_X1 NAND2_1904( .ZN(N7421), .A1(N7328), .A2(N7229) );
  INV_X1 NOT1_1905( .ZN(N7424), .A(N7245) );
  INV_X1 NOT1_1906( .ZN(N7425), .A(N7242) );
  INV_X2 NOT1_1907( .ZN(N7426), .A(N7239) );
  INV_X2 NOT1_1908( .ZN(N7427), .A(N7236) );
  INV_X2 NOT1_1909( .ZN(N7428), .A(N7263) );
  INV_X1 NOT1_1910( .ZN(N7429), .A(N7260) );
  INV_X1 NOT1_1911( .ZN(N7430), .A(N7257) );
  INV_X1 NOT1_1912( .ZN(N7431), .A(N7250) );
  INV_X1 NOT1_1913( .ZN(N7432), .A(N7250) );
  AND3_X1 AND3_1914( .ZN(N7433), .A1(N7310), .A2(N2653), .A3(N2664) );
  AND3_X1 AND3_1915( .ZN(N7434), .A1(N7304), .A2(N1161), .A3(N2664) );
  OR4_X1 OR4_1916( .ZN(N7435), .A1(N7011), .A2(N7338), .A3(N3621), .A4(N2591) );
  AND3_X1 AND3_1917( .ZN(N7436), .A1(N7270), .A2(N1185), .A3(N2692) );
  AND3_X1 AND3_1918( .ZN(N7437), .A1(N7288), .A2(N2681), .A3(N2692) );
  AND3_X1 AND3_1919( .ZN(N7438), .A1(N7276), .A2(N1185), .A3(N2692) );
  AND3_X1 AND3_1920( .ZN(N7439), .A1(N7294), .A2(N2681), .A3(N2692) );
  AND3_X1 AND3_1921( .ZN(N7440), .A1(N7282), .A2(N1185), .A3(N2692) );
  AND3_X1 AND3_1922( .ZN(N7441), .A1(N7310), .A2(N2728), .A3(N2739) );
  AND3_X1 AND3_1923( .ZN(N7442), .A1(N7304), .A2(N1223), .A3(N2739) );
  OR4_X1 OR4_1924( .ZN(N7443), .A1(N7012), .A2(N7340), .A3(N3632), .A4(N2600) );
  AND3_X1 AND3_1925( .ZN(N7444), .A1(N7270), .A2(N1247), .A3(N2767) );
  AND3_X1 AND3_1926( .ZN(N7445), .A1(N7288), .A2(N2756), .A3(N2767) );
  AND3_X1 AND3_1927( .ZN(N7446), .A1(N7276), .A2(N1247), .A3(N2767) );
  AND3_X1 AND3_1928( .ZN(N7447), .A1(N7294), .A2(N2756), .A3(N2767) );
  AND3_X1 AND3_1929( .ZN(N7448), .A1(N7282), .A2(N1247), .A3(N2767) );
  OR4_X1 OR4_1930( .ZN(N7449), .A1(N7013), .A2(N7342), .A3(N3641), .A4(N2605) );
  AND3_X1 AND3_1931( .ZN(N7450), .A1(N7310), .A2(N3041), .A3(N3052) );
  AND3_X1 AND3_1932( .ZN(N7451), .A1(N7304), .A2(N1697), .A3(N3052) );
  AND3_X1 AND3_1933( .ZN(N7452), .A1(N7294), .A2(N2779), .A3(N2790) );
  AND3_X1 AND3_1934( .ZN(N7453), .A1(N7282), .A2(N1327), .A3(N2790) );
  AND3_X1 AND3_1935( .ZN(N7454), .A1(N7288), .A2(N2779), .A3(N2790) );
  AND3_X1 AND3_1936( .ZN(N7455), .A1(N7276), .A2(N1327), .A3(N2790) );
  AND3_X2 AND3_1937( .ZN(N7456), .A1(N7270), .A2(N1327), .A3(N2790) );
  AND3_X2 AND3_1938( .ZN(N7457), .A1(N7310), .A2(N3075), .A3(N3086) );
  AND3_X2 AND3_1939( .ZN(N7458), .A1(N7304), .A2(N1731), .A3(N3086) );
  AND3_X2 AND3_1940( .ZN(N7459), .A1(N7294), .A2(N2801), .A3(N2812) );
  AND3_X1 AND3_1941( .ZN(N7460), .A1(N7282), .A2(N1351), .A3(N2812) );
  AND3_X1 AND3_1942( .ZN(N7461), .A1(N7288), .A2(N2801), .A3(N2812) );
  AND3_X1 AND3_1943( .ZN(N7462), .A1(N7276), .A2(N1351), .A3(N2812) );
  AND3_X1 AND3_1944( .ZN(N7463), .A1(N7270), .A2(N1351), .A3(N2812) );
  AND3_X1 AND3_1945( .ZN(N7464), .A1(N7250), .A2(N603), .A3(N599) );
  INV_X1 NOT1_1946( .ZN(N7465), .A(N7310) );
  INV_X1 NOT1_1947( .ZN(N7466), .A(N7294) );
  INV_X1 NOT1_1948( .ZN(N7467), .A(N7288) );
  INV_X1 NOT1_1949( .ZN(N7468), .A(N7301) );
  OR4_X1 OR4_1950( .ZN(N7469), .A1(N7016), .A2(N7364), .A3(N3660), .A4(N2626) );
  INV_X1 NOT1_1951( .ZN(N7470), .A(N7304) );
  INV_X1 NOT1_1952( .ZN(N7471), .A(N7282) );
  INV_X1 NOT1_1953( .ZN(N7472), .A(N7276) );
  INV_X1 NOT1_1954( .ZN(N7473), .A(N7270) );
  BUF_X1 BUFF1_1955( .Z(N7474), .A(N7394) );
  BUF_X1 BUFF1_1956( .Z(N7476), .A(N7397) );
  AND2_X1 AND2_1957( .ZN(N7479), .A1(N7301), .A2(N3068) );
  AND3_X1 AND3_1958( .ZN(N7481), .A1(N7245), .A2(N1793), .A3(N3158) );
  AND3_X1 AND3_1959( .ZN(N7482), .A1(N7242), .A2(N1793), .A3(N3158) );
  AND3_X1 AND3_1960( .ZN(N7483), .A1(N7239), .A2(N1793), .A3(N3158) );
  AND3_X1 AND3_1961( .ZN(N7484), .A1(N7236), .A2(N1793), .A3(N3158) );
  AND3_X1 AND3_1962( .ZN(N7485), .A1(N7263), .A2(N1807), .A3(N3180) );
  AND3_X1 AND3_1963( .ZN(N7486), .A1(N7260), .A2(N1807), .A3(N3180) );
  AND3_X1 AND3_1964( .ZN(N7487), .A1(N7257), .A2(N1807), .A3(N3180) );
  AND3_X1 AND3_1965( .ZN(N7488), .A1(N7250), .A2(N1807), .A3(N3180) );
  NAND2_X1 NAND2_1966( .ZN(N7489), .A1(N6979), .A2(N7250) );
  NAND2_X1 NAND2_1967( .ZN(N7492), .A1(N6516), .A2(N7405) );
  NAND2_X1 NAND2_1968( .ZN(N7493), .A1(N6526), .A2(N7407) );
  NAND2_X1 NAND2_1969( .ZN(N7498), .A1(N6592), .A2(N7415) );
  NAND2_X1 NAND2_1970( .ZN(N7499), .A1(N6599), .A2(N7417) );
  NAND2_X1 NAND2_1971( .ZN(N7500), .A1(N6609), .A2(N7419) );
  AND4_X1 AND9_1972_A( .ZN(extra20), .A1(N7105), .A2(N7166), .A3(N7167), .A4(N7168) );
  AND4_X1 AND9_1972_B( .ZN(extra21), .A1(extra20), .A2(N7169), .A3(N7424), .A4(N7425) );
  AND3_X1 AND9_1972( .ZN(N7503), .A1(extra21), .A2(N7426), .A3(N7427) );
  AND4_X1 AND9_1973_A( .ZN(extra22), .A1(N6640), .A2(N7110), .A3(N7170), .A4(N7171) );
  AND4_X1 AND9_1973_B( .ZN(extra23), .A1(extra22), .A2(N7172), .A3(N7428), .A4(N7429) );
  AND3_X1 AND9_1973( .ZN(N7504), .A1(extra23), .A2(N7430), .A3(N7431) );
  OR4_X1 OR4_1974( .ZN(N7505), .A1(N7433), .A2(N7434), .A3(N3616), .A4(N2585) );
  AND2_X1 AND2_1975( .ZN(N7506), .A1(N7435), .A2(N2675) );
  OR4_X1 OR4_1976( .ZN(N7507), .A1(N7339), .A2(N7436), .A3(N3622), .A4(N2592) );
  OR4_X1 OR4_1977( .ZN(N7508), .A1(N7437), .A2(N7438), .A3(N3623), .A4(N2593) );
  OR4_X1 OR4_1978( .ZN(N7509), .A1(N7439), .A2(N7440), .A3(N3624), .A4(N2594) );
  OR4_X1 OR4_1979( .ZN(N7510), .A1(N7441), .A2(N7442), .A3(N3627), .A4(N2595) );
  AND2_X1 AND2_1980( .ZN(N7511), .A1(N7443), .A2(N2750) );
  OR4_X1 OR4_1981( .ZN(N7512), .A1(N7341), .A2(N7444), .A3(N3633), .A4(N2601) );
  OR4_X1 OR4_1982( .ZN(N7513), .A1(N7445), .A2(N7446), .A3(N3634), .A4(N2602) );
  OR4_X1 OR4_1983( .ZN(N7514), .A1(N7447), .A2(N7448), .A3(N3635), .A4(N2603) );
  OR4_X1 OR4_1984( .ZN(N7515), .A1(N7450), .A2(N7451), .A3(N3646), .A4(N2610) );
  OR4_X1 OR4_1985( .ZN(N7516), .A1(N7452), .A2(N7453), .A3(N3647), .A4(N2611) );
  OR4_X1 OR4_1986( .ZN(N7517), .A1(N7454), .A2(N7455), .A3(N3648), .A4(N2612) );
  OR4_X1 OR4_1987( .ZN(N7518), .A1(N7349), .A2(N7456), .A3(N3649), .A4(N2613) );
  OR4_X1 OR4_1988( .ZN(N7519), .A1(N7457), .A2(N7458), .A3(N3654), .A4(N2618) );
  OR4_X1 OR4_1989( .ZN(N7520), .A1(N7459), .A2(N7460), .A3(N3655), .A4(N2619) );
  OR4_X1 OR4_1990( .ZN(N7521), .A1(N7461), .A2(N7462), .A3(N3656), .A4(N2620) );
  OR4_X1 OR4_1991( .ZN(N7522), .A1(N7357), .A2(N7463), .A3(N3657), .A4(N2621) );
  OR4_X1 OR4_1992( .ZN(N7525), .A1(N4741), .A2(N7114), .A3(N2624), .A4(N7464) );
  AND3_X1 AND3_1993( .ZN(N7526), .A1(N7468), .A2(N3119), .A3(N3130) );
  INV_X1 NOT1_1994( .ZN(N7527), .A(N7394) );
  INV_X1 NOT1_1995( .ZN(N7528), .A(N7397) );
  INV_X1 NOT1_1996( .ZN(N7529), .A(N7402) );
  AND2_X1 AND2_1997( .ZN(N7530), .A1(N7402), .A2(N3068) );
  OR3_X1 OR3_1998( .ZN(N7531), .A1(N4981), .A2(N7481), .A3(N3801) );
  OR3_X1 OR3_1999( .ZN(N7537), .A1(N4982), .A2(N7482), .A3(N3802) );
  OR3_X2 OR3_2000( .ZN(N7543), .A1(N4983), .A2(N7483), .A3(N3803) );
  OR3_X2 OR3_2001( .ZN(N7549), .A1(N5165), .A2(N7484), .A3(N3804) );
  OR3_X1 OR3_2002( .ZN(N7555), .A1(N4985), .A2(N7485), .A3(N3806) );
  OR3_X1 OR3_2003( .ZN(N7561), .A1(N4986), .A2(N7486), .A3(N3807) );
  OR3_X1 OR3_2004( .ZN(N7567), .A1(N4547), .A2(N7487), .A3(N3808) );
  OR3_X1 OR3_2005( .ZN(N7573), .A1(N4987), .A2(N7488), .A3(N3809) );
  NAND2_X1 NAND2_2006( .ZN(N7579), .A1(N7492), .A2(N7406) );
  NAND2_X1 NAND2_2007( .ZN(N7582), .A1(N7493), .A2(N7408) );
  INV_X1 NOT1_2008( .ZN(N7585), .A(N7409) );
  NAND2_X1 NAND2_2009( .ZN(N7586), .A1(N7409), .A2(N6894) );
  INV_X1 NOT1_2010( .ZN(N7587), .A(N7412) );
  NAND2_X1 NAND2_2011( .ZN(N7588), .A1(N7412), .A2(N6900) );
  NAND2_X1 NAND2_2012( .ZN(N7589), .A1(N7498), .A2(N7416) );
  NAND2_X1 NAND2_2013( .ZN(N7592), .A1(N7499), .A2(N7418) );
  NAND2_X1 NAND2_2014( .ZN(N7595), .A1(N7500), .A2(N7420) );
  INV_X1 NOT1_2015( .ZN(N7598), .A(N7421) );
  NAND2_X1 NAND2_2016( .ZN(N7599), .A1(N7421), .A2(N6919) );
  AND2_X1 AND2_2017( .ZN(N7600), .A1(N7505), .A2(N2647) );
  AND2_X1 AND2_2018( .ZN(N7601), .A1(N7507), .A2(N2675) );
  AND2_X1 AND2_2019( .ZN(N7602), .A1(N7508), .A2(N2675) );
  AND2_X1 AND2_2020( .ZN(N7603), .A1(N7509), .A2(N2675) );
  AND2_X1 AND2_2021( .ZN(N7604), .A1(N7510), .A2(N2722) );
  AND2_X1 AND2_2022( .ZN(N7605), .A1(N7512), .A2(N2750) );
  AND2_X2 AND2_2023( .ZN(N7606), .A1(N7513), .A2(N2750) );
  AND2_X2 AND2_2024( .ZN(N7607), .A1(N7514), .A2(N2750) );
  AND2_X2 AND2_2025( .ZN(N7624), .A1(N6979), .A2(N7489) );
  AND2_X1 AND2_2026( .ZN(N7625), .A1(N7489), .A2(N7250) );
  AND2_X1 AND2_2027( .ZN(N7626), .A1(N1149), .A2(N7525) );
  AND4_X1 AND5_2028_A( .ZN(extra24), .A1(N562), .A2(N7527), .A3(N7528), .A4(N6805) );
  AND2_X1 AND5_2028( .ZN(N7631), .A1(extra24), .A2(N6930) );
  AND3_X1 AND3_2029( .ZN(N7636), .A1(N7529), .A2(N3097), .A3(N3108) );
  NAND2_X1 NAND2_2030( .ZN(N7657), .A1(N6539), .A2(N7585) );
  NAND2_X1 NAND2_2031( .ZN(N7658), .A1(N6556), .A2(N7587) );
  NAND2_X1 NAND2_2032( .ZN(N7665), .A1(N6622), .A2(N7598) );
  AND3_X1 AND3_2033( .ZN(N7666), .A1(N7555), .A2(N2653), .A3(N2664) );
  AND3_X1 AND3_2034( .ZN(N7667), .A1(N7531), .A2(N1161), .A3(N2664) );
  AND3_X1 AND3_2035( .ZN(N7668), .A1(N7561), .A2(N2653), .A3(N2664) );
  AND3_X1 AND3_2036( .ZN(N7669), .A1(N7537), .A2(N1161), .A3(N2664) );
  AND3_X1 AND3_2037( .ZN(N7670), .A1(N7567), .A2(N2653), .A3(N2664) );
  AND3_X1 AND3_2038( .ZN(N7671), .A1(N7543), .A2(N1161), .A3(N2664) );
  AND3_X1 AND3_2039( .ZN(N7672), .A1(N7573), .A2(N2653), .A3(N2664) );
  AND3_X1 AND3_2040( .ZN(N7673), .A1(N7549), .A2(N1161), .A3(N2664) );
  AND3_X1 AND3_2041( .ZN(N7674), .A1(N7555), .A2(N2728), .A3(N2739) );
  AND3_X1 AND3_2042( .ZN(N7675), .A1(N7531), .A2(N1223), .A3(N2739) );
  AND3_X1 AND3_2043( .ZN(N7676), .A1(N7561), .A2(N2728), .A3(N2739) );
  AND3_X1 AND3_2044( .ZN(N7677), .A1(N7537), .A2(N1223), .A3(N2739) );
  AND3_X1 AND3_2045( .ZN(N7678), .A1(N7567), .A2(N2728), .A3(N2739) );
  AND3_X1 AND3_2046( .ZN(N7679), .A1(N7543), .A2(N1223), .A3(N2739) );
  AND3_X1 AND3_2047( .ZN(N7680), .A1(N7573), .A2(N2728), .A3(N2739) );
  AND3_X1 AND3_2048( .ZN(N7681), .A1(N7549), .A2(N1223), .A3(N2739) );
  AND3_X1 AND3_2049( .ZN(N7682), .A1(N7573), .A2(N3075), .A3(N3086) );
  AND3_X1 AND3_2050( .ZN(N7683), .A1(N7549), .A2(N1731), .A3(N3086) );
  AND3_X2 AND3_2051( .ZN(N7684), .A1(N7573), .A2(N3041), .A3(N3052) );
  AND3_X2 AND3_2052( .ZN(N7685), .A1(N7549), .A2(N1697), .A3(N3052) );
  AND3_X2 AND3_2053( .ZN(N7686), .A1(N7567), .A2(N3041), .A3(N3052) );
  AND3_X2 AND3_2054( .ZN(N7687), .A1(N7543), .A2(N1697), .A3(N3052) );
  AND3_X1 AND3_2055( .ZN(N7688), .A1(N7561), .A2(N3041), .A3(N3052) );
  AND3_X1 AND3_2056( .ZN(N7689), .A1(N7537), .A2(N1697), .A3(N3052) );
  AND3_X1 AND3_2057( .ZN(N7690), .A1(N7555), .A2(N3041), .A3(N3052) );
  AND3_X1 AND3_2058( .ZN(N7691), .A1(N7531), .A2(N1697), .A3(N3052) );
  AND3_X1 AND3_2059( .ZN(N7692), .A1(N7567), .A2(N3075), .A3(N3086) );
  AND3_X1 AND3_2060( .ZN(N7693), .A1(N7543), .A2(N1731), .A3(N3086) );
  AND3_X1 AND3_2061( .ZN(N7694), .A1(N7561), .A2(N3075), .A3(N3086) );
  AND3_X1 AND3_2062( .ZN(N7695), .A1(N7537), .A2(N1731), .A3(N3086) );
  AND3_X1 AND3_2063( .ZN(N7696), .A1(N7555), .A2(N3075), .A3(N3086) );
  AND3_X1 AND3_2064( .ZN(N7697), .A1(N7531), .A2(N1731), .A3(N3086) );
  OR2_X1 OR2_2065( .ZN(N7698), .A1(N7624), .A2(N7625) );
  INV_X1 NOT1_2066( .ZN(N7699), .A(N7573) );
  INV_X1 NOT1_2067( .ZN(N7700), .A(N7567) );
  INV_X1 NOT1_2068( .ZN(N7701), .A(N7561) );
  INV_X1 NOT1_2069( .ZN(N7702), .A(N7555) );
  AND3_X1 AND3_2070( .ZN(N7703), .A1(N1156), .A2(N7631), .A3(N245) );
  INV_X1 NOT1_2071( .ZN(N7704), .A(N7549) );
  INV_X1 NOT1_2072( .ZN(N7705), .A(N7543) );
  INV_X1 NOT1_2073( .ZN(N7706), .A(N7537) );
  INV_X1 NOT1_2074( .ZN(N7707), .A(N7531) );
  INV_X1 NOT1_2075( .ZN(N7708), .A(N7579) );
  NAND2_X1 NAND2_2076( .ZN(N7709), .A1(N7579), .A2(N6739) );
  INV_X1 NOT1_2077( .ZN(N7710), .A(N7582) );
  NAND2_X1 NAND2_2078( .ZN(N7711), .A1(N7582), .A2(N6744) );
  NAND2_X1 NAND2_2079( .ZN(N7712), .A1(N7657), .A2(N7586) );
  NAND2_X1 NAND2_2080( .ZN(N7715), .A1(N7658), .A2(N7588) );
  INV_X1 NOT1_2081( .ZN(N7718), .A(N7589) );
  NAND2_X1 NAND2_2082( .ZN(N7719), .A1(N7589), .A2(N6772) );
  INV_X1 NOT1_2083( .ZN(N7720), .A(N7592) );
  NAND2_X1 NAND2_2084( .ZN(N7721), .A1(N7592), .A2(N6776) );
  INV_X1 NOT1_2085( .ZN(N7722), .A(N7595) );
  NAND2_X1 NAND2_2086( .ZN(N7723), .A1(N7595), .A2(N5733) );
  NAND2_X1 NAND2_2087( .ZN(N7724), .A1(N7665), .A2(N7599) );
  OR4_X1 OR4_2088( .ZN(N7727), .A1(N7666), .A2(N7667), .A3(N3617), .A4(N2586) );
  OR4_X1 OR4_2089( .ZN(N7728), .A1(N7668), .A2(N7669), .A3(N3618), .A4(N2587) );
  OR4_X1 OR4_2090( .ZN(N7729), .A1(N7670), .A2(N7671), .A3(N3619), .A4(N2588) );
  OR4_X1 OR4_2091( .ZN(N7730), .A1(N7672), .A2(N7673), .A3(N3620), .A4(N2589) );
  OR4_X1 OR4_2092( .ZN(N7731), .A1(N7674), .A2(N7675), .A3(N3628), .A4(N2596) );
  OR4_X1 OR4_2093( .ZN(N7732), .A1(N7676), .A2(N7677), .A3(N3629), .A4(N2597) );
  OR4_X1 OR4_2094( .ZN(N7733), .A1(N7678), .A2(N7679), .A3(N3630), .A4(N2598) );
  OR4_X1 OR4_2095( .ZN(N7734), .A1(N7680), .A2(N7681), .A3(N3631), .A4(N2599) );
  OR4_X1 OR4_2096( .ZN(N7735), .A1(N7682), .A2(N7683), .A3(N3638), .A4(N2604) );
  OR4_X1 OR4_2097( .ZN(N7736), .A1(N7684), .A2(N7685), .A3(N3642), .A4(N2606) );
  OR4_X1 OR4_2098( .ZN(N7737), .A1(N7686), .A2(N7687), .A3(N3643), .A4(N2607) );
  OR4_X1 OR4_2099( .ZN(N7738), .A1(N7688), .A2(N7689), .A3(N3644), .A4(N2608) );
  OR4_X1 OR4_2100( .ZN(N7739), .A1(N7690), .A2(N7691), .A3(N3645), .A4(N2609) );
  OR4_X1 OR4_2101( .ZN(N7740), .A1(N7692), .A2(N7693), .A3(N3651), .A4(N2615) );
  OR4_X1 OR4_2102( .ZN(N7741), .A1(N7694), .A2(N7695), .A3(N3652), .A4(N2616) );
  OR4_X1 OR4_2103( .ZN(N7742), .A1(N7696), .A2(N7697), .A3(N3653), .A4(N2617) );
  NAND2_X1 NAND2_2104( .ZN(N7743), .A1(N6271), .A2(N7708) );
  NAND2_X1 NAND2_2105( .ZN(N7744), .A1(N6283), .A2(N7710) );
  NAND2_X1 NAND2_2106( .ZN(N7749), .A1(N6341), .A2(N7718) );
  NAND2_X1 NAND2_2107( .ZN(N7750), .A1(N6347), .A2(N7720) );
  NAND2_X1 NAND2_2108( .ZN(N7751), .A1(N5214), .A2(N7722) );
  AND2_X1 AND2_2109( .ZN(N7754), .A1(N7727), .A2(N2647) );
  AND2_X1 AND2_2110( .ZN(N7755), .A1(N7728), .A2(N2647) );
  AND2_X1 AND2_2111( .ZN(N7756), .A1(N7729), .A2(N2647) );
  AND2_X4 AND2_2112( .ZN(N7757), .A1(N7730), .A2(N2647) );
  AND2_X1 AND2_2113( .ZN(N7758), .A1(N7731), .A2(N2722) );
  AND2_X1 AND2_2114( .ZN(N7759), .A1(N7732), .A2(N2722) );
  AND2_X1 AND2_2115( .ZN(N7760), .A1(N7733), .A2(N2722) );
  AND2_X1 AND2_2116( .ZN(N7761), .A1(N7734), .A2(N2722) );
  NAND2_X1 NAND2_2117( .ZN(N7762), .A1(N7743), .A2(N7709) );
  NAND2_X1 NAND2_2118( .ZN(N7765), .A1(N7744), .A2(N7711) );
  INV_X1 NOT1_2119( .ZN(N7768), .A(N7712) );
  NAND2_X1 NAND2_2120( .ZN(N7769), .A1(N7712), .A2(N6751) );
  INV_X1 NOT1_2121( .ZN(N7770), .A(N7715) );
  NAND2_X1 NAND2_2122( .ZN(N7771), .A1(N7715), .A2(N6760) );
  NAND2_X1 NAND2_2123( .ZN(N7772), .A1(N7749), .A2(N7719) );
  NAND2_X1 NAND2_2124( .ZN(N7775), .A1(N7750), .A2(N7721) );
  NAND2_X1 NAND2_2125( .ZN(N7778), .A1(N7751), .A2(N7723) );
  INV_X1 NOT1_2126( .ZN(N7781), .A(N7724) );
  NAND2_X1 NAND2_2127( .ZN(N7782), .A1(N7724), .A2(N5735) );
  NAND2_X1 NAND2_2128( .ZN(N7787), .A1(N6295), .A2(N7768) );
  NAND2_X1 NAND2_2129( .ZN(N7788), .A1(N6313), .A2(N7770) );
  NAND2_X1 NAND2_2130( .ZN(N7795), .A1(N5220), .A2(N7781) );
  INV_X1 NOT1_2131( .ZN(N7796), .A(N7762) );
  NAND2_X1 NAND2_2132( .ZN(N7797), .A1(N7762), .A2(N6740) );
  INV_X1 NOT1_2133( .ZN(N7798), .A(N7765) );
  NAND2_X1 NAND2_2134( .ZN(N7799), .A1(N7765), .A2(N6745) );
  NAND2_X1 NAND2_2135( .ZN(N7800), .A1(N7787), .A2(N7769) );
  NAND2_X1 NAND2_2136( .ZN(N7803), .A1(N7788), .A2(N7771) );
  INV_X1 NOT1_2137( .ZN(N7806), .A(N7772) );
  NAND2_X1 NAND2_2138( .ZN(N7807), .A1(N7772), .A2(N6773) );
  INV_X1 NOT1_2139( .ZN(N7808), .A(N7775) );
  NAND2_X1 NAND2_2140( .ZN(N7809), .A1(N7775), .A2(N6777) );
  INV_X1 NOT1_2141( .ZN(N7810), .A(N7778) );
  NAND2_X1 NAND2_2142( .ZN(N7811), .A1(N7778), .A2(N6782) );
  NAND2_X1 NAND2_2143( .ZN(N7812), .A1(N7795), .A2(N7782) );
  NAND2_X1 NAND2_2144( .ZN(N7815), .A1(N6274), .A2(N7796) );
  NAND2_X1 NAND2_2145( .ZN(N7816), .A1(N6286), .A2(N7798) );
  NAND2_X1 NAND2_2146( .ZN(N7821), .A1(N6344), .A2(N7806) );
  NAND2_X1 NAND2_2147( .ZN(N7822), .A1(N6350), .A2(N7808) );
  NAND2_X1 NAND2_2148( .ZN(N7823), .A1(N6353), .A2(N7810) );
  NAND2_X1 NAND2_2149( .ZN(N7826), .A1(N7815), .A2(N7797) );
  NAND2_X1 NAND2_2150( .ZN(N7829), .A1(N7816), .A2(N7799) );
  INV_X1 NOT1_2151( .ZN(N7832), .A(N7800) );
  NAND2_X1 NAND2_2152( .ZN(N7833), .A1(N7800), .A2(N6752) );
  INV_X1 NOT1_2153( .ZN(N7834), .A(N7803) );
  NAND2_X1 NAND2_2154( .ZN(N7835), .A1(N7803), .A2(N6761) );
  NAND2_X1 NAND2_2155( .ZN(N7836), .A1(N7821), .A2(N7807) );
  NAND2_X1 NAND2_2156( .ZN(N7839), .A1(N7822), .A2(N7809) );
  NAND2_X1 NAND2_2157( .ZN(N7842), .A1(N7823), .A2(N7811) );
  INV_X1 NOT1_2158( .ZN(N7845), .A(N7812) );
  NAND2_X1 NAND2_2159( .ZN(N7846), .A1(N7812), .A2(N6790) );
  NAND2_X1 NAND2_2160( .ZN(N7851), .A1(N6298), .A2(N7832) );
  NAND2_X1 NAND2_2161( .ZN(N7852), .A1(N6316), .A2(N7834) );
  NAND2_X1 NAND2_2162( .ZN(N7859), .A1(N6364), .A2(N7845) );
  INV_X1 NOT1_2163( .ZN(N7860), .A(N7826) );
  NAND2_X1 NAND2_2164( .ZN(N7861), .A1(N7826), .A2(N6741) );
  INV_X1 NOT1_2165( .ZN(N7862), .A(N7829) );
  NAND2_X1 NAND2_2166( .ZN(N7863), .A1(N7829), .A2(N6746) );
  NAND2_X1 NAND2_2167( .ZN(N7864), .A1(N7851), .A2(N7833) );
  NAND2_X1 NAND2_2168( .ZN(N7867), .A1(N7852), .A2(N7835) );
  INV_X1 NOT1_2169( .ZN(N7870), .A(N7836) );
  NAND2_X1 NAND2_2170( .ZN(N7871), .A1(N7836), .A2(N5730) );
  INV_X1 NOT1_2171( .ZN(N7872), .A(N7839) );
  NAND2_X1 NAND2_2172( .ZN(N7873), .A1(N7839), .A2(N5732) );
  INV_X1 NOT1_2173( .ZN(N7874), .A(N7842) );
  NAND2_X1 NAND2_2174( .ZN(N7875), .A1(N7842), .A2(N6783) );
  NAND2_X1 NAND2_2175( .ZN(N7876), .A1(N7859), .A2(N7846) );
  NAND2_X2 NAND2_2176( .ZN(N7879), .A1(N6277), .A2(N7860) );
  NAND2_X2 NAND2_2177( .ZN(N7880), .A1(N6289), .A2(N7862) );
  NAND2_X4 NAND2_2178( .ZN(N7885), .A1(N5199), .A2(N7870) );
  NAND2_X1 NAND2_2179( .ZN(N7886), .A1(N5208), .A2(N7872) );
  NAND2_X1 NAND2_2180( .ZN(N7887), .A1(N6356), .A2(N7874) );
  NAND2_X1 NAND2_2181( .ZN(N7890), .A1(N7879), .A2(N7861) );
  NAND2_X1 NAND2_2182( .ZN(N7893), .A1(N7880), .A2(N7863) );
  INV_X1 NOT1_2183( .ZN(N7896), .A(N7864) );
  NAND2_X1 NAND2_2184( .ZN(N7897), .A1(N7864), .A2(N6753) );
  INV_X1 NOT1_2185( .ZN(N7898), .A(N7867) );
  NAND2_X1 NAND2_2186( .ZN(N7899), .A1(N7867), .A2(N6762) );
  NAND2_X1 NAND2_2187( .ZN(N7900), .A1(N7885), .A2(N7871) );
  NAND2_X1 NAND2_2188( .ZN(N7903), .A1(N7886), .A2(N7873) );
  NAND2_X1 NAND2_2189( .ZN(N7906), .A1(N7887), .A2(N7875) );
  INV_X1 NOT1_2190( .ZN(N7909), .A(N7876) );
  NAND2_X1 NAND2_2191( .ZN(N7910), .A1(N7876), .A2(N6791) );
  NAND2_X1 NAND2_2192( .ZN(N7917), .A1(N6301), .A2(N7896) );
  NAND2_X1 NAND2_2193( .ZN(N7918), .A1(N6319), .A2(N7898) );
  NAND2_X1 NAND2_2194( .ZN(N7923), .A1(N6367), .A2(N7909) );
  INV_X1 NOT1_2195( .ZN(N7924), .A(N7890) );
  NAND2_X1 NAND2_2196( .ZN(N7925), .A1(N7890), .A2(N6680) );
  INV_X1 NOT1_2197( .ZN(N7926), .A(N7893) );
  NAND2_X1 NAND2_2198( .ZN(N7927), .A1(N7893), .A2(N6681) );
  INV_X1 NOT1_2199( .ZN(N7928), .A(N7900) );
  NAND2_X1 NAND2_2200( .ZN(N7929), .A1(N7900), .A2(N5690) );
  INV_X1 NOT1_2201( .ZN(N7930), .A(N7903) );
  NAND2_X1 NAND2_2202( .ZN(N7931), .A1(N7903), .A2(N5691) );
  NAND2_X1 NAND2_2203( .ZN(N7932), .A1(N7917), .A2(N7897) );
  NAND2_X1 NAND2_2204( .ZN(N7935), .A1(N7918), .A2(N7899) );
  INV_X1 NOT1_2205( .ZN(N7938), .A(N7906) );
  NAND2_X1 NAND2_2206( .ZN(N7939), .A1(N7906), .A2(N6784) );
  NAND2_X1 NAND2_2207( .ZN(N7940), .A1(N7923), .A2(N7910) );
  NAND2_X1 NAND2_2208( .ZN(N7943), .A1(N6280), .A2(N7924) );
  NAND2_X1 NAND2_2209( .ZN(N7944), .A1(N6292), .A2(N7926) );
  NAND2_X1 NAND2_2210( .ZN(N7945), .A1(N5202), .A2(N7928) );
  NAND2_X1 NAND2_2211( .ZN(N7946), .A1(N5211), .A2(N7930) );
  NAND2_X1 NAND2_2212( .ZN(N7951), .A1(N6359), .A2(N7938) );
  NAND2_X1 NAND2_2213( .ZN(N7954), .A1(N7943), .A2(N7925) );
  NAND2_X1 NAND2_2214( .ZN(N7957), .A1(N7944), .A2(N7927) );
  NAND2_X1 NAND2_2215( .ZN(N7960), .A1(N7945), .A2(N7929) );
  NAND2_X1 NAND2_2216( .ZN(N7963), .A1(N7946), .A2(N7931) );
  INV_X1 NOT1_2217( .ZN(N7966), .A(N7932) );
  NAND2_X1 NAND2_2218( .ZN(N7967), .A1(N7932), .A2(N6754) );
  INV_X1 NOT1_2219( .ZN(N7968), .A(N7935) );
  NAND2_X1 NAND2_2220( .ZN(N7969), .A1(N7935), .A2(N6755) );
  NAND2_X1 NAND2_2221( .ZN(N7970), .A1(N7951), .A2(N7939) );
  INV_X1 NOT1_2222( .ZN(N7973), .A(N7940) );
  NAND2_X1 NAND2_2223( .ZN(N7974), .A1(N7940), .A2(N6785) );
  NAND2_X1 NAND2_2224( .ZN(N7984), .A1(N6304), .A2(N7966) );
  NAND2_X1 NAND2_2225( .ZN(N7985), .A1(N6322), .A2(N7968) );
  NAND2_X1 NAND2_2226( .ZN(N7987), .A1(N6370), .A2(N7973) );
  AND3_X1 AND3_2227( .ZN(N7988), .A1(N7957), .A2(N6831), .A3(N1157) );
  AND3_X1 AND3_2228( .ZN(N7989), .A1(N7954), .A2(N6415), .A3(N1157) );
  AND3_X1 AND3_2229( .ZN(N7990), .A1(N7957), .A2(N7041), .A3(N566) );
  AND3_X1 AND3_2230( .ZN(N7991), .A1(N7954), .A2(N7177), .A3(N566) );
  INV_X1 NOT1_2231( .ZN(N7992), .A(N7970) );
  NAND2_X1 NAND2_2232( .ZN(N7993), .A1(N7970), .A2(N6448) );
  AND3_X1 AND3_2233( .ZN(N7994), .A1(N7963), .A2(N6857), .A3(N1219) );
  AND3_X1 AND3_2234( .ZN(N7995), .A1(N7960), .A2(N6441), .A3(N1219) );
  AND3_X1 AND3_2235( .ZN(N7996), .A1(N7963), .A2(N7065), .A3(N583) );
  AND3_X1 AND3_2236( .ZN(N7997), .A1(N7960), .A2(N7182), .A3(N583) );
  NAND2_X1 NAND2_2237( .ZN(N7998), .A1(N7984), .A2(N7967) );
  NAND2_X1 NAND2_2238( .ZN(N8001), .A1(N7985), .A2(N7969) );
  NAND2_X1 NAND2_2239( .ZN(N8004), .A1(N7987), .A2(N7974) );
  NAND2_X1 NAND2_2240( .ZN(N8009), .A1(N6051), .A2(N7992) );
  OR4_X1 OR4_2241( .ZN(N8013), .A1(N7988), .A2(N7989), .A3(N7990), .A4(N7991) );
  OR4_X1 OR4_2242( .ZN(N8017), .A1(N7994), .A2(N7995), .A3(N7996), .A4(N7997) );
  INV_X1 NOT1_2243( .ZN(N8020), .A(N7998) );
  NAND2_X1 NAND2_2244( .ZN(N8021), .A1(N7998), .A2(N6682) );
  INV_X1 NOT1_2245( .ZN(N8022), .A(N8001) );
  NAND2_X1 NAND2_2246( .ZN(N8023), .A1(N8001), .A2(N6683) );
  NAND2_X1 NAND2_2247( .ZN(N8025), .A1(N8009), .A2(N7993) );
  INV_X1 NOT1_2248( .ZN(N8026), .A(N8004) );
  NAND2_X1 NAND2_2249( .ZN(N8027), .A1(N8004), .A2(N6449) );
  NAND2_X1 NAND2_2250( .ZN(N8031), .A1(N6307), .A2(N8020) );
  NAND2_X1 NAND2_2251( .ZN(N8032), .A1(N6310), .A2(N8022) );
  INV_X1 NOT1_2252( .ZN(N8033), .A(N8013) );
  NAND2_X1 NAND2_2253( .ZN(N8034), .A1(N6054), .A2(N8026) );
  AND2_X1 AND2_2254( .ZN(N8035), .A1(N583), .A2(N8025) );
  INV_X1 NOT1_2255( .ZN(N8036), .A(N8017) );
  NAND2_X1 NAND2_2256( .ZN(N8037), .A1(N8031), .A2(N8021) );
  NAND2_X1 NAND2_2257( .ZN(N8038), .A1(N8032), .A2(N8023) );
  NAND2_X1 NAND2_2258( .ZN(N8039), .A1(N8034), .A2(N8027) );
  INV_X1 NOT1_2259( .ZN(N8040), .A(N8038) );
  AND2_X1 AND2_2260( .ZN(N8041), .A1(N566), .A2(N8037) );
  INV_X1 NOT1_2261( .ZN(N8042), .A(N8039) );
  AND2_X1 AND2_2262( .ZN(N8043), .A1(N8040), .A2(N1157) );
  AND2_X1 AND2_2263( .ZN(N8044), .A1(N8042), .A2(N1219) );
  OR2_X1 OR2_2264( .ZN(N8045), .A1(N8043), .A2(N8041) );
  OR2_X1 OR2_2265( .ZN(N8048), .A1(N8044), .A2(N8035) );
  NAND2_X1 NAND2_2266( .ZN(N8055), .A1(N8045), .A2(N8033) );
  INV_X1 NOT1_2267( .ZN(N8056), .A(N8045) );
  NAND2_X1 NAND2_2268( .ZN(N8057), .A1(N8048), .A2(N8036) );
  INV_X1 NOT1_2269( .ZN(N8058), .A(N8048) );
  NAND2_X1 NAND2_2270( .ZN(N8059), .A1(N8013), .A2(N8056) );
  NAND2_X1 NAND2_2271( .ZN(N8060), .A1(N8017), .A2(N8058) );
  NAND2_X2 NAND2_2272( .ZN(N8061), .A1(N8055), .A2(N8059) );
  NAND2_X1 NAND2_2273( .ZN(N8064), .A1(N8057), .A2(N8060) );
  AND3_X1 AND3_2274( .ZN(N8071), .A1(N8064), .A2(N1777), .A3(N3130) );
  AND3_X1 AND3_2275( .ZN(N8072), .A1(N8061), .A2(N1761), .A3(N3108) );
  INV_X1 NOT1_2276( .ZN(N8073), .A(N8061) );
  INV_X1 NOT1_2277( .ZN(N8074), .A(N8064) );
  OR4_X1 OR4_2278( .ZN(N8075), .A1(N7526), .A2(N8071), .A3(N3659), .A4(N2625) );
  OR4_X1 OR4_2279( .ZN(N8076), .A1(N7636), .A2(N8072), .A3(N3661), .A4(N2627) );
  AND2_X1 AND2_2280( .ZN(N8077), .A1(N8073), .A2(N1727) );
  AND2_X1 AND2_2281( .ZN(N8078), .A1(N8074), .A2(N1727) );
  OR2_X1 OR2_2282( .ZN(N8079), .A1(N7530), .A2(N8077) );
  OR2_X1 OR2_2283( .ZN(N8082), .A1(N7479), .A2(N8078) );
  AND2_X1 AND2_2284( .ZN(N8089), .A1(N8079), .A2(N3063) );
  AND2_X1 AND2_2285( .ZN(N8090), .A1(N8082), .A2(N3063) );
  AND2_X1 AND2_2286( .ZN(N8091), .A1(N8079), .A2(N3063) );
  AND2_X1 AND2_2287( .ZN(N8092), .A1(N8082), .A2(N3063) );
  OR2_X1 OR2_2288( .ZN(N8093), .A1(N8089), .A2(N3071) );
  OR2_X1 OR2_2289( .ZN(N8096), .A1(N8090), .A2(N3072) );
  OR2_X1 OR2_2290( .ZN(N8099), .A1(N8091), .A2(N3073) );
  OR2_X1 OR2_2291( .ZN(N8102), .A1(N8092), .A2(N3074) );
  AND3_X1 AND3_2292( .ZN(N8113), .A1(N8102), .A2(N2779), .A3(N2790) );
  AND3_X2 AND3_2293( .ZN(N8114), .A1(N8099), .A2(N1327), .A3(N2790) );
  AND3_X2 AND3_2294( .ZN(N8115), .A1(N8102), .A2(N2801), .A3(N2812) );
  AND3_X2 AND3_2295( .ZN(N8116), .A1(N8099), .A2(N1351), .A3(N2812) );
  AND3_X1 AND3_2296( .ZN(N8117), .A1(N8096), .A2(N2681), .A3(N2692) );
  AND3_X1 AND3_2297( .ZN(N8118), .A1(N8093), .A2(N1185), .A3(N2692) );
  AND3_X1 AND3_2298( .ZN(N8119), .A1(N8096), .A2(N2756), .A3(N2767) );
  AND3_X1 AND3_2299( .ZN(N8120), .A1(N8093), .A2(N1247), .A3(N2767) );
  OR4_X1 OR4_2300( .ZN(N8121), .A1(N8117), .A2(N8118), .A3(N3662), .A4(N2703) );
  OR4_X1 OR4_2301( .ZN(N8122), .A1(N8119), .A2(N8120), .A3(N3663), .A4(N2778) );
  OR4_X1 OR4_2302( .ZN(N8123), .A1(N8113), .A2(N8114), .A3(N3650), .A4(N2614) );
  OR4_X1 OR4_2303( .ZN(N8124), .A1(N8115), .A2(N8116), .A3(N3658), .A4(N2622) );
  AND2_X1 AND2_2304( .ZN(N8125), .A1(N8121), .A2(N2675) );
  AND2_X1 AND2_2305( .ZN(N8126), .A1(N8122), .A2(N2750) );
  INV_X1 NOT1_2306( .ZN(N8127), .A(N8125) );
  INV_X1 NOT1_2307( .ZN(N8128), .A(N8126) );

endmodule
