
module c1355(G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,
  G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,
  G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,
  G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,
  G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
  G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,
  G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;

  wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,G284,G287,
    G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,G329,G332,G335,
    G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,G366,G367,G368,G369,
    G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,G381,G382,G383,G384,G385,
    G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,G401,
    G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,
    G418,G419,G420,G421,G422,G423,G424,G425,G426,G429,G432,G435,G438,G441,G444,G447,
    G450,G453,G456,G459,G462,G465,G468,G471,G474,G477,G480,G483,G486,G489,G492,G495,
    G498,G501,G504,G507,G510,G513,G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,
    G546,G549,G552,G555,G558,G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,
    G578,G579,G580,G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,
    G594,G595,G596,G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,
    G642,G645,G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,
    G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,
    G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,G751,
    G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,G768,G769,
    G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,G809,G812,G815,
    G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,
    G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,G941,G942,G943,G944,G945,
    G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,G961,
    G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,
    G978,G979,G980,G981,G982,G983,G984,G985,G986,G991,G996,G1001,G1006,G1011,G1016,G1021,
    G1026,G1031,G1036,G1039,G1042,G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,
    G1078,G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,G1117,G1120,G1123,
    G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,G1153,G1156,G1159,G1162,G1165,G1168,G1171,
    G1174,G1177,G1180,G1183,G1186,G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,
    G1222,G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,G1241,
    G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,
    G1258,G1259,G1260,G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,
    G1274,G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,
    G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,G1301,G1302,G1303,G1304,G1305,
    G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,
    G1322,G1323,extra0,extra1,extra2,extra3,extra4,extra5,extra6,extra7;

  AND2_X1 AND2_0( .ZN(G242), .A1(G33), .A2(G41) );
  AND2_X1 AND2_1( .ZN(G245), .A1(G34), .A2(G41) );
  AND2_X1 AND2_2( .ZN(G248), .A1(G35), .A2(G41) );
  AND2_X1 AND2_3( .ZN(G251), .A1(G36), .A2(G41) );
  AND2_X1 AND2_4( .ZN(G254), .A1(G37), .A2(G41) );
  AND2_X1 AND2_5( .ZN(G257), .A1(G38), .A2(G41) );
  AND2_X1 AND2_6( .ZN(G260), .A1(G39), .A2(G41) );
  AND2_X1 AND2_7( .ZN(G263), .A1(G40), .A2(G41) );
  NAND2_X2 NAND2_0( .ZN(G266), .A1(G1), .A2(G2) );
  NAND2_X2 NAND2_1( .ZN(G269), .A1(G3), .A2(G4) );
  NAND2_X2 NAND2_2( .ZN(G272), .A1(G5), .A2(G6) );
  NAND2_X2 NAND2_3( .ZN(G275), .A1(G7), .A2(G8) );
  NAND2_X1 NAND2_4( .ZN(G278), .A1(G9), .A2(G10) );
  NAND2_X1 NAND2_5( .ZN(G281), .A1(G11), .A2(G12) );
  NAND2_X1 NAND2_6( .ZN(G284), .A1(G13), .A2(G14) );
  NAND2_X1 NAND2_7( .ZN(G287), .A1(G15), .A2(G16) );
  NAND2_X1 NAND2_8( .ZN(G290), .A1(G17), .A2(G18) );
  NAND2_X1 NAND2_9( .ZN(G293), .A1(G19), .A2(G20) );
  NAND2_X1 NAND2_10( .ZN(G296), .A1(G21), .A2(G22) );
  NAND2_X1 NAND2_11( .ZN(G299), .A1(G23), .A2(G24) );
  NAND2_X1 NAND2_12( .ZN(G302), .A1(G25), .A2(G26) );
  NAND2_X2 NAND2_13( .ZN(G305), .A1(G27), .A2(G28) );
  NAND2_X2 NAND2_14( .ZN(G308), .A1(G29), .A2(G30) );
  NAND2_X2 NAND2_15( .ZN(G311), .A1(G31), .A2(G32) );
  NAND2_X2 NAND2_16( .ZN(G314), .A1(G1), .A2(G5) );
  NAND2_X1 NAND2_17( .ZN(G317), .A1(G9), .A2(G13) );
  NAND2_X1 NAND2_18( .ZN(G320), .A1(G2), .A2(G6) );
  NAND2_X1 NAND2_19( .ZN(G323), .A1(G10), .A2(G14) );
  NAND2_X1 NAND2_20( .ZN(G326), .A1(G3), .A2(G7) );
  NAND2_X1 NAND2_21( .ZN(G329), .A1(G11), .A2(G15) );
  NAND2_X1 NAND2_22( .ZN(G332), .A1(G4), .A2(G8) );
  NAND2_X1 NAND2_23( .ZN(G335), .A1(G12), .A2(G16) );
  NAND2_X1 NAND2_24( .ZN(G338), .A1(G17), .A2(G21) );
  NAND2_X1 NAND2_25( .ZN(G341), .A1(G25), .A2(G29) );
  NAND2_X1 NAND2_26( .ZN(G344), .A1(G18), .A2(G22) );
  NAND2_X1 NAND2_27( .ZN(G347), .A1(G26), .A2(G30) );
  NAND2_X1 NAND2_28( .ZN(G350), .A1(G19), .A2(G23) );
  NAND2_X1 NAND2_29( .ZN(G353), .A1(G27), .A2(G31) );
  NAND2_X1 NAND2_30( .ZN(G356), .A1(G20), .A2(G24) );
  NAND2_X1 NAND2_31( .ZN(G359), .A1(G28), .A2(G32) );
  NAND2_X1 NAND2_32( .ZN(G362), .A1(G1), .A2(G266) );
  NAND2_X1 NAND2_33( .ZN(G363), .A1(G2), .A2(G266) );
  NAND2_X1 NAND2_34( .ZN(G364), .A1(G3), .A2(G269) );
  NAND2_X1 NAND2_35( .ZN(G365), .A1(G4), .A2(G269) );
  NAND2_X1 NAND2_36( .ZN(G366), .A1(G5), .A2(G272) );
  NAND2_X1 NAND2_37( .ZN(G367), .A1(G6), .A2(G272) );
  NAND2_X1 NAND2_38( .ZN(G368), .A1(G7), .A2(G275) );
  NAND2_X1 NAND2_39( .ZN(G369), .A1(G8), .A2(G275) );
  NAND2_X1 NAND2_40( .ZN(G370), .A1(G9), .A2(G278) );
  NAND2_X1 NAND2_41( .ZN(G371), .A1(G10), .A2(G278) );
  NAND2_X1 NAND2_42( .ZN(G372), .A1(G11), .A2(G281) );
  NAND2_X1 NAND2_43( .ZN(G373), .A1(G12), .A2(G281) );
  NAND2_X1 NAND2_44( .ZN(G374), .A1(G13), .A2(G284) );
  NAND2_X1 NAND2_45( .ZN(G375), .A1(G14), .A2(G284) );
  NAND2_X1 NAND2_46( .ZN(G376), .A1(G15), .A2(G287) );
  NAND2_X1 NAND2_47( .ZN(G377), .A1(G16), .A2(G287) );
  NAND2_X1 NAND2_48( .ZN(G378), .A1(G17), .A2(G290) );
  NAND2_X1 NAND2_49( .ZN(G379), .A1(G18), .A2(G290) );
  NAND2_X1 NAND2_50( .ZN(G380), .A1(G19), .A2(G293) );
  NAND2_X1 NAND2_51( .ZN(G381), .A1(G20), .A2(G293) );
  NAND2_X1 NAND2_52( .ZN(G382), .A1(G21), .A2(G296) );
  NAND2_X1 NAND2_53( .ZN(G383), .A1(G22), .A2(G296) );
  NAND2_X1 NAND2_54( .ZN(G384), .A1(G23), .A2(G299) );
  NAND2_X1 NAND2_55( .ZN(G385), .A1(G24), .A2(G299) );
  NAND2_X1 NAND2_56( .ZN(G386), .A1(G25), .A2(G302) );
  NAND2_X1 NAND2_57( .ZN(G387), .A1(G26), .A2(G302) );
  NAND2_X1 NAND2_58( .ZN(G388), .A1(G27), .A2(G305) );
  NAND2_X1 NAND2_59( .ZN(G389), .A1(G28), .A2(G305) );
  NAND2_X1 NAND2_60( .ZN(G390), .A1(G29), .A2(G308) );
  NAND2_X1 NAND2_61( .ZN(G391), .A1(G30), .A2(G308) );
  NAND2_X1 NAND2_62( .ZN(G392), .A1(G31), .A2(G311) );
  NAND2_X1 NAND2_63( .ZN(G393), .A1(G32), .A2(G311) );
  NAND2_X1 NAND2_64( .ZN(G394), .A1(G1), .A2(G314) );
  NAND2_X1 NAND2_65( .ZN(G395), .A1(G5), .A2(G314) );
  NAND2_X1 NAND2_66( .ZN(G396), .A1(G9), .A2(G317) );
  NAND2_X1 NAND2_67( .ZN(G397), .A1(G13), .A2(G317) );
  NAND2_X1 NAND2_68( .ZN(G398), .A1(G2), .A2(G320) );
  NAND2_X1 NAND2_69( .ZN(G399), .A1(G6), .A2(G320) );
  NAND2_X1 NAND2_70( .ZN(G400), .A1(G10), .A2(G323) );
  NAND2_X1 NAND2_71( .ZN(G401), .A1(G14), .A2(G323) );
  NAND2_X1 NAND2_72( .ZN(G402), .A1(G3), .A2(G326) );
  NAND2_X1 NAND2_73( .ZN(G403), .A1(G7), .A2(G326) );
  NAND2_X1 NAND2_74( .ZN(G404), .A1(G11), .A2(G329) );
  NAND2_X1 NAND2_75( .ZN(G405), .A1(G15), .A2(G329) );
  NAND2_X1 NAND2_76( .ZN(G406), .A1(G4), .A2(G332) );
  NAND2_X1 NAND2_77( .ZN(G407), .A1(G8), .A2(G332) );
  NAND2_X1 NAND2_78( .ZN(G408), .A1(G12), .A2(G335) );
  NAND2_X1 NAND2_79( .ZN(G409), .A1(G16), .A2(G335) );
  NAND2_X1 NAND2_80( .ZN(G410), .A1(G17), .A2(G338) );
  NAND2_X1 NAND2_81( .ZN(G411), .A1(G21), .A2(G338) );
  NAND2_X1 NAND2_82( .ZN(G412), .A1(G25), .A2(G341) );
  NAND2_X1 NAND2_83( .ZN(G413), .A1(G29), .A2(G341) );
  NAND2_X1 NAND2_84( .ZN(G414), .A1(G18), .A2(G344) );
  NAND2_X1 NAND2_85( .ZN(G415), .A1(G22), .A2(G344) );
  NAND2_X1 NAND2_86( .ZN(G416), .A1(G26), .A2(G347) );
  NAND2_X1 NAND2_87( .ZN(G417), .A1(G30), .A2(G347) );
  NAND2_X1 NAND2_88( .ZN(G418), .A1(G19), .A2(G350) );
  NAND2_X1 NAND2_89( .ZN(G419), .A1(G23), .A2(G350) );
  NAND2_X2 NAND2_90( .ZN(G420), .A1(G27), .A2(G353) );
  NAND2_X2 NAND2_91( .ZN(G421), .A1(G31), .A2(G353) );
  NAND2_X2 NAND2_92( .ZN(G422), .A1(G20), .A2(G356) );
  NAND2_X2 NAND2_93( .ZN(G423), .A1(G24), .A2(G356) );
  NAND2_X2 NAND2_94( .ZN(G424), .A1(G28), .A2(G359) );
  NAND2_X2 NAND2_95( .ZN(G425), .A1(G32), .A2(G359) );
  NAND2_X1 NAND2_96( .ZN(G426), .A1(G362), .A2(G363) );
  NAND2_X1 NAND2_97( .ZN(G429), .A1(G364), .A2(G365) );
  NAND2_X1 NAND2_98( .ZN(G432), .A1(G366), .A2(G367) );
  NAND2_X1 NAND2_99( .ZN(G435), .A1(G368), .A2(G369) );
  NAND2_X1 NAND2_100( .ZN(G438), .A1(G370), .A2(G371) );
  NAND2_X1 NAND2_101( .ZN(G441), .A1(G372), .A2(G373) );
  NAND2_X1 NAND2_102( .ZN(G444), .A1(G374), .A2(G375) );
  NAND2_X1 NAND2_103( .ZN(G447), .A1(G376), .A2(G377) );
  NAND2_X1 NAND2_104( .ZN(G450), .A1(G378), .A2(G379) );
  NAND2_X1 NAND2_105( .ZN(G453), .A1(G380), .A2(G381) );
  NAND2_X1 NAND2_106( .ZN(G456), .A1(G382), .A2(G383) );
  NAND2_X1 NAND2_107( .ZN(G459), .A1(G384), .A2(G385) );
  NAND2_X1 NAND2_108( .ZN(G462), .A1(G386), .A2(G387) );
  NAND2_X1 NAND2_109( .ZN(G465), .A1(G388), .A2(G389) );
  NAND2_X1 NAND2_110( .ZN(G468), .A1(G390), .A2(G391) );
  NAND2_X1 NAND2_111( .ZN(G471), .A1(G392), .A2(G393) );
  NAND2_X1 NAND2_112( .ZN(G474), .A1(G394), .A2(G395) );
  NAND2_X1 NAND2_113( .ZN(G477), .A1(G396), .A2(G397) );
  NAND2_X1 NAND2_114( .ZN(G480), .A1(G398), .A2(G399) );
  NAND2_X1 NAND2_115( .ZN(G483), .A1(G400), .A2(G401) );
  NAND2_X1 NAND2_116( .ZN(G486), .A1(G402), .A2(G403) );
  NAND2_X1 NAND2_117( .ZN(G489), .A1(G404), .A2(G405) );
  NAND2_X1 NAND2_118( .ZN(G492), .A1(G406), .A2(G407) );
  NAND2_X1 NAND2_119( .ZN(G495), .A1(G408), .A2(G409) );
  NAND2_X1 NAND2_120( .ZN(G498), .A1(G410), .A2(G411) );
  NAND2_X1 NAND2_121( .ZN(G501), .A1(G412), .A2(G413) );
  NAND2_X1 NAND2_122( .ZN(G504), .A1(G414), .A2(G415) );
  NAND2_X1 NAND2_123( .ZN(G507), .A1(G416), .A2(G417) );
  NAND2_X1 NAND2_124( .ZN(G510), .A1(G418), .A2(G419) );
  NAND2_X1 NAND2_125( .ZN(G513), .A1(G420), .A2(G421) );
  NAND2_X1 NAND2_126( .ZN(G516), .A1(G422), .A2(G423) );
  NAND2_X1 NAND2_127( .ZN(G519), .A1(G424), .A2(G425) );
  NAND2_X1 NAND2_128( .ZN(G522), .A1(G426), .A2(G429) );
  NAND2_X1 NAND2_129( .ZN(G525), .A1(G432), .A2(G435) );
  NAND2_X1 NAND2_130( .ZN(G528), .A1(G438), .A2(G441) );
  NAND2_X1 NAND2_131( .ZN(G531), .A1(G444), .A2(G447) );
  NAND2_X1 NAND2_132( .ZN(G534), .A1(G450), .A2(G453) );
  NAND2_X1 NAND2_133( .ZN(G537), .A1(G456), .A2(G459) );
  NAND2_X1 NAND2_134( .ZN(G540), .A1(G462), .A2(G465) );
  NAND2_X1 NAND2_135( .ZN(G543), .A1(G468), .A2(G471) );
  NAND2_X1 NAND2_136( .ZN(G546), .A1(G474), .A2(G477) );
  NAND2_X1 NAND2_137( .ZN(G549), .A1(G480), .A2(G483) );
  NAND2_X1 NAND2_138( .ZN(G552), .A1(G486), .A2(G489) );
  NAND2_X1 NAND2_139( .ZN(G555), .A1(G492), .A2(G495) );
  NAND2_X1 NAND2_140( .ZN(G558), .A1(G498), .A2(G501) );
  NAND2_X1 NAND2_141( .ZN(G561), .A1(G504), .A2(G507) );
  NAND2_X1 NAND2_142( .ZN(G564), .A1(G510), .A2(G513) );
  NAND2_X1 NAND2_143( .ZN(G567), .A1(G516), .A2(G519) );
  NAND2_X1 NAND2_144( .ZN(G570), .A1(G426), .A2(G522) );
  NAND2_X1 NAND2_145( .ZN(G571), .A1(G429), .A2(G522) );
  NAND2_X1 NAND2_146( .ZN(G572), .A1(G432), .A2(G525) );
  NAND2_X1 NAND2_147( .ZN(G573), .A1(G435), .A2(G525) );
  NAND2_X1 NAND2_148( .ZN(G574), .A1(G438), .A2(G528) );
  NAND2_X1 NAND2_149( .ZN(G575), .A1(G441), .A2(G528) );
  NAND2_X1 NAND2_150( .ZN(G576), .A1(G444), .A2(G531) );
  NAND2_X1 NAND2_151( .ZN(G577), .A1(G447), .A2(G531) );
  NAND2_X1 NAND2_152( .ZN(G578), .A1(G450), .A2(G534) );
  NAND2_X1 NAND2_153( .ZN(G579), .A1(G453), .A2(G534) );
  NAND2_X1 NAND2_154( .ZN(G580), .A1(G456), .A2(G537) );
  NAND2_X1 NAND2_155( .ZN(G581), .A1(G459), .A2(G537) );
  NAND2_X1 NAND2_156( .ZN(G582), .A1(G462), .A2(G540) );
  NAND2_X1 NAND2_157( .ZN(G583), .A1(G465), .A2(G540) );
  NAND2_X1 NAND2_158( .ZN(G584), .A1(G468), .A2(G543) );
  NAND2_X1 NAND2_159( .ZN(G585), .A1(G471), .A2(G543) );
  NAND2_X1 NAND2_160( .ZN(G586), .A1(G474), .A2(G546) );
  NAND2_X1 NAND2_161( .ZN(G587), .A1(G477), .A2(G546) );
  NAND2_X1 NAND2_162( .ZN(G588), .A1(G480), .A2(G549) );
  NAND2_X1 NAND2_163( .ZN(G589), .A1(G483), .A2(G549) );
  NAND2_X1 NAND2_164( .ZN(G590), .A1(G486), .A2(G552) );
  NAND2_X1 NAND2_165( .ZN(G591), .A1(G489), .A2(G552) );
  NAND2_X1 NAND2_166( .ZN(G592), .A1(G492), .A2(G555) );
  NAND2_X1 NAND2_167( .ZN(G593), .A1(G495), .A2(G555) );
  NAND2_X1 NAND2_168( .ZN(G594), .A1(G498), .A2(G558) );
  NAND2_X1 NAND2_169( .ZN(G595), .A1(G501), .A2(G558) );
  NAND2_X1 NAND2_170( .ZN(G596), .A1(G504), .A2(G561) );
  NAND2_X1 NAND2_171( .ZN(G597), .A1(G507), .A2(G561) );
  NAND2_X1 NAND2_172( .ZN(G598), .A1(G510), .A2(G564) );
  NAND2_X1 NAND2_173( .ZN(G599), .A1(G513), .A2(G564) );
  NAND2_X1 NAND2_174( .ZN(G600), .A1(G516), .A2(G567) );
  NAND2_X1 NAND2_175( .ZN(G601), .A1(G519), .A2(G567) );
  NAND2_X1 NAND2_176( .ZN(G602), .A1(G570), .A2(G571) );
  NAND2_X1 NAND2_177( .ZN(G607), .A1(G572), .A2(G573) );
  NAND2_X1 NAND2_178( .ZN(G612), .A1(G574), .A2(G575) );
  NAND2_X1 NAND2_179( .ZN(G617), .A1(G576), .A2(G577) );
  NAND2_X1 NAND2_180( .ZN(G622), .A1(G578), .A2(G579) );
  NAND2_X1 NAND2_181( .ZN(G627), .A1(G580), .A2(G581) );
  NAND2_X1 NAND2_182( .ZN(G632), .A1(G582), .A2(G583) );
  NAND2_X1 NAND2_183( .ZN(G637), .A1(G584), .A2(G585) );
  NAND2_X1 NAND2_184( .ZN(G642), .A1(G586), .A2(G587) );
  NAND2_X1 NAND2_185( .ZN(G645), .A1(G588), .A2(G589) );
  NAND2_X1 NAND2_186( .ZN(G648), .A1(G590), .A2(G591) );
  NAND2_X1 NAND2_187( .ZN(G651), .A1(G592), .A2(G593) );
  NAND2_X1 NAND2_188( .ZN(G654), .A1(G594), .A2(G595) );
  NAND2_X1 NAND2_189( .ZN(G657), .A1(G596), .A2(G597) );
  NAND2_X1 NAND2_190( .ZN(G660), .A1(G598), .A2(G599) );
  NAND2_X1 NAND2_191( .ZN(G663), .A1(G600), .A2(G601) );
  NAND2_X1 NAND2_192( .ZN(G666), .A1(G602), .A2(G607) );
  NAND2_X1 NAND2_193( .ZN(G669), .A1(G612), .A2(G617) );
  NAND2_X1 NAND2_194( .ZN(G672), .A1(G602), .A2(G612) );
  NAND2_X1 NAND2_195( .ZN(G675), .A1(G607), .A2(G617) );
  NAND2_X1 NAND2_196( .ZN(G678), .A1(G622), .A2(G627) );
  NAND2_X1 NAND2_197( .ZN(G681), .A1(G632), .A2(G637) );
  NAND2_X1 NAND2_198( .ZN(G684), .A1(G622), .A2(G632) );
  NAND2_X1 NAND2_199( .ZN(G687), .A1(G627), .A2(G637) );
  NAND2_X1 NAND2_200( .ZN(G690), .A1(G602), .A2(G666) );
  NAND2_X1 NAND2_201( .ZN(G691), .A1(G607), .A2(G666) );
  NAND2_X1 NAND2_202( .ZN(G692), .A1(G612), .A2(G669) );
  NAND2_X1 NAND2_203( .ZN(G693), .A1(G617), .A2(G669) );
  NAND2_X1 NAND2_204( .ZN(G694), .A1(G602), .A2(G672) );
  NAND2_X1 NAND2_205( .ZN(G695), .A1(G612), .A2(G672) );
  NAND2_X1 NAND2_206( .ZN(G696), .A1(G607), .A2(G675) );
  NAND2_X1 NAND2_207( .ZN(G697), .A1(G617), .A2(G675) );
  NAND2_X1 NAND2_208( .ZN(G698), .A1(G622), .A2(G678) );
  NAND2_X1 NAND2_209( .ZN(G699), .A1(G627), .A2(G678) );
  NAND2_X1 NAND2_210( .ZN(G700), .A1(G632), .A2(G681) );
  NAND2_X1 NAND2_211( .ZN(G701), .A1(G637), .A2(G681) );
  NAND2_X1 NAND2_212( .ZN(G702), .A1(G622), .A2(G684) );
  NAND2_X1 NAND2_213( .ZN(G703), .A1(G632), .A2(G684) );
  NAND2_X1 NAND2_214( .ZN(G704), .A1(G627), .A2(G687) );
  NAND2_X1 NAND2_215( .ZN(G705), .A1(G637), .A2(G687) );
  NAND2_X1 NAND2_216( .ZN(G706), .A1(G690), .A2(G691) );
  NAND2_X1 NAND2_217( .ZN(G709), .A1(G692), .A2(G693) );
  NAND2_X1 NAND2_218( .ZN(G712), .A1(G694), .A2(G695) );
  NAND2_X1 NAND2_219( .ZN(G715), .A1(G696), .A2(G697) );
  NAND2_X1 NAND2_220( .ZN(G718), .A1(G698), .A2(G699) );
  NAND2_X1 NAND2_221( .ZN(G721), .A1(G700), .A2(G701) );
  NAND2_X1 NAND2_222( .ZN(G724), .A1(G702), .A2(G703) );
  NAND2_X1 NAND2_223( .ZN(G727), .A1(G704), .A2(G705) );
  NAND2_X1 NAND2_224( .ZN(G730), .A1(G242), .A2(G718) );
  NAND2_X1 NAND2_225( .ZN(G733), .A1(G245), .A2(G721) );
  NAND2_X1 NAND2_226( .ZN(G736), .A1(G248), .A2(G724) );
  NAND2_X1 NAND2_227( .ZN(G739), .A1(G251), .A2(G727) );
  NAND2_X1 NAND2_228( .ZN(G742), .A1(G254), .A2(G706) );
  NAND2_X1 NAND2_229( .ZN(G745), .A1(G257), .A2(G709) );
  NAND2_X1 NAND2_230( .ZN(G748), .A1(G260), .A2(G712) );
  NAND2_X1 NAND2_231( .ZN(G751), .A1(G263), .A2(G715) );
  NAND2_X1 NAND2_232( .ZN(G754), .A1(G242), .A2(G730) );
  NAND2_X1 NAND2_233( .ZN(G755), .A1(G718), .A2(G730) );
  NAND2_X1 NAND2_234( .ZN(G756), .A1(G245), .A2(G733) );
  NAND2_X1 NAND2_235( .ZN(G757), .A1(G721), .A2(G733) );
  NAND2_X1 NAND2_236( .ZN(G758), .A1(G248), .A2(G736) );
  NAND2_X1 NAND2_237( .ZN(G759), .A1(G724), .A2(G736) );
  NAND2_X1 NAND2_238( .ZN(G760), .A1(G251), .A2(G739) );
  NAND2_X1 NAND2_239( .ZN(G761), .A1(G727), .A2(G739) );
  NAND2_X1 NAND2_240( .ZN(G762), .A1(G254), .A2(G742) );
  NAND2_X1 NAND2_241( .ZN(G763), .A1(G706), .A2(G742) );
  NAND2_X1 NAND2_242( .ZN(G764), .A1(G257), .A2(G745) );
  NAND2_X1 NAND2_243( .ZN(G765), .A1(G709), .A2(G745) );
  NAND2_X1 NAND2_244( .ZN(G766), .A1(G260), .A2(G748) );
  NAND2_X1 NAND2_245( .ZN(G767), .A1(G712), .A2(G748) );
  NAND2_X1 NAND2_246( .ZN(G768), .A1(G263), .A2(G751) );
  NAND2_X1 NAND2_247( .ZN(G769), .A1(G715), .A2(G751) );
  NAND2_X1 NAND2_248( .ZN(G770), .A1(G754), .A2(G755) );
  NAND2_X1 NAND2_249( .ZN(G773), .A1(G756), .A2(G757) );
  NAND2_X1 NAND2_250( .ZN(G776), .A1(G758), .A2(G759) );
  NAND2_X1 NAND2_251( .ZN(G779), .A1(G760), .A2(G761) );
  NAND2_X1 NAND2_252( .ZN(G782), .A1(G762), .A2(G763) );
  NAND2_X1 NAND2_253( .ZN(G785), .A1(G764), .A2(G765) );
  NAND2_X1 NAND2_254( .ZN(G788), .A1(G766), .A2(G767) );
  NAND2_X1 NAND2_255( .ZN(G791), .A1(G768), .A2(G769) );
  NAND2_X1 NAND2_256( .ZN(G794), .A1(G642), .A2(G770) );
  NAND2_X1 NAND2_257( .ZN(G797), .A1(G645), .A2(G773) );
  NAND2_X1 NAND2_258( .ZN(G800), .A1(G648), .A2(G776) );
  NAND2_X1 NAND2_259( .ZN(G803), .A1(G651), .A2(G779) );
  NAND2_X1 NAND2_260( .ZN(G806), .A1(G654), .A2(G782) );
  NAND2_X1 NAND2_261( .ZN(G809), .A1(G657), .A2(G785) );
  NAND2_X1 NAND2_262( .ZN(G812), .A1(G660), .A2(G788) );
  NAND2_X1 NAND2_263( .ZN(G815), .A1(G663), .A2(G791) );
  NAND2_X1 NAND2_264( .ZN(G818), .A1(G642), .A2(G794) );
  NAND2_X1 NAND2_265( .ZN(G819), .A1(G770), .A2(G794) );
  NAND2_X1 NAND2_266( .ZN(G820), .A1(G645), .A2(G797) );
  NAND2_X1 NAND2_267( .ZN(G821), .A1(G773), .A2(G797) );
  NAND2_X1 NAND2_268( .ZN(G822), .A1(G648), .A2(G800) );
  NAND2_X1 NAND2_269( .ZN(G823), .A1(G776), .A2(G800) );
  NAND2_X1 NAND2_270( .ZN(G824), .A1(G651), .A2(G803) );
  NAND2_X1 NAND2_271( .ZN(G825), .A1(G779), .A2(G803) );
  NAND2_X2 NAND2_272( .ZN(G826), .A1(G654), .A2(G806) );
  NAND2_X2 NAND2_273( .ZN(G827), .A1(G782), .A2(G806) );
  NAND2_X2 NAND2_274( .ZN(G828), .A1(G657), .A2(G809) );
  NAND2_X2 NAND2_275( .ZN(G829), .A1(G785), .A2(G809) );
  NAND2_X2 NAND2_276( .ZN(G830), .A1(G660), .A2(G812) );
  NAND2_X2 NAND2_277( .ZN(G831), .A1(G788), .A2(G812) );
  NAND2_X2 NAND2_278( .ZN(G832), .A1(G663), .A2(G815) );
  NAND2_X1 NAND2_279( .ZN(G833), .A1(G791), .A2(G815) );
  NAND2_X1 NAND2_280( .ZN(G834), .A1(G818), .A2(G819) );
  NAND2_X1 NAND2_281( .ZN(G847), .A1(G820), .A2(G821) );
  NAND2_X1 NAND2_282( .ZN(G860), .A1(G822), .A2(G823) );
  NAND2_X1 NAND2_283( .ZN(G873), .A1(G824), .A2(G825) );
  NAND2_X1 NAND2_284( .ZN(G886), .A1(G828), .A2(G829) );
  NAND2_X1 NAND2_285( .ZN(G899), .A1(G832), .A2(G833) );
  NAND2_X1 NAND2_286( .ZN(G912), .A1(G830), .A2(G831) );
  NAND2_X1 NAND2_287( .ZN(G925), .A1(G826), .A2(G827) );
  INV_X1 NOT_0( .ZN(G938), .A(G834) );
  INV_X1 NOT_1( .ZN(G939), .A(G847) );
  INV_X4 NOT_2( .ZN(G940), .A(G860) );
  INV_X4 NOT_3( .ZN(G941), .A(G834) );
  INV_X4 NOT_4( .ZN(G942), .A(G847) );
  INV_X4 NOT_5( .ZN(G943), .A(G873) );
  INV_X1 NOT_6( .ZN(G944), .A(G834) );
  INV_X1 NOT_7( .ZN(G945), .A(G860) );
  INV_X1 NOT_8( .ZN(G946), .A(G873) );
  INV_X1 NOT_9( .ZN(G947), .A(G847) );
  INV_X1 NOT_10( .ZN(G948), .A(G860) );
  INV_X1 NOT_11( .ZN(G949), .A(G873) );
  INV_X1 NOT_12( .ZN(G950), .A(G886) );
  INV_X1 NOT_13( .ZN(G951), .A(G899) );
  INV_X1 NOT_14( .ZN(G952), .A(G886) );
  INV_X1 NOT_15( .ZN(G953), .A(G912) );
  INV_X1 NOT_16( .ZN(G954), .A(G925) );
  INV_X1 NOT_17( .ZN(G955), .A(G899) );
  INV_X1 NOT_18( .ZN(G956), .A(G925) );
  INV_X1 NOT_19( .ZN(G957), .A(G912) );
  INV_X1 NOT_20( .ZN(G958), .A(G925) );
  INV_X1 NOT_21( .ZN(G959), .A(G886) );
  INV_X1 NOT_22( .ZN(G960), .A(G912) );
  INV_X1 NOT_23( .ZN(G961), .A(G925) );
  INV_X1 NOT_24( .ZN(G962), .A(G886) );
  INV_X1 NOT_25( .ZN(G963), .A(G899) );
  INV_X1 NOT_26( .ZN(G964), .A(G925) );
  INV_X1 NOT_27( .ZN(G965), .A(G912) );
  INV_X1 NOT_28( .ZN(G966), .A(G899) );
  INV_X1 NOT_29( .ZN(G967), .A(G886) );
  INV_X1 NOT_30( .ZN(G968), .A(G912) );
  INV_X1 NOT_31( .ZN(G969), .A(G899) );
  INV_X1 NOT_32( .ZN(G970), .A(G847) );
  INV_X4 NOT_33( .ZN(G971), .A(G873) );
  INV_X4 NOT_34( .ZN(G972), .A(G847) );
  INV_X4 NOT_35( .ZN(G973), .A(G860) );
  INV_X1 NOT_36( .ZN(G974), .A(G834) );
  INV_X1 NOT_37( .ZN(G975), .A(G873) );
  INV_X1 NOT_38( .ZN(G976), .A(G834) );
  INV_X1 NOT_39( .ZN(G977), .A(G860) );
  AND4_X1 AND4_0( .ZN(G978), .A1(G938), .A2(G939), .A3(G940), .A4(G873) );
  AND4_X1 AND4_1( .ZN(G979), .A1(G941), .A2(G942), .A3(G860), .A4(G943) );
  AND4_X1 AND4_2( .ZN(G980), .A1(G944), .A2(G847), .A3(G945), .A4(G946) );
  AND4_X1 AND4_3( .ZN(G981), .A1(G834), .A2(G947), .A3(G948), .A4(G949) );
  AND4_X1 AND4_4( .ZN(G982), .A1(G958), .A2(G959), .A3(G960), .A4(G899) );
  AND4_X1 AND4_5( .ZN(G983), .A1(G961), .A2(G962), .A3(G912), .A4(G963) );
  AND4_X1 AND4_6( .ZN(G984), .A1(G964), .A2(G886), .A3(G965), .A4(G966) );
  AND4_X1 AND4_7( .ZN(G985), .A1(G925), .A2(G967), .A3(G968), .A4(G969) );
  OR4_X1 OR4_0( .ZN(G986), .A1(G978), .A2(G979), .A3(G980), .A4(G981) );
  OR4_X1 OR4_1( .ZN(G991), .A1(G982), .A2(G983), .A3(G984), .A4(G985) );
  AND4_X1 AND5_0_A( .ZN(extra0), .A1(G925), .A2(G950), .A3(G912), .A4(G951) );
  AND2_X1 AND5_0( .ZN(G996), .A1(extra0), .A2(G986) );
  AND4_X1 AND5_1_A( .ZN(extra1), .A1(G925), .A2(G952), .A3(G953), .A4(G899) );
  AND2_X1 AND5_1( .ZN(G1001), .A1(extra1), .A2(G986) );
  AND4_X1 AND5_2_A( .ZN(extra2), .A1(G954), .A2(G886), .A3(G912), .A4(G955) );
  AND2_X1 AND5_2( .ZN(G1006), .A1(extra2), .A2(G986) );
  AND4_X1 AND5_3_A( .ZN(extra3), .A1(G956), .A2(G886), .A3(G957), .A4(G899) );
  AND2_X1 AND5_3( .ZN(G1011), .A1(extra3), .A2(G986) );
  AND4_X1 AND5_4_A( .ZN(extra4), .A1(G834), .A2(G970), .A3(G860), .A4(G971) );
  AND2_X1 AND5_4( .ZN(G1016), .A1(extra4), .A2(G991) );
  AND4_X1 AND5_5_A( .ZN(extra5), .A1(G834), .A2(G972), .A3(G973), .A4(G873) );
  AND2_X1 AND5_5( .ZN(G1021), .A1(extra5), .A2(G991) );
  AND4_X1 AND5_6_A( .ZN(extra6), .A1(G974), .A2(G847), .A3(G860), .A4(G975) );
  AND2_X1 AND5_6( .ZN(G1026), .A1(extra6), .A2(G991) );
  AND4_X1 AND5_7_A( .ZN(extra7), .A1(G976), .A2(G847), .A3(G977), .A4(G873) );
  AND2_X1 AND5_7( .ZN(G1031), .A1(extra7), .A2(G991) );
  AND2_X1 AND2_8( .ZN(G1036), .A1(G834), .A2(G996) );
  AND2_X1 AND2_9( .ZN(G1039), .A1(G847), .A2(G996) );
  AND2_X4 AND2_10( .ZN(G1042), .A1(G860), .A2(G996) );
  AND2_X4 AND2_11( .ZN(G1045), .A1(G873), .A2(G996) );
  AND2_X1 AND2_12( .ZN(G1048), .A1(G834), .A2(G1001) );
  AND2_X1 AND2_13( .ZN(G1051), .A1(G847), .A2(G1001) );
  AND2_X1 AND2_14( .ZN(G1054), .A1(G860), .A2(G1001) );
  AND2_X1 AND2_15( .ZN(G1057), .A1(G873), .A2(G1001) );
  AND2_X1 AND2_16( .ZN(G1060), .A1(G834), .A2(G1006) );
  AND2_X1 AND2_17( .ZN(G1063), .A1(G847), .A2(G1006) );
  AND2_X1 AND2_18( .ZN(G1066), .A1(G860), .A2(G1006) );
  AND2_X1 AND2_19( .ZN(G1069), .A1(G873), .A2(G1006) );
  AND2_X1 AND2_20( .ZN(G1072), .A1(G834), .A2(G1011) );
  AND2_X1 AND2_21( .ZN(G1075), .A1(G847), .A2(G1011) );
  AND2_X1 AND2_22( .ZN(G1078), .A1(G860), .A2(G1011) );
  AND2_X1 AND2_23( .ZN(G1081), .A1(G873), .A2(G1011) );
  AND2_X1 AND2_24( .ZN(G1084), .A1(G925), .A2(G1016) );
  AND2_X1 AND2_25( .ZN(G1087), .A1(G886), .A2(G1016) );
  AND2_X1 AND2_26( .ZN(G1090), .A1(G912), .A2(G1016) );
  AND2_X1 AND2_27( .ZN(G1093), .A1(G899), .A2(G1016) );
  AND2_X1 AND2_28( .ZN(G1096), .A1(G925), .A2(G1021) );
  AND2_X1 AND2_29( .ZN(G1099), .A1(G886), .A2(G1021) );
  AND2_X1 AND2_30( .ZN(G1102), .A1(G912), .A2(G1021) );
  AND2_X1 AND2_31( .ZN(G1105), .A1(G899), .A2(G1021) );
  AND2_X4 AND2_32( .ZN(G1108), .A1(G925), .A2(G1026) );
  AND2_X4 AND2_33( .ZN(G1111), .A1(G886), .A2(G1026) );
  AND2_X4 AND2_34( .ZN(G1114), .A1(G912), .A2(G1026) );
  AND2_X4 AND2_35( .ZN(G1117), .A1(G899), .A2(G1026) );
  AND2_X1 AND2_36( .ZN(G1120), .A1(G925), .A2(G1031) );
  AND2_X1 AND2_37( .ZN(G1123), .A1(G886), .A2(G1031) );
  AND2_X1 AND2_38( .ZN(G1126), .A1(G912), .A2(G1031) );
  AND2_X1 AND2_39( .ZN(G1129), .A1(G899), .A2(G1031) );
  NAND2_X1 NAND2_288( .ZN(G1132), .A1(G1), .A2(G1036) );
  NAND2_X1 NAND2_289( .ZN(G1135), .A1(G2), .A2(G1039) );
  NAND2_X1 NAND2_290( .ZN(G1138), .A1(G3), .A2(G1042) );
  NAND2_X1 NAND2_291( .ZN(G1141), .A1(G4), .A2(G1045) );
  NAND2_X1 NAND2_292( .ZN(G1144), .A1(G5), .A2(G1048) );
  NAND2_X1 NAND2_293( .ZN(G1147), .A1(G6), .A2(G1051) );
  NAND2_X1 NAND2_294( .ZN(G1150), .A1(G7), .A2(G1054) );
  NAND2_X1 NAND2_295( .ZN(G1153), .A1(G8), .A2(G1057) );
  NAND2_X1 NAND2_296( .ZN(G1156), .A1(G9), .A2(G1060) );
  NAND2_X1 NAND2_297( .ZN(G1159), .A1(G10), .A2(G1063) );
  NAND2_X1 NAND2_298( .ZN(G1162), .A1(G11), .A2(G1066) );
  NAND2_X1 NAND2_299( .ZN(G1165), .A1(G12), .A2(G1069) );
  NAND2_X1 NAND2_300( .ZN(G1168), .A1(G13), .A2(G1072) );
  NAND2_X1 NAND2_301( .ZN(G1171), .A1(G14), .A2(G1075) );
  NAND2_X1 NAND2_302( .ZN(G1174), .A1(G15), .A2(G1078) );
  NAND2_X1 NAND2_303( .ZN(G1177), .A1(G16), .A2(G1081) );
  NAND2_X1 NAND2_304( .ZN(G1180), .A1(G17), .A2(G1084) );
  NAND2_X1 NAND2_305( .ZN(G1183), .A1(G18), .A2(G1087) );
  NAND2_X1 NAND2_306( .ZN(G1186), .A1(G19), .A2(G1090) );
  NAND2_X1 NAND2_307( .ZN(G1189), .A1(G20), .A2(G1093) );
  NAND2_X1 NAND2_308( .ZN(G1192), .A1(G21), .A2(G1096) );
  NAND2_X1 NAND2_309( .ZN(G1195), .A1(G22), .A2(G1099) );
  NAND2_X1 NAND2_310( .ZN(G1198), .A1(G23), .A2(G1102) );
  NAND2_X1 NAND2_311( .ZN(G1201), .A1(G24), .A2(G1105) );
  NAND2_X1 NAND2_312( .ZN(G1204), .A1(G25), .A2(G1108) );
  NAND2_X1 NAND2_313( .ZN(G1207), .A1(G26), .A2(G1111) );
  NAND2_X1 NAND2_314( .ZN(G1210), .A1(G27), .A2(G1114) );
  NAND2_X1 NAND2_315( .ZN(G1213), .A1(G28), .A2(G1117) );
  NAND2_X1 NAND2_316( .ZN(G1216), .A1(G29), .A2(G1120) );
  NAND2_X1 NAND2_317( .ZN(G1219), .A1(G30), .A2(G1123) );
  NAND2_X1 NAND2_318( .ZN(G1222), .A1(G31), .A2(G1126) );
  NAND2_X1 NAND2_319( .ZN(G1225), .A1(G32), .A2(G1129) );
  NAND2_X1 NAND2_320( .ZN(G1228), .A1(G1), .A2(G1132) );
  NAND2_X1 NAND2_321( .ZN(G1229), .A1(G1036), .A2(G1132) );
  NAND2_X1 NAND2_322( .ZN(G1230), .A1(G2), .A2(G1135) );
  NAND2_X1 NAND2_323( .ZN(G1231), .A1(G1039), .A2(G1135) );
  NAND2_X1 NAND2_324( .ZN(G1232), .A1(G3), .A2(G1138) );
  NAND2_X1 NAND2_325( .ZN(G1233), .A1(G1042), .A2(G1138) );
  NAND2_X1 NAND2_326( .ZN(G1234), .A1(G4), .A2(G1141) );
  NAND2_X1 NAND2_327( .ZN(G1235), .A1(G1045), .A2(G1141) );
  NAND2_X1 NAND2_328( .ZN(G1236), .A1(G5), .A2(G1144) );
  NAND2_X1 NAND2_329( .ZN(G1237), .A1(G1048), .A2(G1144) );
  NAND2_X1 NAND2_330( .ZN(G1238), .A1(G6), .A2(G1147) );
  NAND2_X1 NAND2_331( .ZN(G1239), .A1(G1051), .A2(G1147) );
  NAND2_X1 NAND2_332( .ZN(G1240), .A1(G7), .A2(G1150) );
  NAND2_X1 NAND2_333( .ZN(G1241), .A1(G1054), .A2(G1150) );
  NAND2_X1 NAND2_334( .ZN(G1242), .A1(G8), .A2(G1153) );
  NAND2_X1 NAND2_335( .ZN(G1243), .A1(G1057), .A2(G1153) );
  NAND2_X1 NAND2_336( .ZN(G1244), .A1(G9), .A2(G1156) );
  NAND2_X1 NAND2_337( .ZN(G1245), .A1(G1060), .A2(G1156) );
  NAND2_X1 NAND2_338( .ZN(G1246), .A1(G10), .A2(G1159) );
  NAND2_X1 NAND2_339( .ZN(G1247), .A1(G1063), .A2(G1159) );
  NAND2_X1 NAND2_340( .ZN(G1248), .A1(G11), .A2(G1162) );
  NAND2_X1 NAND2_341( .ZN(G1249), .A1(G1066), .A2(G1162) );
  NAND2_X1 NAND2_342( .ZN(G1250), .A1(G12), .A2(G1165) );
  NAND2_X1 NAND2_343( .ZN(G1251), .A1(G1069), .A2(G1165) );
  NAND2_X1 NAND2_344( .ZN(G1252), .A1(G13), .A2(G1168) );
  NAND2_X1 NAND2_345( .ZN(G1253), .A1(G1072), .A2(G1168) );
  NAND2_X1 NAND2_346( .ZN(G1254), .A1(G14), .A2(G1171) );
  NAND2_X1 NAND2_347( .ZN(G1255), .A1(G1075), .A2(G1171) );
  NAND2_X1 NAND2_348( .ZN(G1256), .A1(G15), .A2(G1174) );
  NAND2_X1 NAND2_349( .ZN(G1257), .A1(G1078), .A2(G1174) );
  NAND2_X1 NAND2_350( .ZN(G1258), .A1(G16), .A2(G1177) );
  NAND2_X1 NAND2_351( .ZN(G1259), .A1(G1081), .A2(G1177) );
  NAND2_X1 NAND2_352( .ZN(G1260), .A1(G17), .A2(G1180) );
  NAND2_X1 NAND2_353( .ZN(G1261), .A1(G1084), .A2(G1180) );
  NAND2_X1 NAND2_354( .ZN(G1262), .A1(G18), .A2(G1183) );
  NAND2_X1 NAND2_355( .ZN(G1263), .A1(G1087), .A2(G1183) );
  NAND2_X1 NAND2_356( .ZN(G1264), .A1(G19), .A2(G1186) );
  NAND2_X1 NAND2_357( .ZN(G1265), .A1(G1090), .A2(G1186) );
  NAND2_X1 NAND2_358( .ZN(G1266), .A1(G20), .A2(G1189) );
  NAND2_X1 NAND2_359( .ZN(G1267), .A1(G1093), .A2(G1189) );
  NAND2_X1 NAND2_360( .ZN(G1268), .A1(G21), .A2(G1192) );
  NAND2_X1 NAND2_361( .ZN(G1269), .A1(G1096), .A2(G1192) );
  NAND2_X1 NAND2_362( .ZN(G1270), .A1(G22), .A2(G1195) );
  NAND2_X1 NAND2_363( .ZN(G1271), .A1(G1099), .A2(G1195) );
  NAND2_X1 NAND2_364( .ZN(G1272), .A1(G23), .A2(G1198) );
  NAND2_X1 NAND2_365( .ZN(G1273), .A1(G1102), .A2(G1198) );
  NAND2_X1 NAND2_366( .ZN(G1274), .A1(G24), .A2(G1201) );
  NAND2_X1 NAND2_367( .ZN(G1275), .A1(G1105), .A2(G1201) );
  NAND2_X1 NAND2_368( .ZN(G1276), .A1(G25), .A2(G1204) );
  NAND2_X1 NAND2_369( .ZN(G1277), .A1(G1108), .A2(G1204) );
  NAND2_X1 NAND2_370( .ZN(G1278), .A1(G26), .A2(G1207) );
  NAND2_X1 NAND2_371( .ZN(G1279), .A1(G1111), .A2(G1207) );
  NAND2_X1 NAND2_372( .ZN(G1280), .A1(G27), .A2(G1210) );
  NAND2_X1 NAND2_373( .ZN(G1281), .A1(G1114), .A2(G1210) );
  NAND2_X1 NAND2_374( .ZN(G1282), .A1(G28), .A2(G1213) );
  NAND2_X1 NAND2_375( .ZN(G1283), .A1(G1117), .A2(G1213) );
  NAND2_X1 NAND2_376( .ZN(G1284), .A1(G29), .A2(G1216) );
  NAND2_X1 NAND2_377( .ZN(G1285), .A1(G1120), .A2(G1216) );
  NAND2_X1 NAND2_378( .ZN(G1286), .A1(G30), .A2(G1219) );
  NAND2_X1 NAND2_379( .ZN(G1287), .A1(G1123), .A2(G1219) );
  NAND2_X1 NAND2_380( .ZN(G1288), .A1(G31), .A2(G1222) );
  NAND2_X1 NAND2_381( .ZN(G1289), .A1(G1126), .A2(G1222) );
  NAND2_X1 NAND2_382( .ZN(G1290), .A1(G32), .A2(G1225) );
  NAND2_X1 NAND2_383( .ZN(G1291), .A1(G1129), .A2(G1225) );
  NAND2_X1 NAND2_384( .ZN(G1292), .A1(G1228), .A2(G1229) );
  NAND2_X1 NAND2_385( .ZN(G1293), .A1(G1230), .A2(G1231) );
  NAND2_X1 NAND2_386( .ZN(G1294), .A1(G1232), .A2(G1233) );
  NAND2_X1 NAND2_387( .ZN(G1295), .A1(G1234), .A2(G1235) );
  NAND2_X1 NAND2_388( .ZN(G1296), .A1(G1236), .A2(G1237) );
  NAND2_X1 NAND2_389( .ZN(G1297), .A1(G1238), .A2(G1239) );
  NAND2_X1 NAND2_390( .ZN(G1298), .A1(G1240), .A2(G1241) );
  NAND2_X1 NAND2_391( .ZN(G1299), .A1(G1242), .A2(G1243) );
  NAND2_X2 NAND2_392( .ZN(G1300), .A1(G1244), .A2(G1245) );
  NAND2_X2 NAND2_393( .ZN(G1301), .A1(G1246), .A2(G1247) );
  NAND2_X2 NAND2_394( .ZN(G1302), .A1(G1248), .A2(G1249) );
  NAND2_X2 NAND2_395( .ZN(G1303), .A1(G1250), .A2(G1251) );
  NAND2_X2 NAND2_396( .ZN(G1304), .A1(G1252), .A2(G1253) );
  NAND2_X1 NAND2_397( .ZN(G1305), .A1(G1254), .A2(G1255) );
  NAND2_X1 NAND2_398( .ZN(G1306), .A1(G1256), .A2(G1257) );
  NAND2_X1 NAND2_399( .ZN(G1307), .A1(G1258), .A2(G1259) );
  NAND2_X1 NAND2_400( .ZN(G1308), .A1(G1260), .A2(G1261) );
  NAND2_X1 NAND2_401( .ZN(G1309), .A1(G1262), .A2(G1263) );
  NAND2_X1 NAND2_402( .ZN(G1310), .A1(G1264), .A2(G1265) );
  NAND2_X1 NAND2_403( .ZN(G1311), .A1(G1266), .A2(G1267) );
  NAND2_X1 NAND2_404( .ZN(G1312), .A1(G1268), .A2(G1269) );
  NAND2_X1 NAND2_405( .ZN(G1313), .A1(G1270), .A2(G1271) );
  NAND2_X1 NAND2_406( .ZN(G1314), .A1(G1272), .A2(G1273) );
  NAND2_X1 NAND2_407( .ZN(G1315), .A1(G1274), .A2(G1275) );
  NAND2_X1 NAND2_408( .ZN(G1316), .A1(G1276), .A2(G1277) );
  NAND2_X1 NAND2_409( .ZN(G1317), .A1(G1278), .A2(G1279) );
  NAND2_X1 NAND2_410( .ZN(G1318), .A1(G1280), .A2(G1281) );
  NAND2_X1 NAND2_411( .ZN(G1319), .A1(G1282), .A2(G1283) );
  NAND2_X1 NAND2_412( .ZN(G1320), .A1(G1284), .A2(G1285) );
  NAND2_X1 NAND2_413( .ZN(G1321), .A1(G1286), .A2(G1287) );
  NAND2_X1 NAND2_414( .ZN(G1322), .A1(G1288), .A2(G1289) );
  NAND2_X1 NAND2_415( .ZN(G1323), .A1(G1290), .A2(G1291) );
  INV_X1 NOT_40( .ZN(G1324), .A(G1292) );
  INV_X1 NOT_41( .ZN(G1325), .A(G1293) );
  INV_X32 NOT_42( .ZN(G1326), .A(G1294) );
  INV_X32 NOT_43( .ZN(G1327), .A(G1295) );
  INV_X32 NOT_44( .ZN(G1328), .A(G1296) );
  INV_X32 NOT_45( .ZN(G1329), .A(G1297) );
  INV_X32 NOT_46( .ZN(G1330), .A(G1298) );
  INV_X1 NOT_47( .ZN(G1331), .A(G1299) );
  INV_X1 NOT_48( .ZN(G1332), .A(G1300) );
  INV_X1 NOT_49( .ZN(G1333), .A(G1301) );
  INV_X1 NOT_50( .ZN(G1334), .A(G1302) );
  INV_X1 NOT_51( .ZN(G1335), .A(G1303) );
  INV_X1 NOT_52( .ZN(G1336), .A(G1304) );
  INV_X8 NOT_53( .ZN(G1337), .A(G1305) );
  INV_X8 NOT_54( .ZN(G1338), .A(G1306) );
  INV_X8 NOT_55( .ZN(G1339), .A(G1307) );
  INV_X8 NOT_56( .ZN(G1340), .A(G1308) );
  INV_X1 NOT_57( .ZN(G1341), .A(G1309) );
  INV_X1 NOT_58( .ZN(G1342), .A(G1310) );
  INV_X1 NOT_59( .ZN(G1343), .A(G1311) );
  INV_X1 NOT_60( .ZN(G1344), .A(G1312) );
  INV_X1 NOT_61( .ZN(G1345), .A(G1313) );
  INV_X1 NOT_62( .ZN(G1346), .A(G1314) );
  INV_X1 NOT_63( .ZN(G1347), .A(G1315) );
  INV_X1 NOT_64( .ZN(G1348), .A(G1316) );
  INV_X1 NOT_65( .ZN(G1349), .A(G1317) );
  INV_X1 NOT_66( .ZN(G1350), .A(G1318) );
  INV_X1 NOT_67( .ZN(G1351), .A(G1319) );
  INV_X1 NOT_68( .ZN(G1352), .A(G1320) );
  INV_X4 NOT_69( .ZN(G1353), .A(G1321) );
  INV_X1 NOT_70( .ZN(G1354), .A(G1322) );
  INV_X1 NOT_71( .ZN(G1355), .A(G1323) );

endmodule
