//# 18 inputs
//# 1 outputs
//# 16 D-type flipflops
//# 78 inverters
//# 140 gates (49 ANDs + 29 NANDs + 28 ORs + 34 NORs)

module s420(CK,C_0,C_1,C_10,C_11,C_12,C_13,C_14,C_15,C_16,C_2,C_3,C_4,C_5,C_6,C_7,
  C_8,C_9,P_0,Z);
input CK,P_0,C_16,C_15,C_14,C_13,C_12,C_11,C_10,C_9,C_8,C_7,C_6,C_5,C_4,C_3,C_2,C_1,
  C_0;
output Z;

  wire X_4,I12,X_3,I13,X_2,I14,X_1,I15,X_8,I110,X_7,I111,X_6,I112,X_5,I113,
    X_12,I208,X_11,I209,X_10,I210,X_9,I211,X_16,I306,X_15,I307,X_14,I308,X_13,I309,
    I73_1,I69,I73_2,I7_1,I66,I7_2,I88_1,I88_2,I48,I49,I50,I68,I171_1,I167,I171_2,I105_1,
    I164,I105_2,I186_1,I186_2,I1_2,I146,I147,I148,I166,I269_1,I265,I269_2,I203_1,I262,I203_2,I284_1,
    I284_2,I1_3,I244,I245,I246,I264,I301_1,I359,I301_2,I378_1,I378_2,I1_4,I344,I345,I357,I358,
    I360,I410,I411,I412,I413,I414,I423,I422,I438,I439,I440,I441,I442,I451,I450,I466,
    I467,I468,I469,I470,I479,I478,I494,I495,I496,I497,I498,I506,I505,I546,P_2,I547,
    P_3,I550,I551,I570,P_6,I571,P_7,I574,I575,I594,P_10,I595,P_11,I598,I599,I618,
    P_14,I619,P_15,I622,I623,I73_3,I73_4,I7_3,I7_4,I88_3,I88_4,I171_3,I171_4,I105_3,I105_4,I186_3,
    I186_4,I269_3,I269_4,I203_3,I203_4,I284_3,I284_4,I301_3,I301_4,I378_3,I378_4,I387_1,I2_1,I2_2,I2_3,I408_2,
    I407_1,I407_2,I408_3,I407_3,P_5,I403_2,I404_2,I405_2,P_8,I406_2,P_9,I403_3,I404_3,I405_3,P_12,I406_3,
    P_13,I403_4,I404_4,I405_4,P_16,I406_4,I559_1,P_1,I559_2,I583_1,I583_2,P_4,I607_1,I607_2,I631_1,I631_2,
    I534_5,I70_1,I95_1,I64,I168_1,I193_1,I162,I266_1,I291_1,I260,I363_1,I361,I366_1,I384_1,I555_1,I555_2,
    I579_1,I579_2,I603_1,I603_2,I627_1,I627_2,I534_2,I533_1,I533_2,I534_3,I533_3,I534_4,I533_4,I62,I160,I258,
    I355,I420,I448,I476,I503,I554,I578,I602,I626,extra0,extra1,extra2;

  DFF_X2 DFF_0( .CK(CK), .Q(X_4), .D(I12) );
  DFF_X2 DFF_1( .CK(CK), .Q(X_3), .D(I13) );
  DFF_X1 DFF_2( .CK(CK), .Q(X_2), .D(I14) );
  DFF_X1 DFF_3( .CK(CK), .Q(X_1), .D(I15) );
  DFF_X1 DFF_4( .CK(CK), .Q(X_8), .D(I110) );
  DFF_X1 DFF_5( .CK(CK), .Q(X_7), .D(I111) );
  DFF_X1 DFF_6( .CK(CK), .Q(X_6), .D(I112) );
  DFF_X1 DFF_7( .CK(CK), .Q(X_5), .D(I113) );
  DFF_X1 DFF_8( .CK(CK), .Q(X_12), .D(I208) );
  DFF_X1 DFF_9( .CK(CK), .Q(X_11), .D(I209) );
  DFF_X1 DFF_10( .CK(CK), .Q(X_10), .D(I210) );
  DFF_X1 DFF_11( .CK(CK), .Q(X_9), .D(I211) );
  DFF_X2 DFF_12( .CK(CK), .Q(X_16), .D(I306) );
  DFF_X1 DFF_13( .CK(CK), .Q(X_15), .D(I307) );
  DFF_X1 DFF_14( .CK(CK), .Q(X_14), .D(I308) );
  DFF_X1 DFF_15( .CK(CK), .Q(X_13), .D(I309) );
  INV_X1 NOT_0( .ZN(I73_1), .A(I69) );
  INV_X1 NOT_1( .ZN(I73_2), .A(X_3) );
  INV_X1 NOT_2( .ZN(I7_1), .A(I66) );
  INV_X1 NOT_3( .ZN(I7_2), .A(X_2) );
  INV_X1 NOT_4( .ZN(I88_1), .A(X_1) );
  INV_X1 NOT_5( .ZN(I88_2), .A(P_0) );
  INV_X1 NOT_6( .ZN(I48), .A(P_0) );
  INV_X1 NOT_7( .ZN(I49), .A(X_4) );
  INV_X1 NOT_8( .ZN(I50), .A(X_3) );
  INV_X1 NOT_9( .ZN(I68), .A(I69) );
  INV_X1 NOT_10( .ZN(I171_1), .A(I167) );
  INV_X1 NOT_11( .ZN(I171_2), .A(X_7) );
  INV_X1 NOT_12( .ZN(I105_1), .A(I164) );
  INV_X1 NOT_13( .ZN(I105_2), .A(X_6) );
  INV_X1 NOT_14( .ZN(I186_1), .A(X_5) );
  INV_X1 NOT_15( .ZN(I186_2), .A(I1_2) );
  INV_X1 NOT_16( .ZN(I146), .A(I1_2) );
  INV_X1 NOT_17( .ZN(I147), .A(X_8) );
  INV_X2 NOT_18( .ZN(I148), .A(X_7) );
  INV_X2 NOT_19( .ZN(I166), .A(I167) );
  INV_X2 NOT_20( .ZN(I269_1), .A(I265) );
  INV_X1 NOT_21( .ZN(I269_2), .A(X_11) );
  INV_X1 NOT_22( .ZN(I203_1), .A(I262) );
  INV_X1 NOT_23( .ZN(I203_2), .A(X_10) );
  INV_X1 NOT_24( .ZN(I284_1), .A(X_9) );
  INV_X1 NOT_25( .ZN(I284_2), .A(I1_3) );
  INV_X1 NOT_26( .ZN(I244), .A(I1_3) );
  INV_X1 NOT_27( .ZN(I245), .A(X_12) );
  INV_X1 NOT_28( .ZN(I246), .A(X_11) );
  INV_X1 NOT_29( .ZN(I264), .A(I265) );
  INV_X1 NOT_30( .ZN(I301_1), .A(I359) );
  INV_X1 NOT_31( .ZN(I301_2), .A(X_14) );
  INV_X1 NOT_32( .ZN(I378_1), .A(X_13) );
  INV_X1 NOT_33( .ZN(I378_2), .A(I1_4) );
  INV_X1 NOT_34( .ZN(I344), .A(X_15) );
  INV_X1 NOT_35( .ZN(I345), .A(X_14) );
  INV_X1 NOT_36( .ZN(I357), .A(I358) );
  INV_X1 NOT_37( .ZN(I360), .A(I359) );
  INV_X1 NOT_38( .ZN(I410), .A(P_0) );
  INV_X1 NOT_39( .ZN(I411), .A(X_1) );
  INV_X1 NOT_40( .ZN(I412), .A(X_2) );
  INV_X1 NOT_41( .ZN(I413), .A(X_3) );
  INV_X1 NOT_42( .ZN(I414), .A(X_4) );
  INV_X1 NOT_43( .ZN(I423), .A(I422) );
  INV_X1 NOT_44( .ZN(I438), .A(P_0) );
  INV_X1 NOT_45( .ZN(I439), .A(X_5) );
  INV_X1 NOT_46( .ZN(I440), .A(X_6) );
  INV_X1 NOT_47( .ZN(I441), .A(X_7) );
  INV_X1 NOT_48( .ZN(I442), .A(X_8) );
  INV_X2 NOT_49( .ZN(I451), .A(I450) );
  INV_X2 NOT_50( .ZN(I466), .A(P_0) );
  INV_X2 NOT_51( .ZN(I467), .A(X_9) );
  INV_X1 NOT_52( .ZN(I468), .A(X_10) );
  INV_X1 NOT_53( .ZN(I469), .A(X_11) );
  INV_X1 NOT_54( .ZN(I470), .A(X_12) );
  INV_X1 NOT_55( .ZN(I479), .A(I478) );
  INV_X1 NOT_56( .ZN(I494), .A(P_0) );
  INV_X1 NOT_57( .ZN(I495), .A(X_13) );
  INV_X1 NOT_58( .ZN(I496), .A(X_14) );
  INV_X1 NOT_59( .ZN(I497), .A(X_15) );
  INV_X1 NOT_60( .ZN(I498), .A(X_16) );
  INV_X1 NOT_61( .ZN(I506), .A(I505) );
  INV_X1 NOT_62( .ZN(I546), .A(P_2) );
  INV_X1 NOT_63( .ZN(I547), .A(P_3) );
  INV_X1 NOT_64( .ZN(I550), .A(C_2) );
  INV_X1 NOT_65( .ZN(I551), .A(C_3) );
  INV_X1 NOT_66( .ZN(I570), .A(P_6) );
  INV_X1 NOT_67( .ZN(I571), .A(P_7) );
  INV_X1 NOT_68( .ZN(I574), .A(C_6) );
  INV_X1 NOT_69( .ZN(I575), .A(C_7) );
  INV_X1 NOT_70( .ZN(I594), .A(P_10) );
  INV_X1 NOT_71( .ZN(I595), .A(P_11) );
  INV_X1 NOT_72( .ZN(I598), .A(C_10) );
  INV_X1 NOT_73( .ZN(I599), .A(C_11) );
  INV_X4 NOT_74( .ZN(I618), .A(P_14) );
  INV_X4 NOT_75( .ZN(I619), .A(P_15) );
  INV_X1 NOT_76( .ZN(I622), .A(C_14) );
  INV_X8 NOT_77( .ZN(I623), .A(C_15) );
  AND2_X1 AND2_0( .ZN(I73_3), .A1(I69), .A2(I73_2) );
  AND2_X1 AND2_1( .ZN(I73_4), .A1(X_3), .A2(I73_1) );
  AND2_X1 AND2_2( .ZN(I7_3), .A1(I66), .A2(I7_2) );
  AND2_X1 AND2_3( .ZN(I7_4), .A1(X_2), .A2(I7_1) );
  AND2_X1 AND2_4( .ZN(I88_3), .A1(X_1), .A2(I88_2) );
  AND2_X1 AND2_5( .ZN(I88_4), .A1(P_0), .A2(I88_1) );
  AND2_X1 AND2_6( .ZN(I171_3), .A1(I167), .A2(I171_2) );
  AND2_X1 AND2_7( .ZN(I171_4), .A1(X_7), .A2(I171_1) );
  AND2_X1 AND2_8( .ZN(I105_3), .A1(I164), .A2(I105_2) );
  AND2_X1 AND2_9( .ZN(I105_4), .A1(X_6), .A2(I105_1) );
  AND2_X1 AND2_10( .ZN(I186_3), .A1(X_5), .A2(I186_2) );
  AND2_X2 AND2_11( .ZN(I186_4), .A1(I1_2), .A2(I186_1) );
  AND2_X2 AND2_12( .ZN(I269_3), .A1(I265), .A2(I269_2) );
  AND2_X2 AND2_13( .ZN(I269_4), .A1(X_11), .A2(I269_1) );
  AND2_X1 AND2_14( .ZN(I203_3), .A1(I262), .A2(I203_2) );
  AND2_X1 AND2_15( .ZN(I203_4), .A1(X_10), .A2(I203_1) );
  AND2_X1 AND2_16( .ZN(I284_3), .A1(X_9), .A2(I284_2) );
  AND2_X1 AND2_17( .ZN(I284_4), .A1(I1_3), .A2(I284_1) );
  AND2_X1 AND2_18( .ZN(I301_3), .A1(I359), .A2(I301_2) );
  AND2_X1 AND2_19( .ZN(I301_4), .A1(X_14), .A2(I301_1) );
  AND2_X1 AND2_20( .ZN(I378_3), .A1(X_13), .A2(I378_2) );
  AND2_X1 AND2_21( .ZN(I378_4), .A1(I1_4), .A2(I378_1) );
  AND2_X1 AND2_22( .ZN(I387_1), .A1(I360), .A2(X_14) );
  AND2_X1 AND2_23( .ZN(I1_2), .A1(I2_1), .A2(P_0) );
  AND2_X1 AND2_24( .ZN(I1_3), .A1(I2_2), .A2(I1_2) );
  AND2_X1 AND2_25( .ZN(I1_4), .A1(I2_3), .A2(I1_3) );
  AND2_X1 AND2_26( .ZN(I408_2), .A1(I407_1), .A2(I407_2) );
  AND2_X1 AND2_27( .ZN(I408_3), .A1(I408_2), .A2(I407_3) );
  AND2_X1 AND2_28( .ZN(P_5), .A1(I407_1), .A2(I403_2) );
  AND2_X1 AND2_29( .ZN(P_6), .A1(I407_1), .A2(I404_2) );
  AND2_X1 AND2_30( .ZN(P_7), .A1(I407_1), .A2(I405_2) );
  AND2_X1 AND2_31( .ZN(P_8), .A1(I407_1), .A2(I406_2) );
  AND2_X1 AND2_32( .ZN(P_9), .A1(I408_2), .A2(I403_3) );
  AND2_X1 AND2_33( .ZN(P_10), .A1(I408_2), .A2(I404_3) );
  AND2_X1 AND2_34( .ZN(P_11), .A1(I408_2), .A2(I405_3) );
  AND2_X1 AND2_35( .ZN(P_12), .A1(I408_2), .A2(I406_3) );
  AND2_X1 AND2_36( .ZN(P_13), .A1(I408_3), .A2(I403_4) );
  AND2_X2 AND2_37( .ZN(P_14), .A1(I408_3), .A2(I404_4) );
  AND2_X2 AND2_38( .ZN(P_15), .A1(I408_3), .A2(I405_4) );
  AND2_X2 AND2_39( .ZN(P_16), .A1(I408_3), .A2(I406_4) );
  AND2_X1 AND2_40( .ZN(I559_1), .A1(P_1), .A2(C_1) );
  AND2_X1 AND2_41( .ZN(I559_2), .A1(P_0), .A2(C_0) );
  AND2_X1 AND2_42( .ZN(I583_1), .A1(P_5), .A2(C_5) );
  AND2_X1 AND2_43( .ZN(I583_2), .A1(P_4), .A2(C_4) );
  AND2_X1 AND2_44( .ZN(I607_1), .A1(P_9), .A2(C_9) );
  AND2_X1 AND2_45( .ZN(I607_2), .A1(P_8), .A2(C_8) );
  AND2_X1 AND2_46( .ZN(I631_1), .A1(P_13), .A2(C_13) );
  AND2_X1 AND2_47( .ZN(I631_2), .A1(P_12), .A2(C_12) );
  AND2_X2 AND2_48( .ZN(I534_5), .A1(P_16), .A2(C_16) );
  OR3_X2 OR3_0( .ZN(I70_1), .A1(I68), .A2(X_4), .A3(I50) );
  OR2_X2 OR2_0( .ZN(I13), .A1(I73_3), .A2(I73_4) );
  OR2_X2 OR2_1( .ZN(I15), .A1(I88_3), .A2(I88_4) );
  OR3_X2 OR3_1( .ZN(I95_1), .A1(I64), .A2(I50), .A3(I48) );
  OR3_X1 OR3_2( .ZN(I168_1), .A1(I166), .A2(X_8), .A3(I148) );
  OR2_X1 OR2_2( .ZN(I111), .A1(I171_3), .A2(I171_4) );
  OR2_X1 OR2_3( .ZN(I113), .A1(I186_3), .A2(I186_4) );
  OR3_X1 OR3_3( .ZN(I193_1), .A1(I162), .A2(I148), .A3(I146) );
  OR3_X1 OR3_4( .ZN(I266_1), .A1(I264), .A2(X_12), .A3(I246) );
  OR2_X1 OR2_4( .ZN(I209), .A1(I269_3), .A2(I269_4) );
  OR2_X1 OR2_5( .ZN(I211), .A1(I284_3), .A2(I284_4) );
  OR3_X1 OR3_5( .ZN(I291_1), .A1(I260), .A2(I246), .A3(I244) );
  OR3_X1 OR3_6( .ZN(I363_1), .A1(I361), .A2(X_16), .A3(I344) );
  OR2_X1 OR2_6( .ZN(I366_1), .A1(I361), .A2(X_15) );
  OR2_X1 OR2_7( .ZN(I309), .A1(I378_3), .A2(I378_4) );
  OR3_X1 OR3_7( .ZN(I384_1), .A1(I359), .A2(I345), .A3(I344) );
  OR2_X1 OR2_8( .ZN(I555_1), .A1(I547), .A2(I551) );
  OR2_X1 OR2_9( .ZN(I555_2), .A1(I546), .A2(I550) );
  OR2_X1 OR2_10( .ZN(I579_1), .A1(I571), .A2(I575) );
  OR2_X1 OR2_11( .ZN(I579_2), .A1(I570), .A2(I574) );
  OR2_X1 OR2_12( .ZN(I603_1), .A1(I595), .A2(I599) );
  OR2_X1 OR2_13( .ZN(I603_2), .A1(I594), .A2(I598) );
  OR2_X1 OR2_14( .ZN(I627_1), .A1(I619), .A2(I623) );
  OR2_X1 OR2_15( .ZN(I627_2), .A1(I618), .A2(I622) );
  OR2_X1 OR2_16( .ZN(I534_2), .A1(I533_1), .A2(I533_2) );
  OR2_X1 OR2_17( .ZN(I534_3), .A1(I534_2), .A2(I533_3) );
  OR2_X4 OR2_18( .ZN(I534_4), .A1(I534_3), .A2(I533_4) );
  OR2_X4 OR2_19( .ZN(Z), .A1(I534_4), .A2(I534_5) );
  NAND2_X1 NAND2_0( .ZN(I12), .A1(I70_1), .A2(I62) );
  NAND2_X1 NAND2_1( .ZN(I62), .A1(I95_1), .A2(X_4) );
  NAND2_X1 NAND2_2( .ZN(I64), .A1(X_1), .A2(X_2) );
  NAND2_X1 NAND2_3( .ZN(I66), .A1(X_1), .A2(P_0) );
  NAND2_X1 NAND2_4( .ZN(I110), .A1(I168_1), .A2(I160) );
  NAND2_X1 NAND2_5( .ZN(I160), .A1(I193_1), .A2(X_8) );
  NAND2_X1 NAND2_6( .ZN(I162), .A1(X_5), .A2(X_6) );
  NAND2_X1 NAND2_7( .ZN(I164), .A1(X_5), .A2(I1_2) );
  NAND2_X2 NAND2_8( .ZN(I208), .A1(I266_1), .A2(I258) );
  NAND2_X1 NAND2_9( .ZN(I258), .A1(I291_1), .A2(X_12) );
  NAND2_X1 NAND2_10( .ZN(I260), .A1(X_9), .A2(X_10) );
  NAND2_X1 NAND2_11( .ZN(I262), .A1(X_9), .A2(I1_3) );
  NAND2_X1 NAND2_12( .ZN(I306), .A1(I363_1), .A2(I355) );
  NAND2_X1 NAND2_13( .ZN(I307), .A1(I366_1), .A2(I357) );
  NAND2_X1 NAND2_14( .ZN(I355), .A1(I384_1), .A2(X_16) );
  NAND2_X1 NAND2_15( .ZN(I359), .A1(X_13), .A2(I1_4) );
  NAND2_X1 NAND2_16( .ZN(I361), .A1(I360), .A2(X_14) );
  NAND2_X1 NAND2_17( .ZN(I420), .A1(I423), .A2(I412) );
  NAND2_X1 NAND2_18( .ZN(I422), .A1(I411), .A2(P_0) );
  NAND2_X1 NAND2_19( .ZN(I448), .A1(I451), .A2(I440) );
  NAND2_X1 NAND2_20( .ZN(I450), .A1(I439), .A2(P_0) );
  NAND2_X2 NAND2_21( .ZN(I476), .A1(I479), .A2(I468) );
  NAND2_X2 NAND2_22( .ZN(I478), .A1(I467), .A2(P_0) );
  NAND2_X2 NAND2_23( .ZN(I503), .A1(I506), .A2(I496) );
  NAND2_X1 NAND2_24( .ZN(I505), .A1(I495), .A2(P_0) );
  NAND3_X1 NAND3_0( .ZN(I533_1), .A1(I555_1), .A2(I555_2), .A3(I554) );
  NAND3_X1 NAND3_1( .ZN(I533_2), .A1(I579_1), .A2(I579_2), .A3(I578) );
  NAND3_X1 NAND3_2( .ZN(I533_3), .A1(I603_1), .A2(I603_2), .A3(I602) );
  NAND3_X1 NAND3_3( .ZN(I533_4), .A1(I627_1), .A2(I627_2), .A3(I626) );
  NOR2_X1 NOR2_0( .ZN(I14), .A1(I7_3), .A2(I7_4) );
  NOR3_X1 NOR3_0( .ZN(I2_1), .A1(I64), .A2(I49), .A3(I50) );
  NOR2_X1 NOR2_1( .ZN(I69), .A1(I64), .A2(I48) );
  NOR2_X1 NOR2_2( .ZN(I112), .A1(I105_3), .A2(I105_4) );
  NOR3_X1 NOR3_1( .ZN(I2_2), .A1(I162), .A2(I147), .A3(I148) );
  NOR2_X1 NOR2_3( .ZN(I167), .A1(I162), .A2(I146) );
  NOR2_X1 NOR2_4( .ZN(I210), .A1(I203_3), .A2(I203_4) );
  NOR3_X1 NOR3_2( .ZN(I2_3), .A1(I260), .A2(I245), .A3(I246) );
  NOR2_X1 NOR2_5( .ZN(I265), .A1(I260), .A2(I244) );
  NOR2_X1 NOR2_6( .ZN(I308), .A1(I301_3), .A2(I301_4) );
  NOR2_X1 NOR2_7( .ZN(I358), .A1(I344), .A2(I387_1) );
  NOR2_X1 NOR2_8( .ZN(P_1), .A1(I410), .A2(I411) );
  NOR2_X1 NOR2_9( .ZN(P_2), .A1(I412), .A2(I422) );
  NOR2_X2 NOR2_10( .ZN(P_3), .A1(I413), .A2(I420) );
  NOR3_X2 NOR3_3( .ZN(P_4), .A1(X_3), .A2(I420), .A3(I414) );
  NOR3_X2 NOR4_0_A( .ZN(extra0), .A1(X_4), .A2(X_2), .A3(X_3) );
  NOR2_X1 NOR4_0( .ZN(I407_1), .A1(extra0), .A2(X_1) );
  NOR2_X1 NOR2_11( .ZN(I403_2), .A1(I438), .A2(I439) );
  NOR2_X1 NOR2_12( .ZN(I404_2), .A1(I440), .A2(I450) );
  NOR2_X1 NOR2_13( .ZN(I405_2), .A1(I441), .A2(I448) );
  NOR3_X1 NOR3_4( .ZN(I406_2), .A1(X_7), .A2(I448), .A3(I442) );
  NOR3_X1 NOR4_1_A( .ZN(extra1), .A1(X_8), .A2(X_6), .A3(X_7) );
  NOR2_X1 NOR4_1( .ZN(I407_2), .A1(extra1), .A2(X_5) );
  NOR2_X1 NOR2_14( .ZN(I403_3), .A1(I466), .A2(I467) );
  NOR2_X4 NOR2_15( .ZN(I404_3), .A1(I468), .A2(I478) );
  NOR2_X2 NOR2_16( .ZN(I405_3), .A1(I469), .A2(I476) );
  NOR3_X1 NOR3_5( .ZN(I406_3), .A1(X_11), .A2(I476), .A3(I470) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(X_12), .A2(X_10), .A3(X_11) );
  NOR2_X1 NOR4_2( .ZN(I407_3), .A1(extra2), .A2(X_9) );
  NOR2_X1 NOR2_17( .ZN(I403_4), .A1(I494), .A2(I495) );
  NOR2_X1 NOR2_18( .ZN(I404_4), .A1(I496), .A2(I505) );
  NOR2_X1 NOR2_19( .ZN(I405_4), .A1(I497), .A2(I503) );
  NOR3_X1 NOR3_6( .ZN(I406_4), .A1(X_15), .A2(I503), .A3(I498) );
  NOR2_X1 NOR2_20( .ZN(I554), .A1(I559_1), .A2(I559_2) );
  NOR2_X1 NOR2_21( .ZN(I578), .A1(I583_1), .A2(I583_2) );
  NOR2_X2 NOR2_22( .ZN(I602), .A1(I607_1), .A2(I607_2) );
  NOR2_X1 NOR2_23( .ZN(I626), .A1(I631_1), .A2(I631_2) );

endmodule
