// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module c880(N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,
  N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,
  N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,
  N255,N259,N260,N261,N267,N268,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,
  N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
  N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
  N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
  N865,N866,N874,N878,N879,N880;

  wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,N290,N291,N292,N293,N294,N295,
    N296,N297,N298,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,N317,N318,
    N319,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
    N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
    N353,N354,N355,N356,N357,N360,N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
    N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
    N415,N416,N417,N424,N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,N460,N463,
    N466,N475,N476,N477,N478,N479,N480,N481,N482,N483,N488,N489,N490,N491,N492,N495,
    N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,
    N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
    N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,N544,N547,N550,N551,N552,N553,
    N557,N561,N565,N569,N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,N596,N597,
    N600,N605,N606,N609,N615,N616,N619,N624,N625,N628,N631,N632,N635,N640,N641,N644,
    N650,N651,N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,N678,N682,N686,N687,
    N692,N696,N697,N700,N704,N705,N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
    N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,
    N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
    N766,N769,N770,N771,N772,N773,N777,N778,N781,N782,N785,N786,N787,N788,N789,N790,
    N791,N792,N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,
    N812,N813,N814,N815,N819,N822,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
    N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N851,
    N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,N870,N871,
    N872,N873,N875,N876,N877;

  NAND4_X2 NAND4_1( .ZN(N269), .A1(N1), .A2(N8), .A3(N13), .A4(N17) );
  NAND4_X2 NAND4_2( .ZN(N270), .A1(N1), .A2(N26), .A3(N13), .A4(N17) );
  AND3_X1 AND3_3( .ZN(N273), .A1(N29), .A2(N36), .A3(N42) );
  AND3_X1 AND3_4( .ZN(N276), .A1(N1), .A2(N26), .A3(N51) );
  NAND4_X1 NAND4_5( .ZN(N279), .A1(N1), .A2(N8), .A3(N51), .A4(N17) );
  NAND4_X1 NAND4_6( .ZN(N280), .A1(N1), .A2(N8), .A3(N13), .A4(N55) );
  NAND4_X1 NAND4_7( .ZN(N284), .A1(N59), .A2(N42), .A3(N68), .A4(N72) );
  NAND2_X1 NAND2_8( .ZN(N285), .A1(N29), .A2(N68) );
  NAND3_X1 NAND3_9( .ZN(N286), .A1(N59), .A2(N68), .A3(N74) );
  AND3_X1 AND3_10( .ZN(N287), .A1(N29), .A2(N75), .A3(N80) );
  AND3_X1 AND3_11( .ZN(N290), .A1(N29), .A2(N75), .A3(N42) );
  AND3_X1 AND3_12( .ZN(N291), .A1(N29), .A2(N36), .A3(N80) );
  AND3_X1 AND3_13( .ZN(N292), .A1(N29), .A2(N36), .A3(N42) );
  AND3_X1 AND3_14( .ZN(N293), .A1(N59), .A2(N75), .A3(N80) );
  AND3_X1 AND3_15( .ZN(N294), .A1(N59), .A2(N75), .A3(N42) );
  AND3_X1 AND3_16( .ZN(N295), .A1(N59), .A2(N36), .A3(N80) );
  AND3_X1 AND3_17( .ZN(N296), .A1(N59), .A2(N36), .A3(N42) );
  AND2_X1 AND2_18( .ZN(N297), .A1(N85), .A2(N86) );
  OR2_X1 OR2_19( .ZN(N298), .A1(N87), .A2(N88) );
  NAND2_X1 NAND2_20( .ZN(N301), .A1(N91), .A2(N96) );
  OR2_X1 OR2_21( .ZN(N302), .A1(N91), .A2(N96) );
  NAND2_X1 NAND2_22( .ZN(N303), .A1(N101), .A2(N106) );
  OR2_X1 OR2_23( .ZN(N304), .A1(N101), .A2(N106) );
  NAND2_X1 NAND2_24( .ZN(N305), .A1(N111), .A2(N116) );
  OR2_X1 OR2_25( .ZN(N306), .A1(N111), .A2(N116) );
  NAND2_X1 NAND2_26( .ZN(N307), .A1(N121), .A2(N126) );
  OR2_X1 OR2_27( .ZN(N308), .A1(N121), .A2(N126) );
  AND2_X1 AND2_28( .ZN(N309), .A1(N8), .A2(N138) );
  INV_X1 NOT1_29( .ZN(N310), .A(N268) );
  AND2_X1 AND2_30( .ZN(N316), .A1(N51), .A2(N138) );
  AND2_X1 AND2_31( .ZN(N317), .A1(N17), .A2(N138) );
  AND2_X1 AND2_32( .ZN(N318), .A1(N152), .A2(N138) );
  NAND2_X1 NAND2_33( .ZN(N319), .A1(N59), .A2(N156) );
  NOR2_X1 NOR2_34( .ZN(N322), .A1(N17), .A2(N42) );
  AND2_X1 AND2_35( .ZN(N323), .A1(N17), .A2(N42) );
  NAND2_X1 NAND2_36( .ZN(N324), .A1(N159), .A2(N165) );
  OR2_X1 OR2_37( .ZN(N325), .A1(N159), .A2(N165) );
  NAND2_X1 NAND2_38( .ZN(N326), .A1(N171), .A2(N177) );
  OR2_X1 OR2_39( .ZN(N327), .A1(N171), .A2(N177) );
  NAND2_X1 NAND2_40( .ZN(N328), .A1(N183), .A2(N189) );
  OR2_X1 OR2_41( .ZN(N329), .A1(N183), .A2(N189) );
  NAND2_X1 NAND2_42( .ZN(N330), .A1(N195), .A2(N201) );
  OR2_X1 OR2_43( .ZN(N331), .A1(N195), .A2(N201) );
  AND2_X1 AND2_44( .ZN(N332), .A1(N210), .A2(N91) );
  AND2_X1 AND2_45( .ZN(N333), .A1(N210), .A2(N96) );
  AND2_X1 AND2_46( .ZN(N334), .A1(N210), .A2(N101) );
  AND2_X2 AND2_47( .ZN(N335), .A1(N210), .A2(N106) );
  AND2_X2 AND2_48( .ZN(N336), .A1(N210), .A2(N111) );
  AND2_X4 AND2_49( .ZN(N337), .A1(N255), .A2(N259) );
  AND2_X1 AND2_50( .ZN(N338), .A1(N210), .A2(N116) );
  AND2_X1 AND2_51( .ZN(N339), .A1(N255), .A2(N260) );
  AND2_X1 AND2_52( .ZN(N340), .A1(N210), .A2(N121) );
  AND2_X1 AND2_53( .ZN(N341), .A1(N255), .A2(N267) );
  INV_X1 NOT1_54( .ZN(N342), .A(N269) );
  INV_X1 NOT1_55( .ZN(N343), .A(N273) );
  OR2_X1 OR2_56( .ZN(N344), .A1(N270), .A2(N273) );
  INV_X1 NOT1_57( .ZN(N345), .A(N276) );
  INV_X1 NOT1_58( .ZN(N346), .A(N276) );
  INV_X1 NOT1_59( .ZN(N347), .A(N279) );
  NOR2_X1 NOR2_60( .ZN(N348), .A1(N280), .A2(N284) );
  OR2_X1 OR2_61( .ZN(N349), .A1(N280), .A2(N285) );
  OR2_X1 OR2_62( .ZN(N350), .A1(N280), .A2(N286) );
  INV_X1 NOT1_63( .ZN(N351), .A(N293) );
  INV_X1 NOT1_64( .ZN(N352), .A(N294) );
  INV_X8 NOT1_65( .ZN(N353), .A(N295) );
  INV_X8 NOT1_66( .ZN(N354), .A(N296) );
  NAND2_X1 NAND2_67( .ZN(N355), .A1(N89), .A2(N298) );
  AND2_X1 AND2_68( .ZN(N356), .A1(N90), .A2(N298) );
  NAND2_X1 NAND2_69( .ZN(N357), .A1(N301), .A2(N302) );
  NAND2_X1 NAND2_70( .ZN(N360), .A1(N303), .A2(N304) );
  NAND2_X1 NAND2_71( .ZN(N363), .A1(N305), .A2(N306) );
  NAND2_X1 NAND2_72( .ZN(N366), .A1(N307), .A2(N308) );
  INV_X1 NOT1_73( .ZN(N369), .A(N310) );
  NOR2_X1 NOR2_74( .ZN(N375), .A1(N322), .A2(N323) );
  NAND2_X1 NAND2_75( .ZN(N376), .A1(N324), .A2(N325) );
  NAND2_X1 NAND2_76( .ZN(N379), .A1(N326), .A2(N327) );
  NAND2_X1 NAND2_77( .ZN(N382), .A1(N328), .A2(N329) );
  NAND2_X1 NAND2_78( .ZN(N385), .A1(N330), .A2(N331) );
  BUF_X1 BUFF1_79( .Z(N388), .A(N290) );
  BUF_X1 BUFF1_80( .Z(N389), .A(N291) );
  BUF_X1 BUFF1_81( .Z(N390), .A(N292) );
  BUF_X1 BUFF1_82( .Z(N391), .A(N297) );
  OR2_X1 OR2_83( .ZN(N392), .A1(N270), .A2(N343) );
  INV_X1 NOT1_84( .ZN(N393), .A(N345) );
  INV_X1 NOT1_85( .ZN(N399), .A(N346) );
  AND2_X1 AND2_86( .ZN(N400), .A1(N348), .A2(N73) );
  INV_X1 NOT1_87( .ZN(N401), .A(N349) );
  INV_X1 NOT1_88( .ZN(N402), .A(N350) );
  INV_X2 NOT1_89( .ZN(N403), .A(N355) );
  INV_X1 NOT1_90( .ZN(N404), .A(N357) );
  INV_X1 NOT1_91( .ZN(N405), .A(N360) );
  AND2_X1 AND2_92( .ZN(N406), .A1(N357), .A2(N360) );
  INV_X1 NOT1_93( .ZN(N407), .A(N363) );
  INV_X1 NOT1_94( .ZN(N408), .A(N366) );
  AND2_X1 AND2_95( .ZN(N409), .A1(N363), .A2(N366) );
  NAND2_X1 NAND2_96( .ZN(N410), .A1(N347), .A2(N352) );
  INV_X1 NOT1_97( .ZN(N411), .A(N376) );
  INV_X1 NOT1_98( .ZN(N412), .A(N379) );
  AND2_X1 AND2_99( .ZN(N413), .A1(N376), .A2(N379) );
  INV_X1 NOT1_100( .ZN(N414), .A(N382) );
  INV_X1 NOT1_101( .ZN(N415), .A(N385) );
  AND2_X1 AND2_102( .ZN(N416), .A1(N382), .A2(N385) );
  AND2_X1 AND2_103( .ZN(N417), .A1(N210), .A2(N369) );
  BUF_X4 BUFF1_104( .Z(N418), .A(N342) );
  BUF_X4 BUFF1_105( .Z(N419), .A(N344) );
  BUF_X1 BUFF1_106( .Z(N420), .A(N351) );
  BUF_X1 BUFF1_107( .Z(N421), .A(N353) );
  BUF_X1 BUFF1_108( .Z(N422), .A(N354) );
  BUF_X1 BUFF1_109( .Z(N423), .A(N356) );
  INV_X1 NOT1_110( .ZN(N424), .A(N400) );
  AND2_X1 AND2_111( .ZN(N425), .A1(N404), .A2(N405) );
  AND2_X1 AND2_112( .ZN(N426), .A1(N407), .A2(N408) );
  AND3_X1 AND3_113( .ZN(N427), .A1(N319), .A2(N393), .A3(N55) );
  AND3_X1 AND3_114( .ZN(N432), .A1(N393), .A2(N17), .A3(N287) );
  NAND3_X1 NAND3_115( .ZN(N437), .A1(N393), .A2(N287), .A3(N55) );
  NAND4_X1 NAND4_116( .ZN(N442), .A1(N375), .A2(N59), .A3(N156), .A4(N393) );
  NAND3_X1 NAND3_117( .ZN(N443), .A1(N393), .A2(N319), .A3(N17) );
  AND2_X1 AND2_118( .ZN(N444), .A1(N411), .A2(N412) );
  AND2_X1 AND2_119( .ZN(N445), .A1(N414), .A2(N415) );
  BUF_X1 BUFF1_120( .Z(N446), .A(N392) );
  BUF_X1 BUFF1_121( .Z(N447), .A(N399) );
  BUF_X1 BUFF1_122( .Z(N448), .A(N401) );
  BUF_X1 BUFF1_123( .Z(N449), .A(N402) );
  BUF_X1 BUFF1_124( .Z(N450), .A(N403) );
  INV_X1 NOT1_125( .ZN(N451), .A(N424) );
  NOR2_X1 NOR2_126( .ZN(N460), .A1(N406), .A2(N425) );
  NOR2_X1 NOR2_127( .ZN(N463), .A1(N409), .A2(N426) );
  NAND2_X1 NAND2_128( .ZN(N466), .A1(N442), .A2(N410) );
  AND2_X1 AND2_129( .ZN(N475), .A1(N143), .A2(N427) );
  AND2_X1 AND2_130( .ZN(N476), .A1(N310), .A2(N432) );
  AND2_X1 AND2_131( .ZN(N477), .A1(N146), .A2(N427) );
  AND2_X1 AND2_132( .ZN(N478), .A1(N310), .A2(N432) );
  AND2_X1 AND2_133( .ZN(N479), .A1(N149), .A2(N427) );
  AND2_X1 AND2_134( .ZN(N480), .A1(N310), .A2(N432) );
  AND2_X1 AND2_135( .ZN(N481), .A1(N153), .A2(N427) );
  AND2_X1 AND2_136( .ZN(N482), .A1(N310), .A2(N432) );
  NAND2_X1 NAND2_137( .ZN(N483), .A1(N443), .A2(N1) );
  OR2_X1 OR2_138( .ZN(N488), .A1(N369), .A2(N437) );
  OR2_X1 OR2_139( .ZN(N489), .A1(N369), .A2(N437) );
  OR2_X1 OR2_140( .ZN(N490), .A1(N369), .A2(N437) );
  OR2_X1 OR2_141( .ZN(N491), .A1(N369), .A2(N437) );
  NOR2_X1 NOR2_142( .ZN(N492), .A1(N413), .A2(N444) );
  NOR2_X1 NOR2_143( .ZN(N495), .A1(N416), .A2(N445) );
  NAND2_X1 NAND2_144( .ZN(N498), .A1(N130), .A2(N460) );
  OR2_X1 OR2_145( .ZN(N499), .A1(N130), .A2(N460) );
  NAND2_X1 NAND2_146( .ZN(N500), .A1(N463), .A2(N135) );
  OR2_X1 OR2_147( .ZN(N501), .A1(N463), .A2(N135) );
  AND2_X1 AND2_148( .ZN(N502), .A1(N91), .A2(N466) );
  NOR2_X1 NOR2_149( .ZN(N503), .A1(N475), .A2(N476) );
  AND2_X1 AND2_150( .ZN(N504), .A1(N96), .A2(N466) );
  NOR2_X1 NOR2_151( .ZN(N505), .A1(N477), .A2(N478) );
  AND2_X2 AND2_152( .ZN(N506), .A1(N101), .A2(N466) );
  NOR2_X2 NOR2_153( .ZN(N507), .A1(N479), .A2(N480) );
  AND2_X2 AND2_154( .ZN(N508), .A1(N106), .A2(N466) );
  NOR2_X2 NOR2_155( .ZN(N509), .A1(N481), .A2(N482) );
  AND2_X1 AND2_156( .ZN(N510), .A1(N143), .A2(N483) );
  AND2_X1 AND2_157( .ZN(N511), .A1(N111), .A2(N466) );
  AND2_X1 AND2_158( .ZN(N512), .A1(N146), .A2(N483) );
  AND2_X1 AND2_159( .ZN(N513), .A1(N116), .A2(N466) );
  AND2_X1 AND2_160( .ZN(N514), .A1(N149), .A2(N483) );
  AND2_X1 AND2_161( .ZN(N515), .A1(N121), .A2(N466) );
  AND2_X1 AND2_162( .ZN(N516), .A1(N153), .A2(N483) );
  AND2_X1 AND2_163( .ZN(N517), .A1(N126), .A2(N466) );
  NAND2_X1 NAND2_164( .ZN(N518), .A1(N130), .A2(N492) );
  OR2_X1 OR2_165( .ZN(N519), .A1(N130), .A2(N492) );
  NAND2_X1 NAND2_166( .ZN(N520), .A1(N495), .A2(N207) );
  OR2_X1 OR2_167( .ZN(N521), .A1(N495), .A2(N207) );
  AND2_X1 AND2_168( .ZN(N522), .A1(N451), .A2(N159) );
  AND2_X1 AND2_169( .ZN(N523), .A1(N451), .A2(N165) );
  AND2_X1 AND2_170( .ZN(N524), .A1(N451), .A2(N171) );
  AND2_X1 AND2_171( .ZN(N525), .A1(N451), .A2(N177) );
  AND2_X1 AND2_172( .ZN(N526), .A1(N451), .A2(N183) );
  NAND2_X1 NAND2_173( .ZN(N527), .A1(N451), .A2(N189) );
  NAND2_X1 NAND2_174( .ZN(N528), .A1(N451), .A2(N195) );
  NAND2_X1 NAND2_175( .ZN(N529), .A1(N451), .A2(N201) );
  NAND2_X1 NAND2_176( .ZN(N530), .A1(N498), .A2(N499) );
  NAND2_X1 NAND2_177( .ZN(N533), .A1(N500), .A2(N501) );
  NOR2_X1 NOR2_178( .ZN(N536), .A1(N309), .A2(N502) );
  NOR2_X1 NOR2_179( .ZN(N537), .A1(N316), .A2(N504) );
  NOR2_X1 NOR2_180( .ZN(N538), .A1(N317), .A2(N506) );
  NOR2_X1 NOR2_181( .ZN(N539), .A1(N318), .A2(N508) );
  NOR2_X1 NOR2_182( .ZN(N540), .A1(N510), .A2(N511) );
  NOR2_X1 NOR2_183( .ZN(N541), .A1(N512), .A2(N513) );
  NOR2_X1 NOR2_184( .ZN(N542), .A1(N514), .A2(N515) );
  NOR2_X1 NOR2_185( .ZN(N543), .A1(N516), .A2(N517) );
  NAND2_X1 NAND2_186( .ZN(N544), .A1(N518), .A2(N519) );
  NAND2_X1 NAND2_187( .ZN(N547), .A1(N520), .A2(N521) );
  INV_X1 NOT1_188( .ZN(N550), .A(N530) );
  INV_X1 NOT1_189( .ZN(N551), .A(N533) );
  AND2_X1 AND2_190( .ZN(N552), .A1(N530), .A2(N533) );
  NAND2_X1 NAND2_191( .ZN(N553), .A1(N536), .A2(N503) );
  NAND2_X1 NAND2_192( .ZN(N557), .A1(N537), .A2(N505) );
  NAND2_X1 NAND2_193( .ZN(N561), .A1(N538), .A2(N507) );
  NAND2_X1 NAND2_194( .ZN(N565), .A1(N539), .A2(N509) );
  NAND2_X1 NAND2_195( .ZN(N569), .A1(N488), .A2(N540) );
  NAND2_X1 NAND2_196( .ZN(N573), .A1(N489), .A2(N541) );
  NAND2_X1 NAND2_197( .ZN(N577), .A1(N490), .A2(N542) );
  NAND2_X1 NAND2_198( .ZN(N581), .A1(N491), .A2(N543) );
  INV_X1 NOT1_199( .ZN(N585), .A(N544) );
  INV_X1 NOT1_200( .ZN(N586), .A(N547) );
  AND2_X1 AND2_201( .ZN(N587), .A1(N544), .A2(N547) );
  AND2_X2 AND2_202( .ZN(N588), .A1(N550), .A2(N551) );
  AND2_X1 AND2_203( .ZN(N589), .A1(N585), .A2(N586) );
  NAND2_X1 NAND2_204( .ZN(N590), .A1(N553), .A2(N159) );
  OR2_X1 OR2_205( .ZN(N593), .A1(N553), .A2(N159) );
  AND2_X1 AND2_206( .ZN(N596), .A1(N246), .A2(N553) );
  NAND2_X1 NAND2_207( .ZN(N597), .A1(N557), .A2(N165) );
  OR2_X1 OR2_208( .ZN(N600), .A1(N557), .A2(N165) );
  AND2_X1 AND2_209( .ZN(N605), .A1(N246), .A2(N557) );
  NAND2_X1 NAND2_210( .ZN(N606), .A1(N561), .A2(N171) );
  OR2_X1 OR2_211( .ZN(N609), .A1(N561), .A2(N171) );
  AND2_X1 AND2_212( .ZN(N615), .A1(N246), .A2(N561) );
  NAND2_X1 NAND2_213( .ZN(N616), .A1(N565), .A2(N177) );
  OR2_X1 OR2_214( .ZN(N619), .A1(N565), .A2(N177) );
  AND2_X1 AND2_215( .ZN(N624), .A1(N246), .A2(N565) );
  NAND2_X1 NAND2_216( .ZN(N625), .A1(N569), .A2(N183) );
  OR2_X1 OR2_217( .ZN(N628), .A1(N569), .A2(N183) );
  AND2_X1 AND2_218( .ZN(N631), .A1(N246), .A2(N569) );
  NAND2_X1 NAND2_219( .ZN(N632), .A1(N573), .A2(N189) );
  OR2_X1 OR2_220( .ZN(N635), .A1(N573), .A2(N189) );
  AND2_X1 AND2_221( .ZN(N640), .A1(N246), .A2(N573) );
  NAND2_X1 NAND2_222( .ZN(N641), .A1(N577), .A2(N195) );
  OR2_X1 OR2_223( .ZN(N644), .A1(N577), .A2(N195) );
  AND2_X1 AND2_224( .ZN(N650), .A1(N246), .A2(N577) );
  NAND2_X1 NAND2_225( .ZN(N651), .A1(N581), .A2(N201) );
  OR2_X1 OR2_226( .ZN(N654), .A1(N581), .A2(N201) );
  AND2_X1 AND2_227( .ZN(N659), .A1(N246), .A2(N581) );
  NOR2_X2 NOR2_228( .ZN(N660), .A1(N552), .A2(N588) );
  NOR2_X1 NOR2_229( .ZN(N661), .A1(N587), .A2(N589) );
  INV_X1 NOT1_230( .ZN(N662), .A(N590) );
  AND2_X1 AND2_231( .ZN(N665), .A1(N593), .A2(N590) );
  NOR2_X1 NOR2_232( .ZN(N669), .A1(N596), .A2(N522) );
  INV_X1 NOT1_233( .ZN(N670), .A(N597) );
  AND2_X1 AND2_234( .ZN(N673), .A1(N600), .A2(N597) );
  NOR2_X1 NOR2_235( .ZN(N677), .A1(N605), .A2(N523) );
  INV_X1 NOT1_236( .ZN(N678), .A(N606) );
  AND2_X1 AND2_237( .ZN(N682), .A1(N609), .A2(N606) );
  NOR2_X1 NOR2_238( .ZN(N686), .A1(N615), .A2(N524) );
  INV_X1 NOT1_239( .ZN(N687), .A(N616) );
  AND2_X1 AND2_240( .ZN(N692), .A1(N619), .A2(N616) );
  NOR2_X1 NOR2_241( .ZN(N696), .A1(N624), .A2(N525) );
  INV_X1 NOT1_242( .ZN(N697), .A(N625) );
  AND2_X1 AND2_243( .ZN(N700), .A1(N628), .A2(N625) );
  NOR2_X1 NOR2_244( .ZN(N704), .A1(N631), .A2(N526) );
  INV_X1 NOT1_245( .ZN(N705), .A(N632) );
  AND2_X1 AND2_246( .ZN(N708), .A1(N635), .A2(N632) );
  NOR2_X1 NOR2_247( .ZN(N712), .A1(N337), .A2(N640) );
  INV_X1 NOT1_248( .ZN(N713), .A(N641) );
  AND2_X1 AND2_249( .ZN(N717), .A1(N644), .A2(N641) );
  NOR2_X1 NOR2_250( .ZN(N721), .A1(N339), .A2(N650) );
  INV_X1 NOT1_251( .ZN(N722), .A(N651) );
  AND2_X1 AND2_252( .ZN(N727), .A1(N654), .A2(N651) );
  NOR2_X1 NOR2_253( .ZN(N731), .A1(N341), .A2(N659) );
  NAND2_X1 NAND2_254( .ZN(N732), .A1(N654), .A2(N261) );
  NAND3_X1 NAND3_255( .ZN(N733), .A1(N644), .A2(N654), .A3(N261) );
  NAND4_X1 NAND4_256( .ZN(N734), .A1(N635), .A2(N644), .A3(N654), .A4(N261) );
  INV_X1 NOT1_257( .ZN(N735), .A(N662) );
  AND2_X1 AND2_258( .ZN(N736), .A1(N228), .A2(N665) );
  AND2_X1 AND2_259( .ZN(N737), .A1(N237), .A2(N662) );
  INV_X1 NOT1_260( .ZN(N738), .A(N670) );
  AND2_X1 AND2_261( .ZN(N739), .A1(N228), .A2(N673) );
  AND2_X1 AND2_262( .ZN(N740), .A1(N237), .A2(N670) );
  INV_X1 NOT1_263( .ZN(N741), .A(N678) );
  AND2_X1 AND2_264( .ZN(N742), .A1(N228), .A2(N682) );
  AND2_X1 AND2_265( .ZN(N743), .A1(N237), .A2(N678) );
  INV_X1 NOT1_266( .ZN(N744), .A(N687) );
  AND2_X1 AND2_267( .ZN(N745), .A1(N228), .A2(N692) );
  AND2_X1 AND2_268( .ZN(N746), .A1(N237), .A2(N687) );
  INV_X1 NOT1_269( .ZN(N747), .A(N697) );
  AND2_X1 AND2_270( .ZN(N748), .A1(N228), .A2(N700) );
  AND2_X1 AND2_271( .ZN(N749), .A1(N237), .A2(N697) );
  INV_X1 NOT1_272( .ZN(N750), .A(N705) );
  AND2_X1 AND2_273( .ZN(N751), .A1(N228), .A2(N708) );
  AND2_X1 AND2_274( .ZN(N752), .A1(N237), .A2(N705) );
  INV_X1 NOT1_275( .ZN(N753), .A(N713) );
  AND2_X1 AND2_276( .ZN(N754), .A1(N228), .A2(N717) );
  AND2_X1 AND2_277( .ZN(N755), .A1(N237), .A2(N713) );
  INV_X1 NOT1_278( .ZN(N756), .A(N722) );
  NOR2_X1 NOR2_279( .ZN(N757), .A1(N727), .A2(N261) );
  AND2_X1 AND2_280( .ZN(N758), .A1(N727), .A2(N261) );
  AND2_X1 AND2_281( .ZN(N759), .A1(N228), .A2(N727) );
  AND2_X1 AND2_282( .ZN(N760), .A1(N237), .A2(N722) );
  NAND2_X1 NAND2_283( .ZN(N761), .A1(N644), .A2(N722) );
  NAND2_X1 NAND2_284( .ZN(N762), .A1(N635), .A2(N713) );
  NAND3_X1 NAND3_285( .ZN(N763), .A1(N635), .A2(N644), .A3(N722) );
  NAND2_X1 NAND2_286( .ZN(N764), .A1(N609), .A2(N687) );
  NAND2_X1 NAND2_287( .ZN(N765), .A1(N600), .A2(N678) );
  NAND3_X1 NAND3_288( .ZN(N766), .A1(N600), .A2(N609), .A3(N687) );
  BUF_X1 BUFF1_289( .Z(N767), .A(N660) );
  BUF_X1 BUFF1_290( .Z(N768), .A(N661) );
  NOR2_X1 NOR2_291( .ZN(N769), .A1(N736), .A2(N737) );
  NOR2_X1 NOR2_292( .ZN(N770), .A1(N739), .A2(N740) );
  NOR2_X1 NOR2_293( .ZN(N771), .A1(N742), .A2(N743) );
  NOR2_X1 NOR2_294( .ZN(N772), .A1(N745), .A2(N746) );
  NAND4_X1 NAND4_295( .ZN(N773), .A1(N750), .A2(N762), .A3(N763), .A4(N734) );
  NOR2_X1 NOR2_296( .ZN(N777), .A1(N748), .A2(N749) );
  NAND3_X1 NAND3_297( .ZN(N778), .A1(N753), .A2(N761), .A3(N733) );
  NOR2_X1 NOR2_298( .ZN(N781), .A1(N751), .A2(N752) );
  NAND2_X1 NAND2_299( .ZN(N782), .A1(N756), .A2(N732) );
  NOR2_X2 NOR2_300( .ZN(N785), .A1(N754), .A2(N755) );
  NOR2_X2 NOR2_301( .ZN(N786), .A1(N757), .A2(N758) );
  NOR2_X2 NOR2_302( .ZN(N787), .A1(N759), .A2(N760) );
  NOR2_X2 NOR2_303( .ZN(N788), .A1(N700), .A2(N773) );
  AND2_X1 AND2_304( .ZN(N789), .A1(N700), .A2(N773) );
  NOR2_X1 NOR2_305( .ZN(N790), .A1(N708), .A2(N778) );
  AND2_X1 AND2_306( .ZN(N791), .A1(N708), .A2(N778) );
  NOR2_X1 NOR2_307( .ZN(N792), .A1(N717), .A2(N782) );
  AND2_X1 AND2_308( .ZN(N793), .A1(N717), .A2(N782) );
  AND2_X1 AND2_309( .ZN(N794), .A1(N219), .A2(N786) );
  NAND2_X1 NAND2_310( .ZN(N795), .A1(N628), .A2(N773) );
  NAND2_X1 NAND2_311( .ZN(N796), .A1(N795), .A2(N747) );
  NOR2_X1 NOR2_312( .ZN(N802), .A1(N788), .A2(N789) );
  NOR2_X1 NOR2_313( .ZN(N803), .A1(N790), .A2(N791) );
  NOR2_X1 NOR2_314( .ZN(N804), .A1(N792), .A2(N793) );
  NOR2_X1 NOR2_315( .ZN(N805), .A1(N340), .A2(N794) );
  NOR2_X1 NOR2_316( .ZN(N806), .A1(N692), .A2(N796) );
  AND2_X1 AND2_317( .ZN(N807), .A1(N692), .A2(N796) );
  AND2_X1 AND2_318( .ZN(N808), .A1(N219), .A2(N802) );
  AND2_X1 AND2_319( .ZN(N809), .A1(N219), .A2(N803) );
  AND2_X1 AND2_320( .ZN(N810), .A1(N219), .A2(N804) );
  NAND4_X1 NAND4_321( .ZN(N811), .A1(N805), .A2(N787), .A3(N731), .A4(N529) );
  NAND2_X1 NAND2_322( .ZN(N812), .A1(N619), .A2(N796) );
  NAND3_X1 NAND3_323( .ZN(N813), .A1(N609), .A2(N619), .A3(N796) );
  NAND4_X1 NAND4_324( .ZN(N814), .A1(N600), .A2(N609), .A3(N619), .A4(N796) );
  NAND4_X1 NAND4_325( .ZN(N815), .A1(N738), .A2(N765), .A3(N766), .A4(N814) );
  NAND3_X1 NAND3_326( .ZN(N819), .A1(N741), .A2(N764), .A3(N813) );
  NAND2_X1 NAND2_327( .ZN(N822), .A1(N744), .A2(N812) );
  NOR2_X1 NOR2_328( .ZN(N825), .A1(N806), .A2(N807) );
  NOR2_X1 NOR2_329( .ZN(N826), .A1(N335), .A2(N808) );
  NOR2_X1 NOR2_330( .ZN(N827), .A1(N336), .A2(N809) );
  NOR2_X1 NOR2_331( .ZN(N828), .A1(N338), .A2(N810) );
  INV_X8 NOT1_332( .ZN(N829), .A(N811) );
  NOR2_X1 NOR2_333( .ZN(N830), .A1(N665), .A2(N815) );
  AND2_X1 AND2_334( .ZN(N831), .A1(N665), .A2(N815) );
  NOR2_X1 NOR2_335( .ZN(N832), .A1(N673), .A2(N819) );
  AND2_X2 AND2_336( .ZN(N833), .A1(N673), .A2(N819) );
  NOR2_X2 NOR2_337( .ZN(N834), .A1(N682), .A2(N822) );
  AND2_X1 AND2_338( .ZN(N835), .A1(N682), .A2(N822) );
  AND2_X1 AND2_339( .ZN(N836), .A1(N219), .A2(N825) );
  NAND3_X1 NAND3_340( .ZN(N837), .A1(N826), .A2(N777), .A3(N704) );
  NAND4_X1 NAND4_341( .ZN(N838), .A1(N827), .A2(N781), .A3(N712), .A4(N527) );
  NAND4_X1 NAND4_342( .ZN(N839), .A1(N828), .A2(N785), .A3(N721), .A4(N528) );
  INV_X1 NOT1_343( .ZN(N840), .A(N829) );
  NAND2_X1 NAND2_344( .ZN(N841), .A1(N815), .A2(N593) );
  NOR2_X1 NOR2_345( .ZN(N842), .A1(N830), .A2(N831) );
  NOR2_X1 NOR2_346( .ZN(N843), .A1(N832), .A2(N833) );
  NOR2_X1 NOR2_347( .ZN(N844), .A1(N834), .A2(N835) );
  NOR2_X1 NOR2_348( .ZN(N845), .A1(N334), .A2(N836) );
  INV_X1 NOT1_349( .ZN(N846), .A(N837) );
  INV_X1 NOT1_350( .ZN(N847), .A(N838) );
  INV_X1 NOT1_351( .ZN(N848), .A(N839) );
  AND2_X1 AND2_352( .ZN(N849), .A1(N735), .A2(N841) );
  BUF_X1 BUFF1_353( .Z(N850), .A(N840) );
  AND2_X1 AND2_354( .ZN(N851), .A1(N219), .A2(N842) );
  AND2_X1 AND2_355( .ZN(N852), .A1(N219), .A2(N843) );
  AND2_X1 AND2_356( .ZN(N853), .A1(N219), .A2(N844) );
  NAND3_X1 NAND3_357( .ZN(N854), .A1(N845), .A2(N772), .A3(N696) );
  INV_X1 NOT1_358( .ZN(N855), .A(N846) );
  INV_X1 NOT1_359( .ZN(N856), .A(N847) );
  INV_X1 NOT1_360( .ZN(N857), .A(N848) );
  INV_X1 NOT1_361( .ZN(N858), .A(N849) );
  NOR2_X1 NOR2_362( .ZN(N859), .A1(N417), .A2(N851) );
  NOR2_X1 NOR2_363( .ZN(N860), .A1(N332), .A2(N852) );
  NOR2_X1 NOR2_364( .ZN(N861), .A1(N333), .A2(N853) );
  INV_X1 NOT1_365( .ZN(N862), .A(N854) );
  BUF_X1 BUFF1_366( .Z(N863), .A(N855) );
  BUF_X1 BUFF1_367( .Z(N864), .A(N856) );
  BUF_X1 BUFF1_368( .Z(N865), .A(N857) );
  BUF_X1 BUFF1_369( .Z(N866), .A(N858) );
  NAND3_X1 NAND3_370( .ZN(N867), .A1(N859), .A2(N769), .A3(N669) );
  NAND3_X1 NAND3_371( .ZN(N868), .A1(N860), .A2(N770), .A3(N677) );
  NAND3_X1 NAND3_372( .ZN(N869), .A1(N861), .A2(N771), .A3(N686) );
  INV_X1 NOT1_373( .ZN(N870), .A(N862) );
  INV_X1 NOT1_374( .ZN(N871), .A(N867) );
  INV_X4 NOT1_375( .ZN(N872), .A(N868) );
  INV_X1 NOT1_376( .ZN(N873), .A(N869) );
  BUF_X1 BUFF1_377( .Z(N874), .A(N870) );
  INV_X1 NOT1_378( .ZN(N875), .A(N871) );
  INV_X1 NOT1_379( .ZN(N876), .A(N872) );
  INV_X1 NOT1_380( .ZN(N877), .A(N873) );
  BUF_X1 BUFF1_381( .Z(N878), .A(N875) );
  BUF_X2 BUFF1_382( .Z(N879), .A(N876) );
  BUF_X1 BUFF1_383( .Z(N880), .A(N877) );

endmodule
