//# 9 inputs
//# 11 outputs
//# 15 D-type flipflops
//# 59 inverters
//# 101 gates (44 ANDs + 18 NANDs + 9 ORs + 30 NORs)

module s344(CK,A0,A1,A2,A3,B0,B1,B2,B3,CNTVCO2,CNTVCON2,P0,P1,P2,P3,P4,
  P5,P6,P7,READY,START);
input CK,START,B0,B1,B2,B3,A0,A1,A2,A3;
output P4,P5,P6,P7,P0,P1,P2,P3,CNTVCON2,CNTVCO2,READY;

  wire CT2,CNTVG3VD,CT1,CNTVG2VD,CT0,CNTVG1VD,ACVQN3,ACVG4VD1,ACVQN2,ACVG3VD1,ACVQN1,ACVG2VD1,ACVQN0,ACVG1VD1,MRVQN3,MRVG4VD,
    MRVQN2,MRVG3VD,MRVQN1,MRVG2VD,MRVQN0,MRVG1VD,AX3,AM3,AX2,AM2,AX1,AM1,AX0,AM0,CNTVG3VQN,CNTVG2VQN,
    CNTVG1VQN,CNTVCON0,CT1N,ACVPCN,CNTVCO0,AMVS0N,IINIIT,READYN,BMVS0N,AMVG5VS0P,AMVG4VS0P,AMVG3VS0P,AMVG2VS0P,AD0,AD0N,AD1,
    AD1N,AD2,AD2N,AD3,AD3N,CNTVG3VD1,CNTVCON1,CNTVG1VD1,BMVG5VS0P,BMVG4VS0P,BMVG3VS0P,BMVG2VS0P,SMVS0N,ADSH,MRVSHLDN,ADDVC1,
    ADDVG1VCN,SMVG5VS0P,SMVG4VS0P,SMVG3VS0P,SMVG2VS0P,CNTVG1VZ,CNTVG1VZ1,AMVG5VX,AMVG4VX,AMVG3VX,AMVG2VX,S0,ADDVG1VP,BM3,BMVG5VX,BM2,
    BMVG4VX,BM1,BMVG3VX,BM0,BMVG2VX,ADDVC2,ADDVG2VCN,S1,ADDVG2VSN,ADDVC3,ADDVG3VCN,S2,ADDVG3VSN,SM0,SMVG2VX,CO,
    ADDVG4VCN,S3,ADDVG4VSN,SM1,SMVG3VX,SM3,SMVG5VX,SM2,SMVG4VX,AMVG5VG1VAD1NF,AMVG4VG1VAD1NF,AMVG3VG1VAD1NF,AMVG2VG1VAD1NF,BMVG5VG1VAD1NF,BMVG4VG1VAD1NF,BMVG3VG1VAD1NF,
    BMVG2VG1VAD1NF,AMVG5VG1VAD2NF,AMVG4VG1VAD2NF,AMVG3VG1VAD2NF,AMVG2VG1VAD2NF,ADDVG2VCNVAD1NF,ADDVG3VCNVAD1NF,ADDVG4VCNVAD1NF,MRVG3VDVAD1NF,MRVG2VDVAD1NF,MRVG1VDVAD1NF,BMVG5VG1VAD2NF,BMVG4VG1VAD2NF,BMVG3VG1VAD2NF,BMVG2VG1VAD2NF,SMVG5VG1VAD1NF,
    SMVG4VG1VAD1NF,SMVG3VG1VAD1NF,SMVG2VG1VAD1NF,ADDVG2VCNVAD4NF,ADDVG2VCNVAD2NF,ADDVG2VCNVOR1NF,MRVG4VDVAD1NF,MRVG4VDVAD2NF,MRVG3VDVAD2NF,MRVG2VDVAD2NF,MRVG1VDVAD2NF,ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG3VCNVAD4NF,ADDVG3VCNVAD2NF,ADDVG3VCNVOR1NF,
    ADDVG3VCNVAD3NF,ADDVG3VCNVOR2NF,SMVG2VG1VAD2NF,ADDVG4VCNVAD4NF,ADDVG4VCNVAD2NF,ADDVG4VCNVOR1NF,ADDVG4VCNVAD3NF,ADDVG4VCNVOR2NF,SMVG3VG1VAD2NF,SMVG5VG1VAD2NF,SMVG4VG1VAD2NF,ADDVG1VPVOR1NF,CNTVG3VG2VOR1NF,CNTVG2VG2VOR1NF,CNTVG2VD1,CNTVCO1,
    CNTVG3VZ1,CNTVG2VZ1,CNTVG3VZ,CNTVG2VZ;

  DFF_X1 DFF_0( .CK(CK), .Q(CT2), .D(CNTVG3VD) );
  DFF_X1 DFF_1( .CK(CK), .Q(CT1), .D(CNTVG2VD) );
  DFF_X1 DFF_2( .CK(CK), .Q(CT0), .D(CNTVG1VD) );
  DFF_X2 DFF_3( .CK(CK), .Q(ACVQN3), .D(ACVG4VD1) );
  DFF_X2 DFF_4( .CK(CK), .Q(ACVQN2), .D(ACVG3VD1) );
  DFF_X2 DFF_5( .CK(CK), .Q(ACVQN1), .D(ACVG2VD1) );
  DFF_X2 DFF_6( .CK(CK), .Q(ACVQN0), .D(ACVG1VD1) );
  DFF_X1 DFF_7( .CK(CK), .Q(MRVQN3), .D(MRVG4VD) );
  DFF_X1 DFF_8( .CK(CK), .Q(MRVQN2), .D(MRVG3VD) );
  DFF_X1 DFF_9( .CK(CK), .Q(MRVQN1), .D(MRVG2VD) );
  DFF_X1 DFF_10( .CK(CK), .Q(MRVQN0), .D(MRVG1VD) );
  DFF_X1 DFF_11( .CK(CK), .Q(AX3), .D(AM3) );
  DFF_X1 DFF_12( .CK(CK), .Q(AX2), .D(AM2) );
  DFF_X1 DFF_13( .CK(CK), .Q(AX1), .D(AM1) );
  DFF_X1 DFF_14( .CK(CK), .Q(AX0), .D(AM0) );
  INV_X1 NOT_0( .ZN(CNTVG3VQN), .A(CT2) );
  INV_X1 NOT_1( .ZN(CNTVG2VQN), .A(CT1) );
  INV_X1 NOT_2( .ZN(CNTVG1VQN), .A(CT0) );
  INV_X1 NOT_3( .ZN(P7), .A(ACVQN3) );
  INV_X1 NOT_4( .ZN(P6), .A(ACVQN2) );
  INV_X1 NOT_5( .ZN(P5), .A(ACVQN1) );
  INV_X1 NOT_6( .ZN(P4), .A(ACVQN0) );
  INV_X1 NOT_7( .ZN(P3), .A(MRVQN3) );
  INV_X1 NOT_8( .ZN(P2), .A(MRVQN2) );
  INV_X1 NOT_9( .ZN(P1), .A(MRVQN1) );
  INV_X1 NOT_10( .ZN(P0), .A(MRVQN0) );
  INV_X1 NOT_11( .ZN(CNTVCON0), .A(CT0) );
  INV_X2 NOT_12( .ZN(CT1N), .A(CT1) );
  INV_X4 NOT_13( .ZN(ACVPCN), .A(START) );
  INV_X2 NOT_14( .ZN(CNTVCO0), .A(CNTVG1VQN) );
  INV_X1 NOT_15( .ZN(AMVS0N), .A(IINIIT) );
  INV_X1 NOT_16( .ZN(READY), .A(READYN) );
  INV_X1 NOT_17( .ZN(BMVS0N), .A(READYN) );
  INV_X1 NOT_18( .ZN(AMVG5VS0P), .A(AMVS0N) );
  INV_X1 NOT_19( .ZN(AMVG4VS0P), .A(AMVS0N) );
  INV_X1 NOT_20( .ZN(AMVG3VS0P), .A(AMVS0N) );
  INV_X1 NOT_21( .ZN(AMVG2VS0P), .A(AMVS0N) );
  INV_X1 NOT_22( .ZN(AD0), .A(AD0N) );
  INV_X1 NOT_23( .ZN(AD1), .A(AD1N) );
  INV_X1 NOT_24( .ZN(AD2), .A(AD2N) );
  INV_X1 NOT_25( .ZN(AD3), .A(AD3N) );
  INV_X1 NOT_26( .ZN(CNTVG3VD1), .A(CNTVCON1) );
  INV_X1 NOT_27( .ZN(CNTVG1VD1), .A(READY) );
  INV_X1 NOT_28( .ZN(BMVG5VS0P), .A(BMVS0N) );
  INV_X1 NOT_29( .ZN(BMVG4VS0P), .A(BMVS0N) );
  INV_X1 NOT_30( .ZN(BMVG3VS0P), .A(BMVS0N) );
  INV_X2 NOT_31( .ZN(BMVG2VS0P), .A(BMVS0N) );
  INV_X2 NOT_32( .ZN(SMVS0N), .A(ADSH) );
  INV_X2 NOT_33( .ZN(MRVSHLDN), .A(ADSH) );
  INV_X8 NOT_34( .ZN(ADDVC1), .A(ADDVG1VCN) );
  INV_X1 NOT_35( .ZN(SMVG5VS0P), .A(SMVS0N) );
  INV_X1 NOT_36( .ZN(SMVG4VS0P), .A(SMVS0N) );
  INV_X1 NOT_37( .ZN(SMVG3VS0P), .A(SMVS0N) );
  INV_X1 NOT_38( .ZN(SMVG2VS0P), .A(SMVS0N) );
  INV_X1 NOT_39( .ZN(CNTVG1VZ), .A(CNTVG1VZ1) );
  INV_X1 NOT_40( .ZN(AM3), .A(AMVG5VX) );
  INV_X1 NOT_41( .ZN(AM2), .A(AMVG4VX) );
  INV_X1 NOT_42( .ZN(AM1), .A(AMVG3VX) );
  INV_X1 NOT_43( .ZN(AM0), .A(AMVG2VX) );
  INV_X1 NOT_44( .ZN(S0), .A(ADDVG1VP) );
  INV_X1 NOT_45( .ZN(BM3), .A(BMVG5VX) );
  INV_X1 NOT_46( .ZN(BM2), .A(BMVG4VX) );
  INV_X1 NOT_47( .ZN(BM1), .A(BMVG3VX) );
  INV_X1 NOT_48( .ZN(BM0), .A(BMVG2VX) );
  INV_X1 NOT_49( .ZN(ADDVC2), .A(ADDVG2VCN) );
  INV_X1 NOT_50( .ZN(S1), .A(ADDVG2VSN) );
  INV_X1 NOT_51( .ZN(ADDVC3), .A(ADDVG3VCN) );
  INV_X1 NOT_52( .ZN(S2), .A(ADDVG3VSN) );
  INV_X1 NOT_53( .ZN(SM0), .A(SMVG2VX) );
  INV_X1 NOT_54( .ZN(CO), .A(ADDVG4VCN) );
  INV_X1 NOT_55( .ZN(S3), .A(ADDVG4VSN) );
  INV_X1 NOT_56( .ZN(SM1), .A(SMVG3VX) );
  INV_X1 NOT_57( .ZN(SM3), .A(SMVG5VX) );
  INV_X1 NOT_58( .ZN(SM2), .A(SMVG4VX) );
  AND2_X1 AND2_0( .ZN(AMVG5VG1VAD1NF), .A1(AMVS0N), .A2(AX3) );
  AND2_X1 AND2_1( .ZN(AMVG4VG1VAD1NF), .A1(AMVS0N), .A2(AX2) );
  AND2_X1 AND2_2( .ZN(AMVG3VG1VAD1NF), .A1(AMVS0N), .A2(AX1) );
  AND2_X1 AND2_3( .ZN(AMVG2VG1VAD1NF), .A1(AMVS0N), .A2(AX0) );
  AND2_X1 AND2_4( .ZN(BMVG5VG1VAD1NF), .A1(BMVS0N), .A2(P3) );
  AND2_X1 AND2_5( .ZN(BMVG4VG1VAD1NF), .A1(BMVS0N), .A2(P2) );
  AND2_X1 AND2_6( .ZN(BMVG3VG1VAD1NF), .A1(BMVS0N), .A2(P1) );
  AND2_X1 AND2_7( .ZN(BMVG2VG1VAD1NF), .A1(BMVS0N), .A2(P0) );
  AND2_X1 AND2_8( .ZN(AMVG5VG1VAD2NF), .A1(AMVG5VS0P), .A2(A3) );
  AND2_X1 AND2_9( .ZN(AMVG4VG1VAD2NF), .A1(AMVG4VS0P), .A2(A2) );
  AND2_X1 AND2_10( .ZN(AMVG3VG1VAD2NF), .A1(AMVG3VS0P), .A2(A1) );
  AND2_X1 AND2_11( .ZN(AMVG2VG1VAD2NF), .A1(AMVG2VS0P), .A2(A0) );
  AND2_X1 AND2_12( .ZN(ADDVG2VCNVAD1NF), .A1(AD1), .A2(P5) );
  AND2_X1 AND2_13( .ZN(ADDVG3VCNVAD1NF), .A1(AD2), .A2(P6) );
  AND2_X1 AND2_14( .ZN(ADDVG4VCNVAD1NF), .A1(AD3), .A2(P7) );
  AND2_X1 AND2_15( .ZN(MRVG3VDVAD1NF), .A1(ADSH), .A2(P3) );
  AND2_X1 AND2_16( .ZN(MRVG2VDVAD1NF), .A1(ADSH), .A2(P2) );
  AND2_X1 AND2_17( .ZN(MRVG1VDVAD1NF), .A1(ADSH), .A2(P1) );
  AND2_X1 AND2_18( .ZN(BMVG5VG1VAD2NF), .A1(BMVG5VS0P), .A2(B3) );
  AND2_X1 AND2_19( .ZN(BMVG4VG1VAD2NF), .A1(BMVG4VS0P), .A2(B2) );
  AND2_X1 AND2_20( .ZN(BMVG3VG1VAD2NF), .A1(BMVG3VS0P), .A2(B1) );
  AND2_X2 AND2_21( .ZN(BMVG2VG1VAD2NF), .A1(BMVG2VS0P), .A2(B0) );
  AND2_X2 AND2_22( .ZN(SMVG5VG1VAD1NF), .A1(SMVS0N), .A2(P7) );
  AND2_X2 AND2_23( .ZN(SMVG4VG1VAD1NF), .A1(SMVS0N), .A2(P6) );
  AND2_X2 AND2_24( .ZN(SMVG3VG1VAD1NF), .A1(SMVS0N), .A2(P5) );
  AND2_X1 AND2_25( .ZN(SMVG2VG1VAD1NF), .A1(SMVS0N), .A2(P4) );
  AND3_X1 AND3_0( .ZN(ADDVG2VCNVAD4NF), .A1(ADDVC1), .A2(AD1), .A3(P5) );
  AND2_X1 AND2_26( .ZN(ADDVG2VCNVAD2NF), .A1(ADDVC1), .A2(ADDVG2VCNVOR1NF) );
  AND2_X1 AND2_27( .ZN(MRVG4VDVAD1NF), .A1(ADSH), .A2(S0) );
  AND2_X1 AND2_28( .ZN(MRVG4VDVAD2NF), .A1(MRVSHLDN), .A2(BM3) );
  AND2_X1 AND2_29( .ZN(MRVG3VDVAD2NF), .A1(MRVSHLDN), .A2(BM2) );
  AND2_X1 AND2_30( .ZN(MRVG2VDVAD2NF), .A1(MRVSHLDN), .A2(BM1) );
  AND2_X1 AND2_31( .ZN(MRVG1VDVAD2NF), .A1(MRVSHLDN), .A2(BM0) );
  AND2_X1 AND2_32( .ZN(ADDVG2VCNVAD3NF), .A1(ADDVG2VCNVOR2NF), .A2(ADDVG2VCN) );
  AND3_X1 AND3_1( .ZN(ADDVG3VCNVAD4NF), .A1(ADDVC2), .A2(AD2), .A3(P6) );
  AND2_X1 AND2_33( .ZN(ADDVG3VCNVAD2NF), .A1(ADDVC2), .A2(ADDVG3VCNVOR1NF) );
  AND2_X1 AND2_34( .ZN(ADDVG3VCNVAD3NF), .A1(ADDVG3VCNVOR2NF), .A2(ADDVG3VCN) );
  AND2_X1 AND2_35( .ZN(SMVG2VG1VAD2NF), .A1(SMVG2VS0P), .A2(S1) );
  AND3_X1 AND3_2( .ZN(ADDVG4VCNVAD4NF), .A1(ADDVC3), .A2(AD3), .A3(P7) );
  AND2_X1 AND2_36( .ZN(ADDVG4VCNVAD2NF), .A1(ADDVC3), .A2(ADDVG4VCNVOR1NF) );
  AND2_X1 AND2_37( .ZN(ADDVG4VCNVAD3NF), .A1(ADDVG4VCNVOR2NF), .A2(ADDVG4VCN) );
  AND2_X1 AND2_38( .ZN(SMVG3VG1VAD2NF), .A1(SMVG3VS0P), .A2(S2) );
  AND2_X1 AND2_39( .ZN(SMVG5VG1VAD2NF), .A1(SMVG5VS0P), .A2(CO) );
  AND2_X1 AND2_40( .ZN(SMVG4VG1VAD2NF), .A1(SMVG4VS0P), .A2(S3) );
  OR2_X1 OR2_0( .ZN(ADDVG1VPVOR1NF), .A1(AD0), .A2(P4) );
  OR2_X1 OR2_1( .ZN(ADDVG2VCNVOR1NF), .A1(AD1), .A2(P5) );
  OR2_X1 OR2_2( .ZN(ADDVG3VCNVOR1NF), .A1(AD2), .A2(P6) );
  OR2_X1 OR2_3( .ZN(ADDVG4VCNVOR1NF), .A1(AD3), .A2(P7) );
  OR2_X1 OR2_4( .ZN(CNTVG3VG2VOR1NF), .A1(CT2), .A2(CNTVG3VD1) );
  OR2_X2 OR2_5( .ZN(CNTVG2VG2VOR1NF), .A1(CT1), .A2(CNTVG2VD1) );
  OR3_X2 OR3_0( .ZN(ADDVG2VCNVOR2NF), .A1(ADDVC1), .A2(AD1), .A3(P5) );
  OR3_X1 OR3_1( .ZN(ADDVG3VCNVOR2NF), .A1(ADDVC2), .A2(AD2), .A3(P6) );
  OR3_X1 OR3_2( .ZN(ADDVG4VCNVOR2NF), .A1(ADDVC3), .A2(AD3), .A3(P7) );
  NAND3_X1 NAND3_0( .ZN(READYN), .A1(CT0), .A2(CT1N), .A3(CT2) );
  NAND2_X1 NAND2_0( .ZN(AD0N), .A1(P0), .A2(AX0) );
  NAND2_X1 NAND2_1( .ZN(AD1N), .A1(P0), .A2(AX1) );
  NAND2_X1 NAND2_2( .ZN(AD2N), .A1(P0), .A2(AX2) );
  NAND2_X1 NAND2_3( .ZN(AD3N), .A1(P0), .A2(AX3) );
  NAND2_X1 NAND2_4( .ZN(CNTVCON1), .A1(CT1), .A2(CNTVCO0) );
  NAND2_X1 NAND2_5( .ZN(CNTVCON2), .A1(CT2), .A2(CNTVCO1) );
  NAND2_X1 NAND2_6( .ZN(ADDVG1VCN), .A1(AD0), .A2(P4) );
  NAND2_X1 NAND2_7( .ZN(CNTVG3VZ1), .A1(CT2), .A2(CNTVG3VD1) );
  NAND2_X1 NAND2_8( .ZN(CNTVG2VZ1), .A1(CT1), .A2(CNTVG2VD1) );
  NAND2_X1 NAND2_9( .ZN(CNTVG1VZ1), .A1(CT0), .A2(CNTVG1VD1) );
  NAND2_X2 NAND2_10( .ZN(ADDVG1VP), .A1(ADDVG1VPVOR1NF), .A2(ADDVG1VCN) );
  NAND2_X2 NAND2_11( .ZN(CNTVG3VZ), .A1(CNTVG3VG2VOR1NF), .A2(CNTVG3VZ1) );
  NAND2_X2 NAND2_12( .ZN(CNTVG2VZ), .A1(CNTVG2VG2VOR1NF), .A2(CNTVG2VZ1) );
  NAND2_X2 NAND2_13( .ZN(ACVG1VD1), .A1(ACVPCN), .A2(SM0) );
  NAND2_X1 NAND2_14( .ZN(ACVG2VD1), .A1(ACVPCN), .A2(SM1) );
  NAND2_X1 NAND2_15( .ZN(ACVG4VD1), .A1(ACVPCN), .A2(SM3) );
  NAND2_X1 NAND2_16( .ZN(ACVG3VD1), .A1(ACVPCN), .A2(SM2) );
  NOR3_X1 NOR3_0( .ZN(IINIIT), .A1(CT0), .A2(CT1), .A3(CT2) );
  NOR2_X1 NOR2_0( .ZN(CNTVCO1), .A1(CNTVG2VQN), .A2(CNTVCON0) );
  NOR2_X1 NOR2_1( .ZN(CNTVCO2), .A1(CNTVG3VQN), .A2(CNTVCON1) );
  NOR2_X1 NOR2_2( .ZN(ADSH), .A1(READY), .A2(IINIIT) );
  NOR2_X1 NOR2_3( .ZN(CNTVG2VD1), .A1(READY), .A2(CNTVCON0) );
  NOR2_X1 NOR2_4( .ZN(AMVG5VX), .A1(AMVG5VG1VAD2NF), .A2(AMVG5VG1VAD1NF) );
  NOR2_X1 NOR2_5( .ZN(AMVG4VX), .A1(AMVG4VG1VAD2NF), .A2(AMVG4VG1VAD1NF) );
  NOR2_X1 NOR2_6( .ZN(AMVG3VX), .A1(AMVG3VG1VAD2NF), .A2(AMVG3VG1VAD1NF) );
  NOR2_X1 NOR2_7( .ZN(AMVG2VX), .A1(AMVG2VG1VAD2NF), .A2(AMVG2VG1VAD1NF) );
  NOR2_X1 NOR2_8( .ZN(BMVG5VX), .A1(BMVG5VG1VAD2NF), .A2(BMVG5VG1VAD1NF) );
  NOR2_X1 NOR2_9( .ZN(BMVG4VX), .A1(BMVG4VG1VAD2NF), .A2(BMVG4VG1VAD1NF) );
  NOR2_X1 NOR2_10( .ZN(BMVG3VX), .A1(BMVG3VG1VAD2NF), .A2(BMVG3VG1VAD1NF) );
  NOR2_X1 NOR2_11( .ZN(BMVG2VX), .A1(BMVG2VG1VAD2NF), .A2(BMVG2VG1VAD1NF) );
  NOR2_X1 NOR2_12( .ZN(CNTVG3VD), .A1(CNTVG3VZ), .A2(START) );
  NOR2_X1 NOR2_13( .ZN(CNTVG2VD), .A1(CNTVG2VZ), .A2(START) );
  NOR2_X1 NOR2_14( .ZN(CNTVG1VD), .A1(CNTVG1VZ), .A2(START) );
  NOR2_X1 NOR2_15( .ZN(ADDVG2VCN), .A1(ADDVG2VCNVAD2NF), .A2(ADDVG2VCNVAD1NF) );
  NOR2_X1 NOR2_16( .ZN(MRVG4VD), .A1(MRVG4VDVAD2NF), .A2(MRVG4VDVAD1NF) );
  NOR2_X1 NOR2_17( .ZN(MRVG3VD), .A1(MRVG3VDVAD2NF), .A2(MRVG3VDVAD1NF) );
  NOR2_X2 NOR2_18( .ZN(MRVG2VD), .A1(MRVG2VDVAD2NF), .A2(MRVG2VDVAD1NF) );
  NOR2_X2 NOR2_19( .ZN(MRVG1VD), .A1(MRVG1VDVAD2NF), .A2(MRVG1VDVAD1NF) );
  NOR2_X2 NOR2_20( .ZN(ADDVG2VSN), .A1(ADDVG2VCNVAD4NF), .A2(ADDVG2VCNVAD3NF) );
  NOR2_X2 NOR2_21( .ZN(ADDVG3VCN), .A1(ADDVG3VCNVAD2NF), .A2(ADDVG3VCNVAD1NF) );
  NOR2_X1 NOR2_22( .ZN(ADDVG3VSN), .A1(ADDVG3VCNVAD4NF), .A2(ADDVG3VCNVAD3NF) );
  NOR2_X1 NOR2_23( .ZN(SMVG2VX), .A1(SMVG2VG1VAD2NF), .A2(SMVG2VG1VAD1NF) );
  NOR2_X1 NOR2_24( .ZN(ADDVG4VCN), .A1(ADDVG4VCNVAD2NF), .A2(ADDVG4VCNVAD1NF) );
  NOR2_X1 NOR2_25( .ZN(ADDVG4VSN), .A1(ADDVG4VCNVAD4NF), .A2(ADDVG4VCNVAD3NF) );
  NOR2_X1 NOR2_26( .ZN(SMVG3VX), .A1(SMVG3VG1VAD2NF), .A2(SMVG3VG1VAD1NF) );
  NOR2_X1 NOR2_27( .ZN(SMVG5VX), .A1(SMVG5VG1VAD2NF), .A2(SMVG5VG1VAD1NF) );
  NOR2_X1 NOR2_28( .ZN(SMVG4VX), .A1(SMVG4VG1VAD2NF), .A2(SMVG4VG1VAD1NF) );

endmodule
