//# 35 inputs
//# 24 outputs
//# 19 D-type flipflops
//# 272 inverters
//# 107 gates (90 ANDs + 4 NANDs + 13 ORs + 0 NORs)

module s641(CK,G1,G10,G100BF,G101BF,G103BF,G104BF,G105BF,G106BF,G107,G11,G12,G13,G138,G14,G15,
  G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,
  G32,G33,G34,G35,G36,G4,G5,G6,G8,G83,G84,G85,G86BF,G87BF,G88BF,G89BF,G9,G90,
  G91,G92,G94,G95BF,G96BF,G97BF,G98BF,G99BF);
input CK,G1,G2,G3,G4,G5,G6,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,
  G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36;
output G91,G94,G107,G83,G84,G85,G100BF,G98BF,G96BF,G92,G87BF,G89BF,G101BF,G106BF,G97BF,G104BF,G88BF,G99BF,G105BF,G138,
  G86BF,G95BF,G103BF,G90;

  wire G64,G380,G65,G262,G66,G394,G67,G250,G68,G122,G69,G133,G70,G71,G139,G72,
    G140,G73,G141,G74,G142,G75,G125,G76,G126,G77,G127,G78,G128,G79,G129,G80,
    G130,G81,G131,G82,G132,IIII633,G366,G379,IIII643,IIII646,IIII649,IIII652,IIII655,IIII660,IIII680,IIII684,
    IIII687,II165,IIII178,II169,II172,II175,II178,II181,II184,II187,II190,II193,II196,II199,II202,II205,
    II208,II211,G352,G360,G361,G362,G363,G364,G367,G386,G388,G389,G113,G115,G117,G219,
    G119,G221,G121,G223,G209,G109,G211,G111,G213,G215,G217,G110,G114,G118,G216,G218,
    G220,G222,G365,G368,G387,G225,G390,IIII356,G289,II254,G324,II257,II260,G338,II263,II266,
    G344,II269,II272,G312,II275,G315,II278,G318,II281,G321,G143,G166,G325,G194,G339,G202,
    G345,G313,G316,G319,G322,II303,IIII299,G281,IIII313,G283,II287,II291,II295,G350,IIII301,IIII315,
    G381,G100,G375,G98,G371,G96,G135,G137,G382,G376,G372,II321,II324,G329,G333,G87,
    IIII406,G89,IIII422,G173,G183,II335,II338,G174,G184,II341,G359,G355,G108,G356,G116,II354,
    G293,II357,II360,G309,II363,G146,G294,G162,G310,II366,G341,II369,II372,G303,II375,II378,
    II382,G198,G342,G154,G304,G383,G101,G396,G106,II386,II390,G384,G397,G373,G97,G392,
    G104,IIII476,IIII279,G278,G374,G393,G224,IIII306,G282,II373,G237,G286,IIII208,IIII308,IIII334,IIII327,
    G285,IIII210,G136,IIII336,IIII329,II442,G331,G88,IIII414,G178,II449,G179,II452,G357,G358,G112,
    II460,G335,II463,II466,G306,II469,G190,G336,G158,G307,II472,II476,G395,G377,G99,IIII272,
    G277,G105,G378,IIII265,G276,IIII292,G280,II440,G235,G284,IIII294,IIII320,IIII285,G279,G134,IIII322,
    IIII287,II517,G327,G86,IIII398,G168,II524,G169,II527,G353,G354,G120,II535,G347,II538,II541,
    G300,II544,G206,G348,G150,G301,II547,II551,G391,G369,G95,G103,G370,IIII258,G275,IIII230,
    G271,II511,G239,G288,IIII237,G272,IIII244,G273,IIII251,G274,IIII348,IIII341,G287,IIII222,G270,IIII350,
    IIII343,IIII224,G124,II608,G298,G231,G232,G233,G234,G247,G248,G263,G264,G214,G210,G266,
    G229,G245,G249,IIII533,G227,G243,G265,G236,G252,IIII527,G212,G228,G244,IIII515,G261,IIII512,
    IIII538,G256,G230,G246,G208,G226,G242,IIII553,IIII518,IIII521,IIII524,IIII495,G257,IIII537,G258,G259,
    G260,G241,G267,G238,G254,IIII546;

  DFF_X2 DFF_0( .CK(CK), .Q(G64), .D(G380) );
  DFF_X2 DFF_1( .CK(CK), .Q(G65), .D(G262) );
  DFF_X1 DFF_2( .CK(CK), .Q(G66), .D(G394) );
  DFF_X1 DFF_3( .CK(CK), .Q(G67), .D(G250) );
  DFF_X1 DFF_4( .CK(CK), .Q(G68), .D(G122) );
  DFF_X1 DFF_5( .CK(CK), .Q(G69), .D(G133) );
  DFF_X1 DFF_6( .CK(CK), .Q(G70), .D(G138) );
  DFF_X1 DFF_7( .CK(CK), .Q(G71), .D(G139) );
  DFF_X1 DFF_8( .CK(CK), .Q(G72), .D(G140) );
  DFF_X1 DFF_9( .CK(CK), .Q(G73), .D(G141) );
  DFF_X1 DFF_10( .CK(CK), .Q(G74), .D(G142) );
  DFF_X1 DFF_11( .CK(CK), .Q(G75), .D(G125) );
  DFF_X1 DFF_12( .CK(CK), .Q(G76), .D(G126) );
  DFF_X1 DFF_13( .CK(CK), .Q(G77), .D(G127) );
  DFF_X1 DFF_14( .CK(CK), .Q(G78), .D(G128) );
  DFF_X1 DFF_15( .CK(CK), .Q(G79), .D(G129) );
  DFF_X1 DFF_16( .CK(CK), .Q(G80), .D(G130) );
  DFF_X1 DFF_17( .CK(CK), .Q(G81), .D(G131) );
  DFF_X2 DFF_18( .CK(CK), .Q(G82), .D(G132) );
  INV_X1 NOT_0( .ZN(IIII633), .A(G1) );
  INV_X1 NOT_1( .ZN(G366), .A(G2) );
  INV_X1 NOT_2( .ZN(G379), .A(G3) );
  INV_X1 NOT_3( .ZN(IIII643), .A(G4) );
  INV_X1 NOT_4( .ZN(IIII646), .A(G5) );
  INV_X1 NOT_5( .ZN(IIII649), .A(G6) );
  INV_X1 NOT_6( .ZN(IIII652), .A(G8) );
  INV_X1 NOT_7( .ZN(IIII655), .A(G9) );
  INV_X1 NOT_8( .ZN(IIII660), .A(G10) );
  INV_X1 NOT_9( .ZN(IIII680), .A(G11) );
  INV_X1 NOT_10( .ZN(IIII684), .A(G12) );
  INV_X1 NOT_11( .ZN(IIII687), .A(G13) );
  INV_X1 NOT_12( .ZN(II165), .A(G27) );
  INV_X1 NOT_13( .ZN(IIII178), .A(G29) );
  INV_X1 NOT_14( .ZN(II169), .A(G70) );
  INV_X1 NOT_15( .ZN(II172), .A(G71) );
  INV_X1 NOT_16( .ZN(II175), .A(G72) );
  INV_X1 NOT_17( .ZN(II178), .A(G80) );
  INV_X1 NOT_18( .ZN(II181), .A(G73) );
  INV_X1 NOT_19( .ZN(II184), .A(G81) );
  INV_X1 NOT_20( .ZN(II187), .A(G74) );
  INV_X1 NOT_21( .ZN(II190), .A(G82) );
  INV_X1 NOT_22( .ZN(II193), .A(G75) );
  INV_X1 NOT_23( .ZN(II196), .A(G68) );
  INV_X2 NOT_24( .ZN(II199), .A(G76) );
  INV_X2 NOT_25( .ZN(II202), .A(G69) );
  INV_X1 NOT_26( .ZN(II205), .A(G77) );
  INV_X1 NOT_27( .ZN(II208), .A(G78) );
  INV_X1 NOT_28( .ZN(II211), .A(G79) );
  INV_X1 NOT_29( .ZN(G352), .A(IIII633) );
  INV_X1 NOT_30( .ZN(G360), .A(IIII643) );
  INV_X1 NOT_31( .ZN(G361), .A(IIII646) );
  INV_X1 NOT_32( .ZN(G362), .A(IIII649) );
  INV_X1 NOT_33( .ZN(G363), .A(IIII652) );
  INV_X1 NOT_34( .ZN(G364), .A(IIII655) );
  INV_X1 NOT_35( .ZN(G367), .A(IIII660) );
  INV_X1 NOT_36( .ZN(G386), .A(IIII680) );
  INV_X1 NOT_37( .ZN(G388), .A(IIII684) );
  INV_X1 NOT_38( .ZN(G389), .A(IIII687) );
  INV_X1 NOT_39( .ZN(G91), .A(II165) );
  INV_X1 NOT_40( .ZN(G94), .A(IIII178) );
  INV_X8 NOT_41( .ZN(G113), .A(II169) );
  INV_X1 NOT_42( .ZN(G115), .A(II172) );
  INV_X1 NOT_43( .ZN(G117), .A(II175) );
  INV_X1 NOT_44( .ZN(G219), .A(II178) );
  INV_X1 NOT_45( .ZN(G119), .A(II181) );
  INV_X1 NOT_46( .ZN(G221), .A(II184) );
  INV_X1 NOT_47( .ZN(G121), .A(II187) );
  INV_X1 NOT_48( .ZN(G223), .A(II190) );
  INV_X1 NOT_49( .ZN(G209), .A(II193) );
  INV_X1 NOT_50( .ZN(G109), .A(II196) );
  INV_X1 NOT_51( .ZN(G211), .A(II199) );
  INV_X1 NOT_52( .ZN(G111), .A(II202) );
  INV_X1 NOT_53( .ZN(G213), .A(II205) );
  INV_X4 NOT_54( .ZN(G215), .A(II208) );
  INV_X1 NOT_55( .ZN(G217), .A(II211) );
  INV_X1 NOT_56( .ZN(G110), .A(G360) );
  INV_X1 NOT_57( .ZN(G114), .A(G360) );
  INV_X1 NOT_58( .ZN(G118), .A(G360) );
  INV_X1 NOT_59( .ZN(G216), .A(G360) );
  INV_X1 NOT_60( .ZN(G218), .A(G360) );
  INV_X1 NOT_61( .ZN(G220), .A(G360) );
  INV_X1 NOT_62( .ZN(G222), .A(G360) );
  INV_X1 NOT_63( .ZN(G365), .A(G364) );
  INV_X1 NOT_64( .ZN(G368), .A(G367) );
  INV_X1 NOT_65( .ZN(G387), .A(G386) );
  INV_X1 NOT_66( .ZN(G225), .A(G388) );
  INV_X1 NOT_67( .ZN(G390), .A(G389) );
  INV_X1 NOT_68( .ZN(IIII356), .A(G289) );
  INV_X1 NOT_69( .ZN(II254), .A(G324) );
  INV_X1 NOT_70( .ZN(II257), .A(G324) );
  INV_X1 NOT_71( .ZN(II260), .A(G338) );
  INV_X1 NOT_72( .ZN(II263), .A(G338) );
  INV_X1 NOT_73( .ZN(II266), .A(G344) );
  INV_X1 NOT_74( .ZN(II269), .A(G344) );
  INV_X1 NOT_75( .ZN(II272), .A(G312) );
  INV_X2 NOT_76( .ZN(II275), .A(G315) );
  INV_X1 NOT_77( .ZN(II278), .A(G318) );
  INV_X1 NOT_78( .ZN(II281), .A(G321) );
  INV_X1 NOT_79( .ZN(G143), .A(IIII356) );
  INV_X1 NOT_80( .ZN(G166), .A(II254) );
  INV_X1 NOT_81( .ZN(G325), .A(II257) );
  INV_X1 NOT_82( .ZN(G194), .A(II260) );
  INV_X1 NOT_83( .ZN(G339), .A(II263) );
  INV_X1 NOT_84( .ZN(G202), .A(II266) );
  INV_X1 NOT_85( .ZN(G345), .A(II269) );
  INV_X1 NOT_86( .ZN(G313), .A(II272) );
  INV_X1 NOT_87( .ZN(G316), .A(II275) );
  INV_X1 NOT_88( .ZN(G319), .A(II278) );
  INV_X1 NOT_89( .ZN(G322), .A(II281) );
  INV_X1 NOT_90( .ZN(II303), .A(G143) );
  INV_X1 NOT_91( .ZN(IIII299), .A(G281) );
  INV_X32 NOT_92( .ZN(IIII313), .A(G283) );
  INV_X1 NOT_93( .ZN(II287), .A(G166) );
  INV_X1 NOT_94( .ZN(II291), .A(G194) );
  INV_X1 NOT_95( .ZN(II295), .A(G202) );
  INV_X1 NOT_96( .ZN(G350), .A(II303) );
  INV_X1 NOT_97( .ZN(IIII301), .A(IIII299) );
  INV_X1 NOT_98( .ZN(IIII315), .A(IIII313) );
  INV_X8 NOT_99( .ZN(G381), .A(II287) );
  INV_X1 NOT_100( .ZN(G100BF), .A(G100) );
  INV_X1 NOT_101( .ZN(G375), .A(II291) );
  INV_X1 NOT_102( .ZN(G98BF), .A(G98) );
  INV_X1 NOT_103( .ZN(G371), .A(II295) );
  INV_X1 NOT_104( .ZN(G96BF), .A(G96) );
  INV_X1 NOT_105( .ZN(G135), .A(IIII301) );
  INV_X1 NOT_106( .ZN(G137), .A(IIII315) );
  INV_X1 NOT_107( .ZN(G382), .A(G381) );
  INV_X1 NOT_108( .ZN(G376), .A(G375) );
  INV_X1 NOT_109( .ZN(G372), .A(G371) );
  INV_X1 NOT_110( .ZN(II321), .A(G135) );
  INV_X1 NOT_111( .ZN(II324), .A(G137) );
  INV_X1 NOT_112( .ZN(G329), .A(II321) );
  INV_X1 NOT_113( .ZN(G333), .A(II324) );
  INV_X1 NOT_114( .ZN(G87BF), .A(G87) );
  INV_X1 NOT_115( .ZN(IIII406), .A(G87) );
  INV_X1 NOT_116( .ZN(G89BF), .A(G89) );
  INV_X1 NOT_117( .ZN(IIII422), .A(G89) );
  INV_X1 NOT_118( .ZN(G173), .A(IIII406) );
  INV_X1 NOT_119( .ZN(G183), .A(IIII422) );
  INV_X1 NOT_120( .ZN(II335), .A(G173) );
  INV_X1 NOT_121( .ZN(II338), .A(G183) );
  INV_X1 NOT_122( .ZN(G174), .A(II335) );
  INV_X1 NOT_123( .ZN(G184), .A(II338) );
  INV_X1 NOT_124( .ZN(II341), .A(G174) );
  INV_X2 NOT_125( .ZN(G359), .A(G184) );
  INV_X2 NOT_126( .ZN(G355), .A(II341) );
  INV_X2 NOT_127( .ZN(G108), .A(G359) );
  INV_X1 NOT_128( .ZN(G356), .A(G355) );
  INV_X1 NOT_129( .ZN(G116), .A(G356) );
  INV_X1 NOT_130( .ZN(II354), .A(G293) );
  INV_X1 NOT_131( .ZN(II357), .A(G293) );
  INV_X1 NOT_132( .ZN(II360), .A(G309) );
  INV_X1 NOT_133( .ZN(II363), .A(G309) );
  INV_X1 NOT_134( .ZN(G146), .A(II354) );
  INV_X1 NOT_135( .ZN(G294), .A(II357) );
  INV_X1 NOT_136( .ZN(G162), .A(II360) );
  INV_X1 NOT_137( .ZN(G310), .A(II363) );
  INV_X1 NOT_138( .ZN(II366), .A(G341) );
  INV_X1 NOT_139( .ZN(II369), .A(G341) );
  INV_X1 NOT_140( .ZN(II372), .A(G303) );
  INV_X1 NOT_141( .ZN(II375), .A(G303) );
  INV_X1 NOT_142( .ZN(II378), .A(G146) );
  INV_X1 NOT_143( .ZN(II382), .A(G162) );
  INV_X1 NOT_144( .ZN(G198), .A(II366) );
  INV_X1 NOT_145( .ZN(G342), .A(II369) );
  INV_X1 NOT_146( .ZN(G154), .A(II372) );
  INV_X1 NOT_147( .ZN(G304), .A(II375) );
  INV_X1 NOT_148( .ZN(G383), .A(II378) );
  INV_X1 NOT_149( .ZN(G101BF), .A(G101) );
  INV_X1 NOT_150( .ZN(G396), .A(II382) );
  INV_X4 NOT_151( .ZN(G106BF), .A(G106) );
  INV_X1 NOT_152( .ZN(II386), .A(G198) );
  INV_X1 NOT_153( .ZN(II390), .A(G154) );
  INV_X1 NOT_154( .ZN(G384), .A(G383) );
  INV_X1 NOT_155( .ZN(G397), .A(G396) );
  INV_X1 NOT_156( .ZN(G373), .A(II386) );
  INV_X1 NOT_157( .ZN(G97BF), .A(G97) );
  INV_X1 NOT_158( .ZN(G392), .A(II390) );
  INV_X1 NOT_159( .ZN(G104BF), .A(G104) );
  INV_X1 NOT_160( .ZN(IIII476), .A(G384) );
  INV_X1 NOT_161( .ZN(IIII279), .A(G278) );
  INV_X1 NOT_162( .ZN(G374), .A(G373) );
  INV_X1 NOT_163( .ZN(G393), .A(G392) );
  INV_X1 NOT_164( .ZN(G224), .A(IIII476) );
  INV_X1 NOT_165( .ZN(G132), .A(IIII279) );
  INV_X1 NOT_166( .ZN(IIII306), .A(G282) );
  INV_X1 NOT_167( .ZN(II373), .A(G237) );
  INV_X1 NOT_168( .ZN(G286), .A(II373) );
  INV_X1 NOT_169( .ZN(IIII208), .A(G224) );
  INV_X1 NOT_170( .ZN(IIII308), .A(IIII306) );
  INV_X1 NOT_171( .ZN(IIII334), .A(G286) );
  INV_X1 NOT_172( .ZN(IIII327), .A(G285) );
  INV_X8 NOT_173( .ZN(IIII210), .A(IIII208) );
  INV_X8 NOT_174( .ZN(G136), .A(IIII308) );
  INV_X1 NOT_175( .ZN(IIII336), .A(IIII334) );
  INV_X1 NOT_176( .ZN(IIII329), .A(IIII327) );
  INV_X1 NOT_177( .ZN(G122), .A(IIII210) );
  INV_X1 NOT_178( .ZN(II442), .A(G136) );
  INV_X1 NOT_179( .ZN(G140), .A(IIII336) );
  INV_X1 NOT_180( .ZN(G139), .A(IIII329) );
  INV_X1 NOT_181( .ZN(G331), .A(II442) );
  INV_X1 NOT_182( .ZN(G88BF), .A(G88) );
  INV_X1 NOT_183( .ZN(IIII414), .A(G88) );
  INV_X1 NOT_184( .ZN(G178), .A(IIII414) );
  INV_X1 NOT_185( .ZN(II449), .A(G178) );
  INV_X1 NOT_186( .ZN(G179), .A(II449) );
  INV_X1 NOT_187( .ZN(II452), .A(G179) );
  INV_X1 NOT_188( .ZN(G357), .A(II452) );
  INV_X1 NOT_189( .ZN(G358), .A(G357) );
  INV_X1 NOT_190( .ZN(G112), .A(G358) );
  INV_X1 NOT_191( .ZN(II460), .A(G335) );
  INV_X1 NOT_192( .ZN(II463), .A(G335) );
  INV_X1 NOT_193( .ZN(II466), .A(G306) );
  INV_X1 NOT_194( .ZN(II469), .A(G306) );
  INV_X1 NOT_195( .ZN(G190), .A(II460) );
  INV_X1 NOT_196( .ZN(G336), .A(II463) );
  INV_X1 NOT_197( .ZN(G158), .A(II466) );
  INV_X1 NOT_198( .ZN(G307), .A(II469) );
  INV_X1 NOT_199( .ZN(II472), .A(G190) );
  INV_X4 NOT_200( .ZN(II476), .A(G158) );
  INV_X1 NOT_201( .ZN(G395), .A(G158) );
  INV_X1 NOT_202( .ZN(G377), .A(II472) );
  INV_X1 NOT_203( .ZN(G99BF), .A(G99) );
  INV_X1 NOT_204( .ZN(G394), .A(II476) );
  INV_X4 NOT_205( .ZN(IIII272), .A(G277) );
  INV_X1 NOT_206( .ZN(G105BF), .A(G105) );
  INV_X1 NOT_207( .ZN(G378), .A(G377) );
  INV_X1 NOT_208( .ZN(G131), .A(IIII272) );
  INV_X1 NOT_209( .ZN(IIII265), .A(G276) );
  INV_X1 NOT_210( .ZN(IIII292), .A(G280) );
  INV_X1 NOT_211( .ZN(G130), .A(IIII265) );
  INV_X1 NOT_212( .ZN(II440), .A(G235) );
  INV_X1 NOT_213( .ZN(G284), .A(II440) );
  INV_X1 NOT_214( .ZN(IIII294), .A(IIII292) );
  INV_X1 NOT_215( .ZN(IIII320), .A(G284) );
  INV_X1 NOT_216( .ZN(IIII285), .A(G279) );
  INV_X1 NOT_217( .ZN(G134), .A(IIII294) );
  INV_X1 NOT_218( .ZN(IIII322), .A(IIII320) );
  INV_X1 NOT_219( .ZN(IIII287), .A(IIII285) );
  INV_X1 NOT_220( .ZN(II517), .A(G134) );
  INV_X1 NOT_221( .ZN(G138), .A(IIII322) );
  INV_X1 NOT_222( .ZN(G133), .A(IIII287) );
  INV_X1 NOT_223( .ZN(G327), .A(II517) );
  INV_X1 NOT_224( .ZN(G86BF), .A(G86) );
  INV_X1 NOT_225( .ZN(IIII398), .A(G86) );
  INV_X1 NOT_226( .ZN(G168), .A(IIII398) );
  INV_X1 NOT_227( .ZN(II524), .A(G168) );
  INV_X1 NOT_228( .ZN(G169), .A(II524) );
  INV_X1 NOT_229( .ZN(II527), .A(G169) );
  INV_X1 NOT_230( .ZN(G353), .A(II527) );
  INV_X1 NOT_231( .ZN(G354), .A(G353) );
  INV_X1 NOT_232( .ZN(G120), .A(G354) );
  INV_X1 NOT_233( .ZN(II535), .A(G347) );
  INV_X1 NOT_234( .ZN(II538), .A(G347) );
  INV_X1 NOT_235( .ZN(II541), .A(G300) );
  INV_X8 NOT_236( .ZN(II544), .A(G300) );
  INV_X8 NOT_237( .ZN(G206), .A(II535) );
  INV_X8 NOT_238( .ZN(G348), .A(II538) );
  INV_X1 NOT_239( .ZN(G150), .A(II541) );
  INV_X1 NOT_240( .ZN(G301), .A(II544) );
  INV_X1 NOT_241( .ZN(II547), .A(G206) );
  INV_X1 NOT_242( .ZN(II551), .A(G150) );
  INV_X1 NOT_243( .ZN(G391), .A(G150) );
  INV_X1 NOT_244( .ZN(G369), .A(II547) );
  INV_X1 NOT_245( .ZN(G95BF), .A(G95) );
  INV_X1 NOT_246( .ZN(G380), .A(II551) );
  INV_X1 NOT_247( .ZN(G103BF), .A(G103) );
  INV_X1 NOT_248( .ZN(G370), .A(G369) );
  INV_X1 NOT_249( .ZN(IIII258), .A(G275) );
  INV_X1 NOT_250( .ZN(G129), .A(IIII258) );
  INV_X1 NOT_251( .ZN(IIII230), .A(G271) );
  INV_X1 NOT_252( .ZN(II511), .A(G239) );
  INV_X1 NOT_253( .ZN(G288), .A(II511) );
  INV_X1 NOT_254( .ZN(IIII237), .A(G272) );
  INV_X1 NOT_255( .ZN(IIII244), .A(G273) );
  INV_X1 NOT_256( .ZN(IIII251), .A(G274) );
  INV_X1 NOT_257( .ZN(G125), .A(IIII230) );
  INV_X1 NOT_258( .ZN(IIII348), .A(G288) );
  INV_X1 NOT_259( .ZN(IIII341), .A(G287) );
  INV_X1 NOT_260( .ZN(G126), .A(IIII237) );
  INV_X1 NOT_261( .ZN(G127), .A(IIII244) );
  INV_X1 NOT_262( .ZN(G128), .A(IIII251) );
  INV_X1 NOT_263( .ZN(IIII222), .A(G270) );
  INV_X1 NOT_264( .ZN(IIII350), .A(IIII348) );
  INV_X1 NOT_265( .ZN(IIII343), .A(IIII341) );
  INV_X1 NOT_266( .ZN(IIII224), .A(IIII222) );
  INV_X1 NOT_267( .ZN(G142), .A(IIII350) );
  INV_X1 NOT_268( .ZN(G141), .A(IIII343) );
  INV_X1 NOT_269( .ZN(G124), .A(IIII224) );
  INV_X1 NOT_270( .ZN(II608), .A(G124) );
  INV_X1 NOT_271( .ZN(G298), .A(II608) );
  AND3_X1 AND3_0( .ZN(G289), .A1(G386), .A2(G388), .A3(G389) );
  AND2_X1 AND2_0( .ZN(G324), .A1(G110), .A2(G111) );
  AND2_X1 AND2_1( .ZN(G338), .A1(G114), .A2(G115) );
  AND2_X1 AND2_2( .ZN(G344), .A1(G118), .A2(G119) );
  AND2_X1 AND2_3( .ZN(G312), .A1(G216), .A2(G217) );
  AND2_X1 AND2_4( .ZN(G315), .A1(G218), .A2(G219) );
  AND2_X1 AND2_5( .ZN(G318), .A1(G220), .A2(G221) );
  AND2_X1 AND2_6( .ZN(G321), .A1(G222), .A2(G223) );
  AND2_X1 AND2_7( .ZN(G231), .A1(G379), .A2(G387) );
  AND2_X1 AND2_8( .ZN(G232), .A1(G379), .A2(G387) );
  AND2_X1 AND2_9( .ZN(G233), .A1(G379), .A2(G387) );
  AND2_X1 AND2_10( .ZN(G234), .A1(G379), .A2(G387) );
  AND4_X1 AND4_0( .ZN(G247), .A1(G379), .A2(G365), .A3(G368), .A4(G390) );
  AND4_X1 AND4_1( .ZN(G248), .A1(G379), .A2(G365), .A3(G367), .A4(G390) );
  AND4_X1 AND4_2( .ZN(G263), .A1(G379), .A2(G364), .A3(G368), .A4(G390) );
  AND4_X2 AND4_3( .ZN(G264), .A1(G379), .A2(G364), .A3(G367), .A4(G390) );
  AND2_X2 AND2_11( .ZN(G100), .A1(G325), .A2(G35) );
  AND2_X2 AND2_12( .ZN(G98), .A1(G339), .A2(G33) );
  AND2_X1 AND2_13( .ZN(G96), .A1(G345), .A2(G31) );
  AND2_X1 AND2_14( .ZN(G107), .A1(G313), .A2(G18) );
  AND2_X1 AND2_15( .ZN(G83), .A1(G316), .A2(G19) );
  AND2_X1 AND2_16( .ZN(G84), .A1(G319), .A2(G20) );
  AND2_X1 AND2_17( .ZN(G85), .A1(G322), .A2(G21) );
  AND2_X1 AND2_18( .ZN(G92), .A1(G350), .A2(G28) );
  AND2_X1 AND2_19( .ZN(G87), .A1(G329), .A2(G23) );
  AND2_X1 AND2_20( .ZN(G89), .A1(G333), .A2(G25) );
  AND2_X1 AND2_21( .ZN(G293), .A1(G108), .A2(G109) );
  AND2_X1 AND2_22( .ZN(G309), .A1(G214), .A2(G215) );
  AND2_X1 AND2_23( .ZN(G341), .A1(G116), .A2(G117) );
  AND2_X1 AND2_24( .ZN(G303), .A1(G210), .A2(G211) );
  AND2_X1 AND2_25( .ZN(G101), .A1(G294), .A2(G36) );
  AND2_X1 AND2_26( .ZN(G106), .A1(G310), .A2(G17) );
  AND2_X1 AND2_27( .ZN(G97), .A1(G342), .A2(G32) );
  AND2_X1 AND2_28( .ZN(G104), .A1(G304), .A2(G15) );
  AND4_X1 AND4_4( .ZN(G266), .A1(G364), .A2(G367), .A3(G383), .A4(G390) );
  AND2_X1 AND2_29( .ZN(G229), .A1(G366), .A2(G396) );
  AND2_X1 AND2_30( .ZN(G245), .A1(G352), .A2(G396) );
  AND2_X1 AND2_31( .ZN(G250), .A1(G366), .A2(G396) );
  AND2_X1 AND2_32( .ZN(G278), .A1(G366), .A2(G396) );
  AND3_X1 AND3_1( .ZN(G249), .A1(G366), .A2(G66), .A3(G397) );
  AND3_X1 AND3_2( .ZN(IIII533), .A1(G365), .A2(G367), .A3(G373) );
  AND2_X1 AND2_33( .ZN(G227), .A1(G366), .A2(G392) );
  AND2_X2 AND2_34( .ZN(G243), .A1(G392), .A2(G361) );
  AND3_X1 AND3_3( .ZN(G265), .A1(G375), .A2(G390), .A3(IIII533) );
  AND2_X1 AND2_35( .ZN(G236), .A1(G374), .A2(G376) );
  AND2_X1 AND2_36( .ZN(G237), .A1(G374), .A2(G375) );
  AND2_X1 AND2_37( .ZN(G252), .A1(G355), .A2(G374) );
  AND3_X1 AND3_4( .ZN(IIII527), .A1(G366), .A2(G64), .A3(G393) );
  AND2_X1 AND2_38( .ZN(G88), .A1(G331), .A2(G24) );
  AND2_X1 AND2_39( .ZN(G335), .A1(G112), .A2(G113) );
  AND2_X1 AND2_40( .ZN(G306), .A1(G212), .A2(G213) );
  AND2_X1 AND2_41( .ZN(G99), .A1(G336), .A2(G34) );
  AND2_X1 AND2_42( .ZN(G228), .A1(G366), .A2(G158) );
  AND2_X1 AND2_43( .ZN(G244), .A1(G158), .A2(G362) );
  AND3_X1 AND3_5( .ZN(G277), .A1(G366), .A2(G158), .A3(G397) );
  AND2_X1 AND2_44( .ZN(G105), .A1(G307), .A2(G16) );
  AND3_X1 AND3_6( .ZN(IIII515), .A1(G393), .A2(G395), .A3(G397) );
  AND3_X1 AND3_7( .ZN(G261), .A1(G395), .A2(G397), .A3(IIII527) );
  AND4_X1 AND4_5( .ZN(G262), .A1(G366), .A2(G392), .A3(G395), .A4(G397) );
  AND4_X1 AND4_6( .ZN(G276), .A1(G366), .A2(G392), .A3(G395), .A4(G397) );
  AND3_X1 AND3_8( .ZN(IIII512), .A1(G364), .A2(G368), .A3(G377) );
  AND4_X1 AND4_7( .ZN(IIII538), .A1(G377), .A2(G381), .A3(G383), .A4(G387) );
  AND3_X1 AND3_9( .ZN(G256), .A1(G381), .A2(G390), .A3(IIII512) );
  AND2_X1 AND2_45( .ZN(G230), .A1(G378), .A2(G382) );
  AND2_X1 AND2_46( .ZN(G235), .A1(G378), .A2(G381) );
  AND2_X1 AND2_47( .ZN(G246), .A1(G357), .A2(G378) );
  AND2_X1 AND2_48( .ZN(G86), .A1(G327), .A2(G22) );
  AND2_X1 AND2_49( .ZN(G347), .A1(G120), .A2(G121) );
  AND2_X1 AND2_50( .ZN(G300), .A1(G208), .A2(G209) );
  AND2_X1 AND2_51( .ZN(G95), .A1(G348), .A2(G30) );
  AND2_X1 AND2_52( .ZN(G226), .A1(G366), .A2(G150) );
  AND2_X1 AND2_53( .ZN(G242), .A1(G150), .A2(G363) );
  AND3_X1 AND3_10( .ZN(IIII553), .A1(G366), .A2(G150), .A3(G393) );
  AND2_X1 AND2_54( .ZN(G103), .A1(G301), .A2(G14) );
  AND3_X4 AND3_11( .ZN(G275), .A1(G395), .A2(G397), .A3(IIII553) );
  AND3_X2 AND3_12( .ZN(IIII518), .A1(G391), .A2(G395), .A3(G397) );
  AND3_X2 AND3_13( .ZN(IIII521), .A1(G391), .A2(G393), .A3(G397) );
  AND3_X1 AND3_14( .ZN(IIII524), .A1(G352), .A2(G391), .A3(G393) );
  AND3_X1 AND3_15( .ZN(IIII495), .A1(G365), .A2(G368), .A3(G369) );
  AND4_X1 AND4_8( .ZN(G257), .A1(G363), .A2(G369), .A3(G371), .A4(IIII515) );
  AND4_X1 AND4_9( .ZN(IIII537), .A1(G369), .A2(G371), .A3(G373), .A4(G375) );
  AND4_X1 AND4_10( .ZN(G258), .A1(G361), .A2(G373), .A3(G375), .A4(IIII518) );
  AND4_X1 AND4_11( .ZN(G259), .A1(G362), .A2(G377), .A3(G381), .A4(IIII521) );
  AND3_X1 AND3_16( .ZN(G260), .A1(G395), .A2(G383), .A3(IIII524) );
  AND3_X1 AND3_17( .ZN(G241), .A1(G371), .A2(G390), .A3(IIII495) );
  AND2_X1 AND2_55( .ZN(G267), .A1(IIII537), .A2(IIII538) );
  AND2_X1 AND2_56( .ZN(G238), .A1(G370), .A2(G372) );
  AND2_X1 AND2_57( .ZN(G239), .A1(G370), .A2(G371) );
  AND2_X1 AND2_58( .ZN(G254), .A1(G353), .A2(G370) );
  AND2_X1 AND2_59( .ZN(G90), .A1(G298), .A2(G26) );
  OR3_X1 OR3_0( .ZN(G281), .A1(G232), .A2(G248), .A3(G65) );
  OR3_X1 OR3_1( .ZN(G283), .A1(G234), .A2(G67), .A3(G264) );
  OR3_X1 OR3_2( .ZN(G282), .A1(G233), .A2(G249), .A3(G263) );
  OR2_X1 OR2_0( .ZN(G285), .A1(G236), .A2(G252) );
  OR3_X1 OR3_3( .ZN(G280), .A1(G231), .A2(G247), .A3(G261) );
  OR2_X2 OR2_1( .ZN(G279), .A1(G230), .A2(G246) );
  OR3_X2 OR3_4( .ZN(G271), .A1(G226), .A2(G242), .A3(G257) );
  OR3_X1 OR3_5( .ZN(G272), .A1(G227), .A2(G243), .A3(G258) );
  OR3_X1 OR3_6( .ZN(G273), .A1(G228), .A2(G244), .A3(G259) );
  OR3_X1 OR3_7( .ZN(G274), .A1(G229), .A2(G245), .A3(G260) );
  OR3_X1 OR3_8( .ZN(IIII546), .A1(G225), .A2(G241), .A3(G256) );
  OR2_X1 OR2_2( .ZN(G287), .A1(G238), .A2(G254) );
  OR4_X1 OR4_0( .ZN(G270), .A1(G265), .A2(G266), .A3(G267), .A4(IIII546) );
  NAND2_X1 NAND2_0( .ZN(G214), .A1(G379), .A2(G359) );
  NAND2_X2 NAND2_1( .ZN(G210), .A1(G379), .A2(G356) );
  NAND2_X2 NAND2_2( .ZN(G212), .A1(G379), .A2(G358) );
  NAND2_X1 NAND2_3( .ZN(G208), .A1(G379), .A2(G354) );

endmodule
