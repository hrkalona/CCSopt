//# 35 inputs
//# 49 outputs
//# 179 D-type flipflops
//# 1775 inverters
//# 1004 gates (0 ANDs + 0 NANDs + 239 ORs + 765 NORs)

module s5378(CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,n3071gat,n3072gat,n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,
  n3080gat,n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,n3088gat,n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,n3097gat,n3098gat,
  n3099gat,n3100gat,n3104gat,n3105gat,n3106gat,n3107gat,n3108gat,n3109gat,n3110gat,n3111gat,n3112gat,n3113gat,n3114gat,n3115gat,n3116gat,n3117gat,n3118gat,n3119gat,
  n3120gat,n3121gat,n3122gat,n3123gat,n3124gat,n3125gat,n3126gat,n3127gat,n3128gat,n3129gat,n3130gat,n3131gat,n3132gat,n3133gat,n3134gat,n3135gat,n3136gat,n3137gat,
  n3138gat,n3139gat,n3140gat,n3141gat,n3142gat,n3143gat,n3144gat,n3145gat,n3146gat,n3147gat,n3148gat,n3149gat,n3150gat,n3151gat,n3152gat);
input CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,n3071gat,n3072gat,n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,n3080gat,n3081gat,
  n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,n3088gat,n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,n3097gat,n3098gat,n3099gat,n3100gat;
output n3104gat,n3105gat,n3106gat,n3107gat,n3108gat,n3109gat,n3110gat,n3111gat,n3112gat,n3113gat,n3114gat,n3115gat,n3116gat,n3117gat,n3118gat,n3119gat,n3120gat,n3121gat,n3122gat,n3123gat,
  n3124gat,n3125gat,n3126gat,n3127gat,n3128gat,n3129gat,n3130gat,n3131gat,n3132gat,n3133gat,n3134gat,n3135gat,n3136gat,n3137gat,n3138gat,n3139gat,n3140gat,n3141gat,n3142gat,n3143gat,
  n3144gat,n3145gat,n3146gat,n3147gat,n3148gat,n3149gat,n3150gat,n3151gat,n3152gat;

  wire n673gat,n2897gat,n398gat,n2782gat,n402gat,n2790gat,n919gat,n2670gat,n846gat,n2793gat,n394gat,n703gat,n722gat,n726gat,n2510gat,n748gat,
    n271gat,n2732gat,n160gat,n2776gat,n337gat,n2735gat,n842gat,n2673gat,n341gat,n2779gat,n2522gat,n43gat,n2472gat,n1620gat,n2319gat,n2470gat,
    n1821gat,n1827gat,n1825gat,n2029gat,n1816gat,n1829gat,n2027gat,n283gat,n165gat,n279gat,n1026gat,n275gat,n2476gat,n55gat,n1068gat,n2914gat,
    n957gat,n2928gat,n861gat,n2927gat,n1294gat,n2896gat,n1241gat,n2922gat,n1298gat,n865gat,n2894gat,n1080gat,n2921gat,n1148gat,n2895gat,n2468gat,
    n933gat,n618gat,n491gat,n622gat,n626gat,n834gat,n3064gat,n707gat,n3055gat,n838gat,n3063gat,n830gat,n3062gat,n614gat,n3056gat,n2526gat,
    n504gat,n680gat,n2913gat,n816gat,n2920gat,n580gat,n2905gat,n824gat,n3057gat,n820gat,n3059gat,n883gat,n3058gat,n584gat,n2898gat,n684gat,
    n3060gat,n699gat,n3061gat,n2464gat,n567gat,n2399gat,n3048gat,n2343gat,n3049gat,n2203gat,n3051gat,n2562gat,n3047gat,n2207gat,n3050gat,n2626gat,
    n3040gat,n2490gat,n3044gat,n2622gat,n3042gat,n2630gat,n3037gat,n2543gat,n3041gat,n2102gat,n1606gat,n1880gat,n3052gat,n1763gat,n1610gat,n2155gat,
    n1858gat,n1035gat,n2918gat,n1121gat,n2952gat,n1072gat,n2919gat,n1282gat,n2910gat,n1226gat,n2907gat,n931gat,n2911gat,n1135gat,n2912gat,n1045gat,
    n2909gat,n1197gat,n2908gat,n2518gat,n2971gat,n667gat,n2904gat,n659gat,n2891gat,n553gat,n2903gat,n777gat,n2915gat,n561gat,n2901gat,n366gat,
    n2890gat,n322gat,n2888gat,n318gat,n2887gat,n314gat,n2886gat,n2599gat,n3010gat,n2588gat,n3016gat,n2640gat,n3054gat,n2658gat,n2579gat,n2495gat,
    n3036gat,n2390gat,n3034gat,n2270gat,n3031gat,n2339gat,n3035gat,n2502gat,n2646gat,n2634gat,n3053gat,n2506gat,n2613gat,n1834gat,n1625gat,n1767gat,
    n1626gat,n2084gat,n1603gat,n2143gat,n2541gat,n2061gat,n2557gat,n2139gat,n2487gat,n1899gat,n2532gat,n1850gat,n2628gat,n2403gat,n2397gat,n2394gat,
    n2341gat,n2440gat,n2560gat,n2407gat,n2205gat,n2347gat,n2201gat,n1389gat,n1793gat,n2021gat,n1781gat,n1394gat,n1516gat,n1496gat,n1392gat,n2091gat,
    n1685gat,n1332gat,n1565gat,n1740gat,n1330gat,n2179gat,n1945gat,n2190gat,n2268gat,n2135gat,n2337gat,n2262gat,n2388gat,n2182gat,n1836gat,n1433gat,
    n2983gat,n1316gat,n1431gat,n1363gat,n1314gat,n1312gat,n1361gat,n1775gat,n1696gat,n1871gat,n2009gat,n2592gat,n1773gat,n1508gat,n1636gat,n1678gat,
    n1712gat,n2309gat,n3000gat,n2450gat,n2307gat,n2446gat,n2661gat,n2095gat,n827gat,n2176gat,n2093gat,n2169gat,n2174gat,n2454gat,n2163gat,n2040gat,
    n1777gat,n2044gat,n2015gat,n2037gat,n2042gat,n2025gat,n2017gat,n2099gat,n2023gat,n2266gat,n2493gat,n2033gat,n2035gat,n2110gat,n2031gat,n2125gat,
    n2108gat,n2121gat,n2123gat,n2117gat,n2119gat,n1975gat,n2632gat,n2644gat,n2638gat,n156gat,n612gat,n152gat,n705gat,n331gat,n822gat,n388gat,
    n881gat,n463gat,n818gat,n327gat,n682gat,n384gat,n697gat,n256gat,n836gat,n470gat,n828gat,n148gat,n832gat,n2458gat,n2590gat,n2514gat,
    n2456gat,n1771gat,n1613gat,n1336gat,n1391gat,n1748gat,n1927gat,n1675gat,n1713gat,n1807gat,n1717gat,n1340gat,n1567gat,n1456gat,n1564gat,n1525gat,
    n1632gat,n1462gat,n1915gat,n1596gat,n1800gat,n1588gat,n1593gat,II1,n2717gat,n2715gat,II5,n2725gat,n2723gat,n296gat,n421gat,II11,
    n2768gat,II14,n2767gat,n373gat,II18,n2671gat,n2669gat,II23,n2845gat,n2844gat,II27,n2668gat,II30,n2667gat,n856gat,II44,
    n672gat,II47,n2783gat,II50,n396gat,II62,n2791gat,II65,II76,n401gat,n1645gat,n1499gat,II81,II92,n918gat,n1553gat,
    n1616gat,II97,n2794gat,II100,II111,n845gat,n1559gat,n1614gat,n1643gat,n1641gat,n1651gat,n1642gat,n1562gat,n1556gat,n1560gat,n1557gat,
    n1640gat,n1639gat,n1566gat,n1605gat,n1554gat,n1555gat,n1722gat,n1558gat,n392gat,II149,n702gat,n1319gat,n1256gat,n720gat,II171,n725gat,
    n1447gat,n1117gat,n1627gat,n1618gat,II178,n721gat,n1380gat,n1114gat,n1628gat,n1621gat,n701gat,n1446gat,n1318gat,n1705gat,n1619gat,n1706gat,
    n1622gat,II192,n2856gat,n2854gat,II196,n1218gat,II199,n2861gat,n2859gat,II203,n1219gat,II206,n2864gat,n2862gat,II210,n1220gat,
    II214,n2860gat,II217,n1221gat,II220,n2863gat,II223,n1222gat,II227,n2855gat,II230,n1223gat,n640gat,n1213gat,II237,n753gat,
    II240,n2716gat,II243,n2869gat,n2867gat,II248,n2868gat,II253,n2906gat,n754gat,II256,n2724gat,II259,n2728gat,n2726gat,II264,
    n2727gat,n422gat,n2889gat,II270,n755gat,n747gat,II275,n756gat,II278,n757gat,II282,n758gat,n2508gat,II297,n2733gat,II300,
    II311,n270gat,II314,n263gat,II317,n2777gat,II320,II331,n159gat,II334,n264gat,II337,n2736gat,II340,II351,n336gat,
    II354,n265gat,n158gat,II359,n266gat,n335gat,II363,n267gat,n269gat,II368,n268gat,n41gat,n258gat,II375,n48gat,II378,
    n1018gat,II381,n2674gat,II384,II395,n841gat,II398,n1019gat,II401,n1020gat,n840gat,II406,n1021gat,II409,n1022gat,n724gat,
    II414,n1023gat,II420,n1013gat,n49gat,II423,n2780gat,II426,II437,n340gat,II440,n480gat,II443,n481gat,II446,n393gat,
    II449,n482gat,II453,n483gat,II456,n484gat,n339gat,II461,n485gat,n42gat,n475gat,II468,n50gat,n162gat,II473,n51gat,
    II476,n52gat,II480,n53gat,n2520gat,n1448gat,n1376gat,n1701gat,n1617gat,n1379gat,n1377gat,n1615gat,n1624gat,n1500gat,n1113gat,n1503gat,
    n1501gat,n1779gat,n1623gat,II509,n2730gat,II512,n2729gat,n2317gat,n1819gat,n1823gat,n1817gat,II572,n1828gat,II576,n2851gat,II579,
    n2850gat,II583,n2786gat,n2785gat,n92gat,n637gat,n529gat,n293gat,n361gat,II591,n2722gat,II594,n2721gat,n297gat,II606,n282gat,
    II609,n172gat,II620,n164gat,II623,n173gat,II634,n278gat,II637,n174gat,n163gat,II642,n175gat,n277gat,II646,n176gat,
    n281gat,II651,n177gat,n54gat,n167gat,II658,n60gat,II661,n911gat,II672,n1025gat,II675,n912gat,II678,n913gat,n1024gat,
    II683,n914gat,n917gat,II687,n915gat,n844gat,II692,n916gat,II698,n906gat,n61gat,II709,n274gat,II712,n348gat,II715,
    n349gat,II718,n397gat,II721,n350gat,n400gat,II726,n351gat,II729,n352gat,n273gat,II734,n353gat,n178gat,n343gat,II741,
    n62gat,n66gat,II746,n63gat,II749,n64gat,II753,n65gat,n2474gat,II768,n2832gat,II771,n2831gat,n2731gat,II776,n2719gat,
    n2718gat,II790,n1067gat,II793,n949gat,II796,n2839gat,n2838gat,n2775gat,II812,n956gat,II815,n950gat,II818,n2712gat,n2711gat,
    n2734gat,II834,n860gat,II837,n951gat,n955gat,II842,n952gat,n859gat,II846,n953gat,n1066gat,II851,n954gat,n857gat,n944gat,
    II858,n938gat,n2792gat,II863,n2847gat,n2846gat,II877,n1293gat,II880,n1233gat,n2672gat,II885,n2853gat,n2852gat,II899,n1240gat,
    II902,n1234gat,II913,n1297gat,II916,n1235gat,n1239gat,II921,n1236gat,n1296gat,II925,n1237gat,n1292gat,II930,n1238gat,II936,
    n1228gat,n939gat,n2778gat,II941,n2837gat,n2836gat,II955,n864gat,II958,n1055gat,n2789gat,II963,n2841gat,n2840gat,II977,n1079gat,
    II980,n1056gat,n2781gat,II985,n2843gat,n2842gat,II999,n1147gat,II1002,n1057gat,n1078gat,II1007,n1058gat,n1146gat,II1011,n1059gat,
    n863gat,II1016,n1060gat,n928gat,n1050gat,II1023,n940gat,n858gat,II1028,n941gat,II1031,n942gat,II1035,n943gat,n2466gat,n2720gat,
    n740gat,n2784gat,n743gat,n746gat,n294gat,n360gat,n374gat,n616gat,II1067,n501gat,n489gat,II1079,n502gat,II1082,n617gat,II1085,
    n499gat,II1088,n490gat,II1091,n500gat,n620gat,II1103,n738gat,n624gat,II1115,n737gat,II1118,n621gat,II1121,n733gat,II1124,
    n625gat,II1127,n735gat,II1138,n833gat,II1141,n714gat,II1152,n706gat,II1155,n715gat,II1166,n837gat,II1169,n716gat,II1174,
    n717gat,II1178,n718gat,II1183,n719gat,n515gat,n709gat,II1190,n509gat,II1201,n829gat,II1204,n734gat,II1209,n736gat,II1216,
    n728gat,n510gat,II1227,n613gat,II1230,n498gat,II1236,n503gat,n404gat,n493gat,II1243,n511gat,n405gat,II1248,n512gat,II1251,
    n513gat,II1255,n514gat,n2524gat,n17gat,n564gat,n79gat,n86gat,n219gat,n78gat,n563gat,II1278,n289gat,n179gat,n287gat,n188gat,
    n288gat,n72gat,n181gat,n111gat,n182gat,II1302,n679gat,II1305,n808gat,II1319,n815gat,II1322,n809gat,II1336,n579gat,II1339,
    n810gat,n814gat,II1344,n811gat,n578gat,II1348,n812gat,n678gat,II1353,n813gat,n677gat,n803gat,II1360,n572gat,II1371,n823gat,
    II1374,n591gat,II1385,n819gat,II1388,n592gat,II1399,n882gat,II1402,n593gat,II1407,n594gat,II1411,n595gat,II1416,n596gat,
    II1422,n586gat,n573gat,II1436,n583gat,II1439,n691gat,II1450,n683gat,II1453,n692gat,II1464,n698gat,II1467,n693gat,II1472,
    n694gat,II1476,n695gat,n582gat,II1481,n696gat,n456gat,n686gat,II1488,n574gat,n565gat,II1493,n575gat,II1496,n576gat,II1500,
    n577gat,n2462gat,n2665gat,II1516,n2596gat,n189gat,n286gat,n194gat,n187gat,n21gat,n15gat,II1538,n2398gat,n2353gat,II1550,n2342gat,
    n2284gat,n2354gat,n2356gat,n2214gat,n2286gat,II1585,n2624gat,II1606,n2489gat,II1617,n2621gat,n2533gat,n2534gat,II1630,n2629gat,n2486gat,
    n2429gat,n2432gat,n2430gat,II1655,n2101gat,n1693gat,II1667,n1879gat,n1698gat,n1934gat,n1543gat,II1683,n1762gat,n1673gat,n2989gat,II1698,
    n2154gat,n2488gat,II1703,n2625gat,n2530gat,n2531gat,II1708,n2542gat,n2482gat,n2426gat,n2480gat,n2153gat,n2355gat,II1719,n2561gat,n2443gat,
    n2289gat,II1724,n2148gat,II1734,n855gat,n759gat,II1749,n1034gat,II1752,n1189gat,n1075gat,II1766,n1120gat,II1769,n1190gat,n760gat,
    II1783,n1071gat,II1786,n1191gat,n1119gat,II1791,n1192gat,n1070gat,II1795,n1193gat,n1033gat,II1800,n1194gat,n1183gat,n1184gat,II1807,
    n1274gat,n644gat,n1280gat,n641gat,II1833,n1225gat,II1837,n1281gat,n1224gat,II1843,n2970gat,n1275gat,n761gat,II1857,n930gat,II1860,
    n1206gat,n762gat,II1874,n1134gat,II1877,n1207gat,n643gat,II1891,n1044gat,II1894,n1208gat,n1133gat,II1899,n1209gat,n1043gat,II1903,
    n1210gat,n929gat,II1908,n1211gat,n1268gat,n1201gat,II1915,n1276gat,n1329gat,II1920,n1277gat,II1923,n1278gat,II1927,n1279gat,n1284gat,
    n1269gat,n642gat,n1195gat,II1947,n1196gat,n2516gat,II1961,n3017gat,n851gat,n853gat,n1725gat,n664gat,n852gat,n854gat,II1981,n666gat,
    n368gat,II1996,n658gat,II1999,n784gat,n662gat,II2014,n552gat,II2017,n785gat,n661gat,II2032,n776gat,II2035,n786gat,n551gat,
    II2040,n787gat,n775gat,II2044,n788gat,n657gat,II2049,n789gat,n35gat,n779gat,II2056,n125gat,n558gat,n559gat,n371gat,II2084,
    n365gat,II2088,n560gat,n364gat,II2094,n2876gat,n126gat,n663gat,II2109,n321gat,II2112,n226gat,n370gat,II2127,n317gat,II2130,
    n227gat,n369gat,II2145,n313gat,II2148,n228gat,n316gat,II2153,n229gat,n312gat,II2157,n230gat,n320gat,II2162,n231gat,n34gat,
    n221gat,II2169,n127gat,n133gat,II2174,n128gat,II2177,n129gat,II2181,n130gat,n665gat,n1601gat,n120gat,n2597gat,n2595gat,n2594gat,
    n2586gat,II2213,n2573gat,II2225,n2574gat,II2228,n2575gat,II2232,n2639gat,II2235,n2576gat,II2238,n2577gat,II2242,n2578gat,II2248,
    n2568gat,n2582gat,II2251,n2206gat,II2254,n2414gat,II2257,n2415gat,II2260,n2202gat,II2263,n2416gat,II2268,n2417gat,II2271,n2418gat,
    II2275,n2419gat,II2281,n2409gat,n2585gat,n2656gat,II2316,n2389gat,II2319,n2494gat,II2324,n3014gat,n2649gat,II2344,n2338gat,II2349,
    n2269gat,II2354,n2880gat,n2652gat,n2500gat,n2620gat,n2612gat,II2372,n2606gat,II2376,n2607gat,n2540gat,II2380,n2608gat,n2536gat,II2385,
    n2609gat,II2389,n2610gat,II2394,n2611gat,II2400,n2601gat,n2616gat,II2403,n2550gat,II2414,n2633gat,II2417,n2551gat,II2420,n2552gat,
    II2425,n2553gat,II2428,n2554gat,II2433,n2555gat,II2439,n2545gat,n2619gat,n2504gat,n2660gat,n2655gat,n1528gat,n2293gat,n1523gat,n2219gat,
    n1592gat,n1529gat,n2666gat,n1704gat,n2422gat,n3013gat,n2290gat,n2081gat,n2218gat,n2285gat,n2359gat,n2358gat,n1414gat,n1415gat,n566gat,n1480gat,
    n2292gat,n1301gat,n1416gat,n1150gat,n873gat,n2011gat,n2306gat,n1478gat,n1481gat,n875gat,n1410gat,n2357gat,n876gat,n1347gat,n1160gat,n1484gat,
    n1084gat,n983gat,n1482gat,n2363gat,n1157gat,n1483gat,n985gat,n1530gat,n2364gat,n1307gat,n1308gat,n1085gat,n1479gat,n2291gat,n1348gat,n1349gat,
    n2217gat,n1591gat,n2223gat,n1437gat,n1438gat,n1832gat,n1765gat,n1878gat,n1442gat,n1831gat,n1444gat,n1378gat,n2975gat,n1322gat,n2974gat,n1439gat,
    n1486gat,n1370gat,n1426gat,n1369gat,n2966gat,n1366gat,n1365gat,n1374gat,n2979gat,n2162gat,n2220gat,n1450gat,n1423gat,n1427gat,n1608gat,n2082gat,
    n1449gat,n1494gat,n1590gat,n1248gat,n2954gat,n1418gat,n1417gat,n1306gat,n2964gat,n1353gat,n1419gat,n1247gat,n2958gat,n1355gat,n1422gat,n1300gat,
    n2963gat,n1487gat,n1485gat,n1164gat,n2953gat,n1356gat,n1354gat,n1436gat,n1435gat,n1106gat,n2949gat,n1425gat,n1421gat,n1105gat,n2934gat,n1424gat,
    n1420gat,n1309gat,n2959gat,II2672,n2142gat,n1788gat,II2684,n2060gat,n1786gat,II2696,n2138gat,n1839gat,n1897gat,n1884gat,n1848gat,n1783gat,
    n1548gat,II2721,n1719gat,n2137gat,n1633gat,n2059gat,n1785gat,II2731,n1849gat,n1784gat,n1716gat,II2736,n1635gat,n2401gat,n1989gat,n2392gat,
    n1918gat,II2771,n2439gat,n1986gat,n1866gat,n1865gat,II2785,n2406gat,n2216gat,n2345gat,n1988gat,n1735gat,n1861gat,n1387gat,n1694gat,II2813,
    n1780gat,n2019gat,n1549gat,II2832,n1551gat,II2837,n2346gat,n2152gat,n2405gat,n2351gat,II2843,n2402gat,n2212gat,II2847,n2393gat,n1991gat,
    n1665gat,n1666gat,n1517gat,n1578gat,II2873,n1495gat,n1604gat,II2885,n2090gat,n1550gat,II2890,n1552gat,n1738gat,II2915,n1739gat,n1925gat,
    n1920gat,n1917gat,n1921gat,n2141gat,n1787gat,II2926,n1859gat,n1922gat,n1798gat,II2935,n1743gat,n1923gat,n1864gat,n1690gat,II2953,n2178gat,
    n1661gat,n1660gat,n1572gat,n1576gat,n2438gat,n2283gat,n1520gat,n1582gat,n1580gat,n1577gat,n1990gat,n2988gat,II2978,n2189gat,II2989,n2134gat,
    II3000,n2261gat,n2128gat,n2129gat,n1695gat,II3016,n2181gat,II3056,n1311gat,n1707gat,n1659gat,n2987gat,n1515gat,n1521gat,n1736gat,n1737gat,
    n1658gat,n1724gat,n1732gat,n1662gat,n1663gat,n1656gat,n1655gat,n1670gat,n1667gat,n1569gat,n1570gat,n1568gat,n1575gat,n1727gat,n1728gat,n1797gat,
    n1801gat,n1730gat,n1731gat,n1561gat,n1571gat,n1668gat,n1734gat,n1742gat,n1671gat,n1669gat,n1652gat,n1657gat,n1648gat,n1729gat,n1790gat,n1726gat,
    n2004gat,n1929gat,n1869gat,II3143,n2591gat,n1584gat,n1714gat,II3149,n1718gat,II3163,n1507gat,n1396gat,n1401gat,II3168,n1393gat,n1409gat,
    n1476gat,II3174,n1898gat,n1838gat,II3179,II3191,n1677gat,n2000gat,n1412gat,n2001gat,n1999gat,II3211,n2663gat,n3018gat,n2448gat,n2662gat,
    n2444gat,II3235,n2238gat,n3019gat,n1310gat,n199gat,n87gat,n195gat,n184gat,n204gat,II3273,n2168gat,n2452gat,n1691gat,II3287,n3020gat,
    II3290,n3021gat,II3293,n3022gat,n1699gat,II3297,n3023gat,II3300,n3024gat,II3303,n3025gat,II3306,n3026gat,II3309,n3027gat,II3312,
    n3028gat,II3315,n3029gat,II3318,n3030gat,n2260gat,n2257gat,n2188gat,n2187gat,n3004gat,II3336,n2039gat,II3339,n1774gat,II3342,n1315gat,
    n2097gat,n1855gat,n2014gat,II3387,n2194gat,II3390,n3032gat,n2256gat,II3394,n3033gat,n2251gat,n2184gat,n3003gat,II3401,n2192gat,n2133gat,
    n2131gat,n2185gat,n2049gat,n3001gat,II3412,n2057gat,n2253gat,n2252gat,n2248gat,n3006gat,n2264gat,II3429,n2265gat,n2492gat,n2329gat,II3436,
    n1709gat,n1845gat,n1891gat,n1963gat,n1886gat,n1968gat,n1958gat,n1629gat,n1895gat,n1631gat,n1711gat,n2990gat,n2200gat,n2078gat,n2437gat,n2195gat,
    II3457,n2556gat,n1956gat,II3461,n3038gat,n1954gat,II3465,n3039gat,n1888gat,n2048gat,n2994gat,II3472,n2539gat,n1969gat,n1893gat,n1892gat,
    n2993gat,II3483,n2436gat,n2056gat,n2998gat,II3491,n2387gat,II3494,n3043gat,n1960gat,n1887gat,n1961gat,n2996gat,II3504,n2330gat,n2199gat,
    n2147gat,II3509,n3045gat,n2332gat,II3513,n3046gat,n2259gat,n2328gat,n3008gat,II3520,n2498gat,n2151gat,n2193gat,n2209gat,n3005gat,II3530,
    n2396gat,n2052gat,n2058gat,n2997gat,II3539,n2198gat,n2349gat,n2215gat,n2281gat,n3009gat,II3549,n2197gat,n2146gat,n3002gat,II3558,n2196gat,
    II3587,n2124gat,n2115gat,II3610,n1882gat,II3621,n1974gat,n1955gat,n1970gat,n1896gat,n1973gat,n2558gat,n2559gat,II3635,II3646,n2643gat,
    n2333gat,n2564gat,n2352gat,n2642gat,n2636gat,n2637gat,II3660,n88gat,n84gat,n375gat,n110gat,II3677,n155gat,n253gat,n1702gat,n150gat,
    II3691,n151gat,n243gat,n233gat,n154gat,n800gat,n2874gat,II3703,n2917gat,n235gat,n2878gat,II3713,n2892gat,n372gat,n212gat,n329gat,
    II3736,n387gat,n334gat,n1700gat,n386gat,II3742,n330gat,n1430gat,n1490gat,n452gat,n2885gat,II3754,n2900gat,n333gat,n2883gat,II3765,
    n2929gat,II3777,n462gat,n325gat,n457gat,n2884gat,n461gat,n458gat,n2902gat,II3801,n2925gat,n144gat,n247gat,II3808,n326gat,n878gat,
    n2879gat,II3817,n2916gat,n382gat,II3831,n383gat,n134gat,n2875gat,II3841,n2899gat,n254gat,n252gat,n2877gat,n468gat,II3867,n469gat,
    n381gat,n2893gat,II3876,n2926gat,n241gat,n140gat,II3882,n255gat,n802gat,n2882gat,II3891,n2924gat,n146gat,II3904,n147gat,n380gat,
    n2881gat,II3914,n2923gat,n69gat,n68gat,n1885gat,II3923,n2710gat,n2707gat,n16gat,n295gat,n357gat,n11gat,n12gat,n1889gat,II3935,
    n2704gat,n2700gat,n2051gat,II3941,n2684gat,n2680gat,n1350gat,II3945,n2696gat,II3948,n2692gat,II3951,n2683gat,II3954,n2679gat,II3957,
    n2449gat,n1754gat,II3962,n2830gat,n2827gat,n2512gat,n1544gat,n1769gat,n1683gat,n1756gat,n2167gat,n2013gat,II4000,n1791gat,n2691gat,n2695gat,
    n1518gat,n2699gat,n2703gat,n2159gat,n2478gat,II4014,n2744gat,n2740gat,n2158gat,n2186gat,II4020,n2800gat,n2797gat,n2288gat,II4024,n1513gat,
    n2537gat,n2538gat,n2442gat,n2483gat,n1334gat,II4055,n1747gat,II4067,n1674gat,n1403gat,n1402gat,II4081,n1806gat,n1634gat,n1338gat,II4105,
    n1455gat,II4108,n1339gat,n1505gat,n2980gat,II4117,n2758gat,n2755gat,n1546gat,II4122,n2752gat,n2748gat,n2012gat,n2016gat,n2002gat,n2008gat,
    II4129,n2858gat,n2857gat,II4135,n2766gat,II4138,n2765gat,n1684gat,n1759gat,II4145,II4157,n1524gat,n1862gat,n1863gat,n1919gat,n1860gat,
    n1460gat,II4185,n1595gat,n1454gat,n1469gat,n1468gat,n1519gat,II4194,n1461gat,n1477gat,n2984gat,n1594gat,II4212,n1587gat,n1681gat,II4217,
    II4222,n1761gat,n2751gat,n2747gat,II4227,n1760gat,n2743gat,n2739gat,n1978gat,II4233,n1721gat,n2808gat,II4236,n2804gat,n517gat,n518gat,
    n417gat,n418gat,n413gat,n411gat,n412gat,n522gat,n406gat,n516gat,n407gat,n355gat,n290gat,n525gat,n527gat,n356gat,n416gat,n415gat,
    n528gat,n521gat,n358gat,n532gat,n639gat,n523gat,n1111gat,n635gat,n524gat,n414gat,n1112gat,n630gat,n741gat,n629gat,n633gat,n634gat,
    n926gat,n632gat,n670gat,n636gat,n1123gat,n1007gat,n1006gat,II4309,n2941gat,n2814gat,II4312,n2811gat,n1002gat,n2946gat,II4329,n2950gat,
    n2813gat,II4332,n2810gat,n888gat,n2933gat,II4349,n2935gat,n2818gat,II4352,n2816gat,n898gat,n2940gat,II4369,n2937gat,n2817gat,II4372,
    n2815gat,n1179gat,n2947gat,II4389,n2956gat,n2824gat,II4392,n2821gat,n897gat,n2939gat,II4409,n2938gat,n2823gat,II4412,n2820gat,n894gat,
    n2932gat,II4429,n2936gat,n2829gat,II4432,n2826gat,n1180gat,n2948gat,II4449,n2955gat,n2828gat,II4452,n2825gat,n671gat,n628gat,n631gat,
    n976gat,II4475,n2951gat,n2807gat,II4478,n2803gat,n2127gat,II4482,n2682gat,II4485,n2678gat,n2046gat,II4489,n2681gat,II4492,n2677gat,
    n1708gat,II4496,n2688gat,II4499,n2686gat,n455gat,n291gat,n2237gat,II4506,n2764gat,n2763gat,n1782gat,II4512,n2762gat,n2760gat,n2325gat,
    II4518,n2761gat,n2759gat,n2245gat,II4524,n2757gat,n2754gat,n2244gat,II4530,n2756gat,n2753gat,n2243gat,II4536,n2750gat,n2746gat,n2246gat,
    II4542,n2749gat,n2745gat,n2384gat,II4548,n2742gat,n2738gat,n2385gat,II4554,n2741gat,n2737gat,n1286gat,II4558,n2687gat,n2685gat,n1328gat,
    n1381gat,n1384gat,II4566,n2694gat,n2690gat,n1382gat,n1451gat,n1453gat,II4573,n2693gat,n2689gat,n927gat,n925gat,n1452gat,II4580,n2702gat,
    n2698gat,n923gat,n921gat,n1890gat,II4587,n2701gat,n2697gat,n850gat,n739gat,n1841gat,II4594,n2709gat,n2706gat,n922gat,n848gat,n2047gat,
    II4601,n2708gat,n2705gat,n924gat,n849gat,n2050gat,II4608,n2799gat,n2796gat,n1118gat,n1032gat,n2054gat,II4615,n2798gat,n2795gat,II4620,
    n1745gat,n2806gat,II4623,n2802gat,II4626,n1870gat,n1086gat,II4630,n2805gat,II4633,n2801gat,n67gat,n85gat,n71gat,n180gat,n1840gat,
    II4642,n2812gat,n2809gat,n76gat,n82gat,n14gat,n186gat,n1842gat,II4651,n2822gat,n2819gat,II4654,II4657,II4660,II4663,II4666,
    II4669,II4672,II4675,II4678,II4681,II4684,II4687,II4690,II4693,II4696,II4699,II4702,II4705,II4708,II4711,II4714,
    II4717,II4720,II4723,II4726,II4729,II4732,II4735,II4738,II4741,II4744,II4747,II4750,II4753,II4756,II4759,II4762,
    II4765,II4768,II4771,II4774,II4777,II4780,II4783,II4786,II4789,II4792,II4795,II4798,n648gat,n442gat,n1214gat,n1215gat,
    n1216gat,n1217gat,n745gat,n638gat,n423gat,n362gat,n749gat,n750gat,n751gat,n752gat,n259gat,n260gat,n261gat,n262gat,n1014gat,n1015gat,
    n1016gat,n1017gat,n476gat,n477gat,n478gat,n479gat,n44gat,n45gat,n46gat,n47gat,n168gat,n169gat,n170gat,n171gat,n907gat,n908gat,
    n909gat,n910gat,n344gat,n345gat,n346gat,n347gat,n56gat,n57gat,n58gat,n59gat,n768gat,n655gat,n963gat,n868gat,n962gat,n959gat,
    n945gat,n946gat,n947gat,n948gat,n647gat,n441gat,n967gat,n792gat,n1229gat,n1230gat,n1231gat,n1232gat,n443gat,n439gat,n966gat,n790gat,
    n444gat,n440gat,n1051gat,n1052gat,n1053gat,n1054gat,n934gat,n935gat,n936gat,n937gat,n710gat,n711gat,n712gat,n713gat,n729gat,n730gat,
    n731gat,n732gat,n494gat,n495gat,n496gat,n497gat,n505gat,n506gat,n507gat,n508gat,II1277,n767gat,n653gat,n867gat,n771gat,n964gat,
    n961gat,n804gat,n805gat,n806gat,n807gat,n587gat,n588gat,n589gat,n590gat,n447gat,n445gat,n687gat,n688gat,n689gat,n690gat,n568gat,
    n569gat,n570gat,n571gat,II1515,II1584,n1692gat,II1723,II1733,n2428gat,n769gat,n1076gat,n766gat,n1185gat,n1186gat,n1187gat,n1188gat,
    n645gat,n646gat,n1383gat,n1327gat,n651gat,n652gat,n765gat,n1202gat,n1203gat,n1204gat,n1205gat,n1270gat,n1271gat,n1272gat,n1273gat,n763gat,
    n1287gat,n1285gat,n793gat,n556gat,n795gat,n656gat,n794gat,n773gat,n965gat,n960gat,n780gat,n781gat,n782gat,n783gat,n555gat,n450gat,
    n654gat,n557gat,n874gat,n132gat,n649gat,n449gat,n791gat,n650gat,n774gat,n764gat,n222gat,n223gat,n224gat,n225gat,n121gat,n122gat,
    n123gat,n124gat,n2460gat,n2423gat,n2569gat,n2570gat,n2571gat,n2572gat,n2410gat,n2411gat,n2412gat,n2413gat,n2580gat,n2581gat,n2567gat,n2499gat,
    n299gat,n207gat,n2647gat,n2648gat,n2602gat,n2603gat,n2604gat,n2605gat,n2546gat,n2547gat,n2548gat,n2549gat,n2614gat,n2615gat,n2461gat,n2421gat,
    n2930gat,n1153gat,n1151gat,n982gat,n877gat,n2957gat,n1159gat,n1158gat,n1156gat,n1155gat,n1443gat,n1325gat,n1321gat,n1320gat,n1368gat,n1258gat,
    n1373gat,n1372gat,n2978gat,n1441gat,n1440gat,n1371gat,n1367gat,n2982gat,n1504gat,n1502gat,n1250gat,n1103gat,n1304gat,n1249gat,n1246gat,n1161gat,
    n1291gat,n1245gat,n2973gat,n1352gat,n1351gat,n1303gat,n1302gat,n1163gat,n1102gat,n1101gat,n996gat,n1104gat,n887gat,n1305gat,n1162gat,n2977gat,
    n1360gat,n1359gat,n1358gat,n1357gat,II2720,II2735,II2812,n1703gat,n1778gat,n1609gat,II2831,II2889,II2925,II2934,n1733gat,n1581gat,
    n2079gat,n2073gat,n1574gat,n1573gat,n2992gat,n1723gat,n1647gat,n1646gat,n2986gat,n1650gat,n1649gat,n1563gat,n2991gat,n1654gat,n1653gat,n1644gat,
    II3148,II3178,n2981gat,n1413gat,n1408gat,n1407gat,n2258gat,n2255gat,n2132gat,n2130gat,n3007gat,n2250gat,n2249gat,n1710gat,n1630gat,n1894gat,
    n1847gat,n1846gat,n2055gat,n1967gat,n1959gat,n1957gat,n2211gat,n2210gat,n2053gat,n1964gat,n2350gat,n2282gat,n2213gat,n2150gat,n2149gat,n2995gat,
    n1962gat,n2999gat,n1972gat,n1971gat,n3011gat,n2331gat,n3015gat,n2566gat,n2565gat,n141gat,n38gat,n37gat,n1074gat,n872gat,n234gat,n137gat,
    n378gat,n377gat,n250gat,n249gat,n248gat,n869gat,n453gat,n448gat,n251gat,n244gat,n974gat,n973gat,n870gat,n246gat,n245gat,n460gat,
    n459gat,n975gat,n972gat,n969gat,n145gat,n143gat,n971gat,n970gat,n968gat,n142gat,n40gat,n39gat,n772gat,n451gat,n446gat,n139gat,
    n136gat,n391gat,n390gat,n1083gat,n1077gat,n242gat,n240gat,n871gat,n797gat,n324gat,n238gat,n237gat,n1082gat,n796gat,n1599gat,II3999,
    n1586gat,n1755gat,II4023,n1470gat,n1400gat,n1399gat,n1398gat,II4144,n1467gat,n1466gat,n2985gat,n1686gat,n1533gat,n1532gat,n1531gat,II4216,
    n2931gat,n1100gat,n994gat,n989gat,n880gat,n2943gat,n1012gat,n905gat,n1003gat,n902gat,n1099gat,n998gat,n995gat,n980gat,n2960gat,n1175gat,
    n1174gat,n1001gat,n999gat,n2969gat,n1323gat,n1264gat,n981gat,n890gat,n889gat,n886gat,n892gat,n891gat,n2942gat,n904gat,n903gat,n1152gat,
    n1092gat,n997gat,n993gat,n900gat,n895gat,n1094gat,n1093gat,n988gat,n984gat,n2965gat,n1267gat,n1257gat,n1178gat,n1116gat,n2961gat,n1375gat,
    n1324gat,n1091gat,n1088gat,n992gat,n987gat,n899gat,n896gat,n2967gat,n1262gat,n1260gat,n1098gat,n1090gat,n986gat,n885gat,n901gat,n893gat,
    n1097gat,n1089gat,n1087gat,n991gat,n2968gat,n1326gat,n1261gat,n1177gat,n1115gat,n2944gat,n977gat,n2945gat,n1096gat,n1095gat,n990gat,n979gat,
    n2962gat,n1176gat,n1173gat,n1004gat,n1000gat,n1029gat,n1028gat,n1031gat,n1030gat,n1011gat,n1181gat,n1010gat,n1005gat,n1182gat,n73gat,n70gat,
    n77gat,n13gat,n1935gat,n197gat,n22gat,n93gat,n2239gat,n2433gat,n2427gat,n2583gat,n2650gat,n2617gat,n1598gat,n1154gat,n1411gat,n1498gat,
    n1607gat,n1428gat,n1794gat,n1796gat,n1792gat,n1406gat,n2664gat,n1926gat,n1916gat,n1994gat,n1924gat,n1758gat,n200gat,n196gat,n2018gat,n89gat,
    n1471gat,n1472gat,n1600gat,n1397gat,n2005gat,n1818gat,n1510gat,n1459gat,n1458gat,n1602gat,n520gat,n519gat,n410gat,n354gat,n408gat,n526gat,
    n531gat,n530gat,n359gat,n420gat,n801gat,n879gat,n1255gat,n1009gat,n409gat,n292gat,n419gat,n1243gat,n1171gat,n1244gat,n1265gat,n1254gat,
    n1008gat,n1253gat,n1266gat,n1200gat,n1172gat,n1251gat,n1259gat,n1212gat,n1263gat,n978gat,n1199gat,n1252gat,n1757gat,extra0,extra1,extra2,
    extra3,extra4,extra5,extra6,extra7,extra8,extra9,extra10,extra11;

  DFF_X1 DFF_0( .CK(CK), .Q(n673gat), .D(n2897gat) );
  DFF_X1 DFF_1( .CK(CK), .Q(n398gat), .D(n2782gat) );
  DFF_X1 DFF_2( .CK(CK), .Q(n402gat), .D(n2790gat) );
  DFF_X2 DFF_3( .CK(CK), .Q(n919gat), .D(n2670gat) );
  DFF_X2 DFF_4( .CK(CK), .Q(n846gat), .D(n2793gat) );
  DFF_X2 DFF_5( .CK(CK), .Q(n394gat), .D(n2782gat) );
  DFF_X1 DFF_6( .CK(CK), .Q(n703gat), .D(n2790gat) );
  DFF_X1 DFF_7( .CK(CK), .Q(n722gat), .D(n2670gat) );
  DFF_X1 DFF_8( .CK(CK), .Q(n726gat), .D(n2793gat) );
  DFF_X1 DFF_9( .CK(CK), .Q(n2510gat), .D(n748gat) );
  DFF_X1 DFF_10( .CK(CK), .Q(n271gat), .D(n2732gat) );
  DFF_X1 DFF_11( .CK(CK), .Q(n160gat), .D(n2776gat) );
  DFF_X1 DFF_12( .CK(CK), .Q(n337gat), .D(n2735gat) );
  DFF_X1 DFF_13( .CK(CK), .Q(n842gat), .D(n2673gat) );
  DFF_X1 DFF_14( .CK(CK), .Q(n341gat), .D(n2779gat) );
  DFF_X1 DFF_15( .CK(CK), .Q(n2522gat), .D(n43gat) );
  DFF_X1 DFF_16( .CK(CK), .Q(n2472gat), .D(n1620gat) );
  DFF_X1 DFF_17( .CK(CK), .Q(n2319gat), .D(n2470gat) );
  DFF_X1 DFF_18( .CK(CK), .Q(n1821gat), .D(n1827gat) );
  DFF_X1 DFF_19( .CK(CK), .Q(n1825gat), .D(n1827gat) );
  DFF_X1 DFF_20( .CK(CK), .Q(n2029gat), .D(n1816gat) );
  DFF_X1 DFF_21( .CK(CK), .Q(n1829gat), .D(n2027gat) );
  DFF_X1 DFF_22( .CK(CK), .Q(n283gat), .D(n2732gat) );
  DFF_X1 DFF_23( .CK(CK), .Q(n165gat), .D(n2776gat) );
  DFF_X1 DFF_24( .CK(CK), .Q(n279gat), .D(n2735gat) );
  DFF_X1 DFF_25( .CK(CK), .Q(n1026gat), .D(n2673gat) );
  DFF_X1 DFF_26( .CK(CK), .Q(n275gat), .D(n2779gat) );
  DFF_X1 DFF_27( .CK(CK), .Q(n2476gat), .D(n55gat) );
  DFF_X1 DFF_28( .CK(CK), .Q(n1068gat), .D(n2914gat) );
  DFF_X1 DFF_29( .CK(CK), .Q(n957gat), .D(n2928gat) );
  DFF_X1 DFF_30( .CK(CK), .Q(n861gat), .D(n2927gat) );
  DFF_X1 DFF_31( .CK(CK), .Q(n1294gat), .D(n2896gat) );
  DFF_X1 DFF_32( .CK(CK), .Q(n1241gat), .D(n2922gat) );
  DFF_X1 DFF_33( .CK(CK), .Q(n1298gat), .D(n2897gat) );
  DFF_X1 DFF_34( .CK(CK), .Q(n865gat), .D(n2894gat) );
  DFF_X1 DFF_35( .CK(CK), .Q(n1080gat), .D(n2921gat) );
  DFF_X1 DFF_36( .CK(CK), .Q(n1148gat), .D(n2895gat) );
  DFF_X1 DFF_37( .CK(CK), .Q(n2468gat), .D(n933gat) );
  DFF_X1 DFF_38( .CK(CK), .Q(n618gat), .D(n2790gat) );
  DFF_X1 DFF_39( .CK(CK), .Q(n491gat), .D(n2782gat) );
  DFF_X2 DFF_40( .CK(CK), .Q(n622gat), .D(n2793gat) );
  DFF_X2 DFF_41( .CK(CK), .Q(n626gat), .D(n2670gat) );
  DFF_X2 DFF_42( .CK(CK), .Q(n834gat), .D(n3064gat) );
  DFF_X1 DFF_43( .CK(CK), .Q(n707gat), .D(n3055gat) );
  DFF_X1 DFF_44( .CK(CK), .Q(n838gat), .D(n3063gat) );
  DFF_X1 DFF_45( .CK(CK), .Q(n830gat), .D(n3062gat) );
  DFF_X1 DFF_46( .CK(CK), .Q(n614gat), .D(n3056gat) );
  DFF_X1 DFF_47( .CK(CK), .Q(n2526gat), .D(n504gat) );
  DFF_X1 DFF_48( .CK(CK), .Q(n680gat), .D(n2913gat) );
  DFF_X1 DFF_49( .CK(CK), .Q(n816gat), .D(n2920gat) );
  DFF_X1 DFF_50( .CK(CK), .Q(n580gat), .D(n2905gat) );
  DFF_X1 DFF_51( .CK(CK), .Q(n824gat), .D(n3057gat) );
  DFF_X1 DFF_52( .CK(CK), .Q(n820gat), .D(n3059gat) );
  DFF_X1 DFF_53( .CK(CK), .Q(n883gat), .D(n3058gat) );
  DFF_X1 DFF_54( .CK(CK), .Q(n584gat), .D(n2898gat) );
  DFF_X1 DFF_55( .CK(CK), .Q(n684gat), .D(n3060gat) );
  DFF_X1 DFF_56( .CK(CK), .Q(n699gat), .D(n3061gat) );
  DFF_X1 DFF_57( .CK(CK), .Q(n2464gat), .D(n567gat) );
  DFF_X1 DFF_58( .CK(CK), .Q(n2399gat), .D(n3048gat) );
  DFF_X1 DFF_59( .CK(CK), .Q(n2343gat), .D(n3049gat) );
  DFF_X1 DFF_60( .CK(CK), .Q(n2203gat), .D(n3051gat) );
  DFF_X1 DFF_61( .CK(CK), .Q(n2562gat), .D(n3047gat) );
  DFF_X1 DFF_62( .CK(CK), .Q(n2207gat), .D(n3050gat) );
  DFF_X1 DFF_63( .CK(CK), .Q(n2626gat), .D(n3040gat) );
  DFF_X1 DFF_64( .CK(CK), .Q(n2490gat), .D(n3044gat) );
  DFF_X1 DFF_65( .CK(CK), .Q(n2622gat), .D(n3042gat) );
  DFF_X1 DFF_66( .CK(CK), .Q(n2630gat), .D(n3037gat) );
  DFF_X1 DFF_67( .CK(CK), .Q(n2543gat), .D(n3041gat) );
  DFF_X1 DFF_68( .CK(CK), .Q(n2102gat), .D(n1606gat) );
  DFF_X1 DFF_69( .CK(CK), .Q(n1880gat), .D(n3052gat) );
  DFF_X1 DFF_70( .CK(CK), .Q(n1763gat), .D(n1610gat) );
  DFF_X1 DFF_71( .CK(CK), .Q(n2155gat), .D(n1858gat) );
  DFF_X1 DFF_72( .CK(CK), .Q(n1035gat), .D(n2918gat) );
  DFF_X1 DFF_73( .CK(CK), .Q(n1121gat), .D(n2952gat) );
  DFF_X1 DFF_74( .CK(CK), .Q(n1072gat), .D(n2919gat) );
  DFF_X1 DFF_75( .CK(CK), .Q(n1282gat), .D(n2910gat) );
  DFF_X1 DFF_76( .CK(CK), .Q(n1226gat), .D(n2907gat) );
  DFF_X1 DFF_77( .CK(CK), .Q(n931gat), .D(n2911gat) );
  DFF_X1 DFF_78( .CK(CK), .Q(n1135gat), .D(n2912gat) );
  DFF_X1 DFF_79( .CK(CK), .Q(n1045gat), .D(n2909gat) );
  DFF_X1 DFF_80( .CK(CK), .Q(n1197gat), .D(n2908gat) );
  DFF_X1 DFF_81( .CK(CK), .Q(n2518gat), .D(n2971gat) );
  DFF_X1 DFF_82( .CK(CK), .Q(n667gat), .D(n2904gat) );
  DFF_X1 DFF_83( .CK(CK), .Q(n659gat), .D(n2891gat) );
  DFF_X1 DFF_84( .CK(CK), .Q(n553gat), .D(n2903gat) );
  DFF_X1 DFF_85( .CK(CK), .Q(n777gat), .D(n2915gat) );
  DFF_X1 DFF_86( .CK(CK), .Q(n561gat), .D(n2901gat) );
  DFF_X1 DFF_87( .CK(CK), .Q(n366gat), .D(n2890gat) );
  DFF_X1 DFF_88( .CK(CK), .Q(n322gat), .D(n2888gat) );
  DFF_X1 DFF_89( .CK(CK), .Q(n318gat), .D(n2887gat) );
  DFF_X1 DFF_90( .CK(CK), .Q(n314gat), .D(n2886gat) );
  DFF_X1 DFF_91( .CK(CK), .Q(n2599gat), .D(n3010gat) );
  DFF_X1 DFF_92( .CK(CK), .Q(n2588gat), .D(n3016gat) );
  DFF_X1 DFF_93( .CK(CK), .Q(n2640gat), .D(n3054gat) );
  DFF_X1 DFF_94( .CK(CK), .Q(n2658gat), .D(n2579gat) );
  DFF_X1 DFF_95( .CK(CK), .Q(n2495gat), .D(n3036gat) );
  DFF_X1 DFF_96( .CK(CK), .Q(n2390gat), .D(n3034gat) );
  DFF_X1 DFF_97( .CK(CK), .Q(n2270gat), .D(n3031gat) );
  DFF_X1 DFF_98( .CK(CK), .Q(n2339gat), .D(n3035gat) );
  DFF_X1 DFF_99( .CK(CK), .Q(n2502gat), .D(n2646gat) );
  DFF_X1 DFF_100( .CK(CK), .Q(n2634gat), .D(n3053gat) );
  DFF_X1 DFF_101( .CK(CK), .Q(n2506gat), .D(n2613gat) );
  DFF_X1 DFF_102( .CK(CK), .Q(n1834gat), .D(n1625gat) );
  DFF_X1 DFF_103( .CK(CK), .Q(n1767gat), .D(n1626gat) );
  DFF_X1 DFF_104( .CK(CK), .Q(n2084gat), .D(n1603gat) );
  DFF_X1 DFF_105( .CK(CK), .Q(n2143gat), .D(n2541gat) );
  DFF_X1 DFF_106( .CK(CK), .Q(n2061gat), .D(n2557gat) );
  DFF_X1 DFF_107( .CK(CK), .Q(n2139gat), .D(n2487gat) );
  DFF_X1 DFF_108( .CK(CK), .Q(n1899gat), .D(n2532gat) );
  DFF_X1 DFF_109( .CK(CK), .Q(n1850gat), .D(n2628gat) );
  DFF_X1 DFF_110( .CK(CK), .Q(n2403gat), .D(n2397gat) );
  DFF_X1 DFF_111( .CK(CK), .Q(n2394gat), .D(n2341gat) );
  DFF_X1 DFF_112( .CK(CK), .Q(n2440gat), .D(n2560gat) );
  DFF_X1 DFF_113( .CK(CK), .Q(n2407gat), .D(n2205gat) );
  DFF_X1 DFF_114( .CK(CK), .Q(n2347gat), .D(n2201gat) );
  DFF_X1 DFF_115( .CK(CK), .Q(n1389gat), .D(n1793gat) );
  DFF_X1 DFF_116( .CK(CK), .Q(n2021gat), .D(n1781gat) );
  DFF_X1 DFF_117( .CK(CK), .Q(n1394gat), .D(n1516gat) );
  DFF_X1 DFF_118( .CK(CK), .Q(n1496gat), .D(n1392gat) );
  DFF_X1 DFF_119( .CK(CK), .Q(n2091gat), .D(n1685gat) );
  DFF_X1 DFF_120( .CK(CK), .Q(n1332gat), .D(n1565gat) );
  DFF_X1 DFF_121( .CK(CK), .Q(n1740gat), .D(n1330gat) );
  DFF_X1 DFF_122( .CK(CK), .Q(n2179gat), .D(n1945gat) );
  DFF_X1 DFF_123( .CK(CK), .Q(n2190gat), .D(n2268gat) );
  DFF_X1 DFF_124( .CK(CK), .Q(n2135gat), .D(n2337gat) );
  DFF_X1 DFF_125( .CK(CK), .Q(n2262gat), .D(n2388gat) );
  DFF_X1 DFF_126( .CK(CK), .Q(n2182gat), .D(n1836gat) );
  DFF_X1 DFF_127( .CK(CK), .Q(n1433gat), .D(n2983gat) );
  DFF_X1 DFF_128( .CK(CK), .Q(n1316gat), .D(n1431gat) );
  DFF_X1 DFF_129( .CK(CK), .Q(n1363gat), .D(n1314gat) );
  DFF_X1 DFF_130( .CK(CK), .Q(n1312gat), .D(n1361gat) );
  DFF_X1 DFF_131( .CK(CK), .Q(n1775gat), .D(n1696gat) );
  DFF_X1 DFF_132( .CK(CK), .Q(n1871gat), .D(n2009gat) );
  DFF_X1 DFF_133( .CK(CK), .Q(n2592gat), .D(n1773gat) );
  DFF_X1 DFF_134( .CK(CK), .Q(n1508gat), .D(n1636gat) );
  DFF_X1 DFF_135( .CK(CK), .Q(n1678gat), .D(n1712gat) );
  DFF_X1 DFF_136( .CK(CK), .Q(n2309gat), .D(n3000gat) );
  DFF_X1 DFF_137( .CK(CK), .Q(n2450gat), .D(n2307gat) );
  DFF_X1 DFF_138( .CK(CK), .Q(n2446gat), .D(n2661gat) );
  DFF_X1 DFF_139( .CK(CK), .Q(n2095gat), .D(n827gat) );
  DFF_X1 DFF_140( .CK(CK), .Q(n2176gat), .D(n2093gat) );
  DFF_X1 DFF_141( .CK(CK), .Q(n2169gat), .D(n2174gat) );
  DFF_X1 DFF_142( .CK(CK), .Q(n2454gat), .D(n2163gat) );
  DFF_X1 DFF_143( .CK(CK), .Q(n2040gat), .D(n1777gat) );
  DFF_X1 DFF_144( .CK(CK), .Q(n2044gat), .D(n2015gat) );
  DFF_X1 DFF_145( .CK(CK), .Q(n2037gat), .D(n2042gat) );
  DFF_X1 DFF_146( .CK(CK), .Q(n2025gat), .D(n2017gat) );
  DFF_X1 DFF_147( .CK(CK), .Q(n2099gat), .D(n2023gat) );
  DFF_X1 DFF_148( .CK(CK), .Q(n2266gat), .D(n2493gat) );
  DFF_X1 DFF_149( .CK(CK), .Q(n2033gat), .D(n2035gat) );
  DFF_X1 DFF_150( .CK(CK), .Q(n2110gat), .D(n2031gat) );
  DFF_X1 DFF_151( .CK(CK), .Q(n2125gat), .D(n2108gat) );
  DFF_X1 DFF_152( .CK(CK), .Q(n2121gat), .D(n2123gat) );
  DFF_X1 DFF_153( .CK(CK), .Q(n2117gat), .D(n2119gat) );
  DFF_X1 DFF_154( .CK(CK), .Q(n1975gat), .D(n2632gat) );
  DFF_X1 DFF_155( .CK(CK), .Q(n2644gat), .D(n2638gat) );
  DFF_X1 DFF_156( .CK(CK), .Q(n156gat), .D(n612gat) );
  DFF_X1 DFF_157( .CK(CK), .Q(n152gat), .D(n705gat) );
  DFF_X1 DFF_158( .CK(CK), .Q(n331gat), .D(n822gat) );
  DFF_X1 DFF_159( .CK(CK), .Q(n388gat), .D(n881gat) );
  DFF_X1 DFF_160( .CK(CK), .Q(n463gat), .D(n818gat) );
  DFF_X1 DFF_161( .CK(CK), .Q(n327gat), .D(n682gat) );
  DFF_X1 DFF_162( .CK(CK), .Q(n384gat), .D(n697gat) );
  DFF_X1 DFF_163( .CK(CK), .Q(n256gat), .D(n836gat) );
  DFF_X1 DFF_164( .CK(CK), .Q(n470gat), .D(n828gat) );
  DFF_X1 DFF_165( .CK(CK), .Q(n148gat), .D(n832gat) );
  DFF_X1 DFF_166( .CK(CK), .Q(n2458gat), .D(n2590gat) );
  DFF_X2 DFF_167( .CK(CK), .Q(n2514gat), .D(n2456gat) );
  DFF_X2 DFF_168( .CK(CK), .Q(n1771gat), .D(n1613gat) );
  DFF_X2 DFF_169( .CK(CK), .Q(n1336gat), .D(n1391gat) );
  DFF_X2 DFF_170( .CK(CK), .Q(n1748gat), .D(n1927gat) );
  DFF_X1 DFF_171( .CK(CK), .Q(n1675gat), .D(n1713gat) );
  DFF_X1 DFF_172( .CK(CK), .Q(n1807gat), .D(n1717gat) );
  DFF_X1 DFF_173( .CK(CK), .Q(n1340gat), .D(n1567gat) );
  DFF_X1 DFF_174( .CK(CK), .Q(n1456gat), .D(n1564gat) );
  DFF_X1 DFF_175( .CK(CK), .Q(n1525gat), .D(n1632gat) );
  DFF_X1 DFF_176( .CK(CK), .Q(n1462gat), .D(n1915gat) );
  DFF_X1 DFF_177( .CK(CK), .Q(n1596gat), .D(n1800gat) );
  DFF_X1 DFF_178( .CK(CK), .Q(n1588gat), .D(n1593gat) );
  INV_X1 NOT_0( .ZN(II1), .A(n3088gat) );
  INV_X1 NOT_1( .ZN(n2717gat), .A(II1) );
  INV_X1 NOT_2( .ZN(n2715gat), .A(n2717gat) );
  INV_X1 NOT_3( .ZN(II5), .A(n3087gat) );
  INV_X1 NOT_4( .ZN(n2725gat), .A(II5) );
  INV_X1 NOT_5( .ZN(n2723gat), .A(n2725gat) );
  INV_X1 NOT_6( .ZN(n296gat), .A(n421gat) );
  INV_X1 NOT_7( .ZN(II11), .A(n3093gat) );
  INV_X1 NOT_8( .ZN(n2768gat), .A(II11) );
  INV_X1 NOT_9( .ZN(II14), .A(n2768gat) );
  INV_X1 NOT_10( .ZN(n2767gat), .A(II14) );
  INV_X1 NOT_11( .ZN(n373gat), .A(n2767gat) );
  INV_X1 NOT_12( .ZN(II18), .A(n3072gat) );
  INV_X1 NOT_13( .ZN(n2671gat), .A(II18) );
  INV_X1 NOT_14( .ZN(n2669gat), .A(n2671gat) );
  INV_X1 NOT_15( .ZN(II23), .A(n3081gat) );
  INV_X1 NOT_16( .ZN(n2845gat), .A(II23) );
  INV_X1 NOT_17( .ZN(n2844gat), .A(n2845gat) );
  INV_X1 NOT_18( .ZN(II27), .A(n3095gat) );
  INV_X2 NOT_19( .ZN(n2668gat), .A(II27) );
  INV_X1 NOT_20( .ZN(II30), .A(n2668gat) );
  INV_X1 NOT_21( .ZN(n2667gat), .A(II30) );
  INV_X1 NOT_22( .ZN(n856gat), .A(n2667gat) );
  INV_X1 NOT_23( .ZN(II44), .A(n673gat) );
  INV_X1 NOT_24( .ZN(n672gat), .A(II44) );
  INV_X1 NOT_25( .ZN(II47), .A(n3069gat) );
  INV_X1 NOT_26( .ZN(n2783gat), .A(II47) );
  INV_X1 NOT_27( .ZN(II50), .A(n2783gat) );
  INV_X1 NOT_28( .ZN(n2782gat), .A(II50) );
  INV_X1 NOT_29( .ZN(n396gat), .A(n398gat) );
  INV_X1 NOT_30( .ZN(II62), .A(n3070gat) );
  INV_X1 NOT_31( .ZN(n2791gat), .A(II62) );
  INV_X1 NOT_32( .ZN(II65), .A(n2791gat) );
  INV_X1 NOT_33( .ZN(n2790gat), .A(II65) );
  INV_X1 NOT_34( .ZN(II76), .A(n402gat) );
  INV_X1 NOT_35( .ZN(n401gat), .A(II76) );
  INV_X1 NOT_36( .ZN(n1645gat), .A(n1499gat) );
  INV_X1 NOT_37( .ZN(II81), .A(n2671gat) );
  INV_X1 NOT_38( .ZN(n2670gat), .A(II81) );
  INV_X1 NOT_39( .ZN(II92), .A(n919gat) );
  INV_X1 NOT_40( .ZN(n918gat), .A(II92) );
  INV_X1 NOT_41( .ZN(n1553gat), .A(n1616gat) );
  INV_X1 NOT_42( .ZN(II97), .A(n3071gat) );
  INV_X1 NOT_43( .ZN(n2794gat), .A(II97) );
  INV_X1 NOT_44( .ZN(II100), .A(n2794gat) );
  INV_X1 NOT_45( .ZN(n2793gat), .A(II100) );
  INV_X1 NOT_46( .ZN(II111), .A(n846gat) );
  INV_X1 NOT_47( .ZN(n845gat), .A(II111) );
  INV_X1 NOT_48( .ZN(n1559gat), .A(n1614gat) );
  INV_X1 NOT_49( .ZN(n1643gat), .A(n1641gat) );
  INV_X1 NOT_50( .ZN(n1651gat), .A(n1642gat) );
  INV_X1 NOT_51( .ZN(n1562gat), .A(n1556gat) );
  INV_X1 NOT_52( .ZN(n1560gat), .A(n1557gat) );
  INV_X1 NOT_53( .ZN(n1640gat), .A(n1639gat) );
  INV_X1 NOT_54( .ZN(n1566gat), .A(n1605gat) );
  INV_X1 NOT_55( .ZN(n1554gat), .A(n1555gat) );
  INV_X1 NOT_56( .ZN(n1722gat), .A(n1558gat) );
  INV_X1 NOT_57( .ZN(n392gat), .A(n394gat) );
  INV_X1 NOT_58( .ZN(II149), .A(n703gat) );
  INV_X1 NOT_59( .ZN(n702gat), .A(II149) );
  INV_X1 NOT_60( .ZN(n1319gat), .A(n1256gat) );
  INV_X1 NOT_61( .ZN(n720gat), .A(n722gat) );
  INV_X1 NOT_62( .ZN(II171), .A(n726gat) );
  INV_X1 NOT_63( .ZN(n725gat), .A(II171) );
  INV_X1 NOT_64( .ZN(n1447gat), .A(n1117gat) );
  INV_X1 NOT_65( .ZN(n1627gat), .A(n1618gat) );
  INV_X1 NOT_66( .ZN(II178), .A(n722gat) );
  INV_X1 NOT_67( .ZN(n721gat), .A(II178) );
  INV_X1 NOT_68( .ZN(n1380gat), .A(n1114gat) );
  INV_X1 NOT_69( .ZN(n1628gat), .A(n1621gat) );
  INV_X1 NOT_70( .ZN(n701gat), .A(n703gat) );
  INV_X1 NOT_71( .ZN(n1446gat), .A(n1318gat) );
  INV_X1 NOT_72( .ZN(n1705gat), .A(n1619gat) );
  INV_X8 NOT_73( .ZN(n1706gat), .A(n1622gat) );
  INV_X8 NOT_74( .ZN(II192), .A(n3083gat) );
  INV_X1 NOT_75( .ZN(n2856gat), .A(II192) );
  INV_X1 NOT_76( .ZN(n2854gat), .A(n2856gat) );
  INV_X1 NOT_77( .ZN(II196), .A(n2854gat) );
  INV_X1 NOT_78( .ZN(n1218gat), .A(II196) );
  INV_X1 NOT_79( .ZN(II199), .A(n3085gat) );
  INV_X1 NOT_80( .ZN(n2861gat), .A(II199) );
  INV_X1 NOT_81( .ZN(n2859gat), .A(n2861gat) );
  INV_X1 NOT_82( .ZN(II203), .A(n2859gat) );
  INV_X1 NOT_83( .ZN(n1219gat), .A(II203) );
  INV_X1 NOT_84( .ZN(II206), .A(n3084gat) );
  INV_X1 NOT_85( .ZN(n2864gat), .A(II206) );
  INV_X1 NOT_86( .ZN(n2862gat), .A(n2864gat) );
  INV_X1 NOT_87( .ZN(II210), .A(n2862gat) );
  INV_X1 NOT_88( .ZN(n1220gat), .A(II210) );
  INV_X1 NOT_89( .ZN(II214), .A(n2861gat) );
  INV_X1 NOT_90( .ZN(n2860gat), .A(II214) );
  INV_X1 NOT_91( .ZN(II217), .A(n2860gat) );
  INV_X1 NOT_92( .ZN(n1221gat), .A(II217) );
  INV_X1 NOT_93( .ZN(II220), .A(n2864gat) );
  INV_X1 NOT_94( .ZN(n2863gat), .A(II220) );
  INV_X1 NOT_95( .ZN(II223), .A(n2863gat) );
  INV_X16 NOT_96( .ZN(n1222gat), .A(II223) );
  INV_X16 NOT_97( .ZN(II227), .A(n2856gat) );
  INV_X1 NOT_98( .ZN(n2855gat), .A(II227) );
  INV_X1 NOT_99( .ZN(II230), .A(n2855gat) );
  INV_X1 NOT_100( .ZN(n1223gat), .A(II230) );
  INV_X1 NOT_101( .ZN(n640gat), .A(n1213gat) );
  INV_X1 NOT_102( .ZN(II237), .A(n640gat) );
  INV_X1 NOT_103( .ZN(n753gat), .A(II237) );
  INV_X1 NOT_104( .ZN(II240), .A(n2717gat) );
  INV_X1 NOT_105( .ZN(n2716gat), .A(II240) );
  INV_X1 NOT_106( .ZN(II243), .A(n3089gat) );
  INV_X1 NOT_107( .ZN(n2869gat), .A(II243) );
  INV_X1 NOT_108( .ZN(n2867gat), .A(n2869gat) );
  INV_X1 NOT_109( .ZN(II248), .A(n2869gat) );
  INV_X1 NOT_110( .ZN(n2868gat), .A(II248) );
  INV_X1 NOT_111( .ZN(II253), .A(n2906gat) );
  INV_X1 NOT_112( .ZN(n754gat), .A(II253) );
  INV_X1 NOT_113( .ZN(II256), .A(n2725gat) );
  INV_X1 NOT_114( .ZN(n2724gat), .A(II256) );
  INV_X1 NOT_115( .ZN(II259), .A(n3086gat) );
  INV_X1 NOT_116( .ZN(n2728gat), .A(II259) );
  INV_X1 NOT_117( .ZN(n2726gat), .A(n2728gat) );
  INV_X1 NOT_118( .ZN(II264), .A(n2728gat) );
  INV_X1 NOT_119( .ZN(n2727gat), .A(II264) );
  INV_X1 NOT_120( .ZN(n422gat), .A(n2889gat) );
  INV_X1 NOT_121( .ZN(II270), .A(n422gat) );
  INV_X1 NOT_122( .ZN(n755gat), .A(II270) );
  INV_X1 NOT_123( .ZN(n747gat), .A(n2906gat) );
  INV_X1 NOT_124( .ZN(II275), .A(n747gat) );
  INV_X1 NOT_125( .ZN(n756gat), .A(II275) );
  INV_X1 NOT_126( .ZN(II278), .A(n2889gat) );
  INV_X1 NOT_127( .ZN(n757gat), .A(II278) );
  INV_X1 NOT_128( .ZN(II282), .A(n1213gat) );
  INV_X1 NOT_129( .ZN(n758gat), .A(II282) );
  INV_X1 NOT_130( .ZN(n2508gat), .A(n2510gat) );
  INV_X1 NOT_131( .ZN(II297), .A(n3065gat) );
  INV_X1 NOT_132( .ZN(n2733gat), .A(II297) );
  INV_X1 NOT_133( .ZN(II300), .A(n2733gat) );
  INV_X1 NOT_134( .ZN(n2732gat), .A(II300) );
  INV_X1 NOT_135( .ZN(II311), .A(n271gat) );
  INV_X1 NOT_136( .ZN(n270gat), .A(II311) );
  INV_X1 NOT_137( .ZN(II314), .A(n270gat) );
  INV_X1 NOT_138( .ZN(n263gat), .A(II314) );
  INV_X1 NOT_139( .ZN(II317), .A(n3067gat) );
  INV_X1 NOT_140( .ZN(n2777gat), .A(II317) );
  INV_X1 NOT_141( .ZN(II320), .A(n2777gat) );
  INV_X1 NOT_142( .ZN(n2776gat), .A(II320) );
  INV_X1 NOT_143( .ZN(II331), .A(n160gat) );
  INV_X1 NOT_144( .ZN(n159gat), .A(II331) );
  INV_X1 NOT_145( .ZN(II334), .A(n159gat) );
  INV_X1 NOT_146( .ZN(n264gat), .A(II334) );
  INV_X1 NOT_147( .ZN(II337), .A(n3066gat) );
  INV_X1 NOT_148( .ZN(n2736gat), .A(II337) );
  INV_X1 NOT_149( .ZN(II340), .A(n2736gat) );
  INV_X1 NOT_150( .ZN(n2735gat), .A(II340) );
  INV_X1 NOT_151( .ZN(II351), .A(n337gat) );
  INV_X1 NOT_152( .ZN(n336gat), .A(II351) );
  INV_X1 NOT_153( .ZN(II354), .A(n336gat) );
  INV_X1 NOT_154( .ZN(n265gat), .A(II354) );
  INV_X1 NOT_155( .ZN(n158gat), .A(n160gat) );
  INV_X1 NOT_156( .ZN(II359), .A(n158gat) );
  INV_X1 NOT_157( .ZN(n266gat), .A(II359) );
  INV_X1 NOT_158( .ZN(n335gat), .A(n337gat) );
  INV_X1 NOT_159( .ZN(II363), .A(n335gat) );
  INV_X1 NOT_160( .ZN(n267gat), .A(II363) );
  INV_X1 NOT_161( .ZN(n269gat), .A(n271gat) );
  INV_X1 NOT_162( .ZN(II368), .A(n269gat) );
  INV_X1 NOT_163( .ZN(n268gat), .A(II368) );
  INV_X1 NOT_164( .ZN(n41gat), .A(n258gat) );
  INV_X1 NOT_165( .ZN(II375), .A(n41gat) );
  INV_X1 NOT_166( .ZN(n48gat), .A(II375) );
  INV_X1 NOT_167( .ZN(II378), .A(n725gat) );
  INV_X1 NOT_168( .ZN(n1018gat), .A(II378) );
  INV_X1 NOT_169( .ZN(II381), .A(n3073gat) );
  INV_X2 NOT_170( .ZN(n2674gat), .A(II381) );
  INV_X2 NOT_171( .ZN(II384), .A(n2674gat) );
  INV_X2 NOT_172( .ZN(n2673gat), .A(II384) );
  INV_X1 NOT_173( .ZN(II395), .A(n842gat) );
  INV_X1 NOT_174( .ZN(n841gat), .A(II395) );
  INV_X1 NOT_175( .ZN(II398), .A(n841gat) );
  INV_X1 NOT_176( .ZN(n1019gat), .A(II398) );
  INV_X1 NOT_177( .ZN(II401), .A(n721gat) );
  INV_X1 NOT_178( .ZN(n1020gat), .A(II401) );
  INV_X1 NOT_179( .ZN(n840gat), .A(n842gat) );
  INV_X1 NOT_180( .ZN(II406), .A(n840gat) );
  INV_X1 NOT_181( .ZN(n1021gat), .A(II406) );
  INV_X1 NOT_182( .ZN(II409), .A(n720gat) );
  INV_X1 NOT_183( .ZN(n1022gat), .A(II409) );
  INV_X1 NOT_184( .ZN(n724gat), .A(n726gat) );
  INV_X1 NOT_185( .ZN(II414), .A(n724gat) );
  INV_X1 NOT_186( .ZN(n1023gat), .A(II414) );
  INV_X1 NOT_187( .ZN(II420), .A(n1013gat) );
  INV_X1 NOT_188( .ZN(n49gat), .A(II420) );
  INV_X1 NOT_189( .ZN(II423), .A(n3068gat) );
  INV_X1 NOT_190( .ZN(n2780gat), .A(II423) );
  INV_X1 NOT_191( .ZN(II426), .A(n2780gat) );
  INV_X1 NOT_192( .ZN(n2779gat), .A(II426) );
  INV_X1 NOT_193( .ZN(II437), .A(n341gat) );
  INV_X1 NOT_194( .ZN(n340gat), .A(II437) );
  INV_X1 NOT_195( .ZN(II440), .A(n340gat) );
  INV_X1 NOT_196( .ZN(n480gat), .A(II440) );
  INV_X1 NOT_197( .ZN(II443), .A(n702gat) );
  INV_X1 NOT_198( .ZN(n481gat), .A(II443) );
  INV_X1 NOT_199( .ZN(II446), .A(n394gat) );
  INV_X1 NOT_200( .ZN(n393gat), .A(II446) );
  INV_X1 NOT_201( .ZN(II449), .A(n393gat) );
  INV_X1 NOT_202( .ZN(n482gat), .A(II449) );
  INV_X1 NOT_203( .ZN(II453), .A(n701gat) );
  INV_X1 NOT_204( .ZN(n483gat), .A(II453) );
  INV_X1 NOT_205( .ZN(II456), .A(n392gat) );
  INV_X1 NOT_206( .ZN(n484gat), .A(II456) );
  INV_X1 NOT_207( .ZN(n339gat), .A(n341gat) );
  INV_X1 NOT_208( .ZN(II461), .A(n339gat) );
  INV_X1 NOT_209( .ZN(n485gat), .A(II461) );
  INV_X1 NOT_210( .ZN(n42gat), .A(n475gat) );
  INV_X1 NOT_211( .ZN(II468), .A(n42gat) );
  INV_X1 NOT_212( .ZN(n50gat), .A(II468) );
  INV_X1 NOT_213( .ZN(n162gat), .A(n1013gat) );
  INV_X1 NOT_214( .ZN(II473), .A(n162gat) );
  INV_X1 NOT_215( .ZN(n51gat), .A(II473) );
  INV_X1 NOT_216( .ZN(II476), .A(n475gat) );
  INV_X1 NOT_217( .ZN(n52gat), .A(II476) );
  INV_X1 NOT_218( .ZN(II480), .A(n258gat) );
  INV_X1 NOT_219( .ZN(n53gat), .A(II480) );
  INV_X1 NOT_220( .ZN(n2520gat), .A(n2522gat) );
  INV_X1 NOT_221( .ZN(n1448gat), .A(n1376gat) );
  INV_X1 NOT_222( .ZN(n1701gat), .A(n1617gat) );
  INV_X8 NOT_223( .ZN(n1379gat), .A(n1377gat) );
  INV_X8 NOT_224( .ZN(n1615gat), .A(n1624gat) );
  INV_X1 NOT_225( .ZN(n1500gat), .A(n1113gat) );
  INV_X1 NOT_226( .ZN(n1503gat), .A(n1501gat) );
  INV_X1 NOT_227( .ZN(n1779gat), .A(n1623gat) );
  INV_X1 NOT_228( .ZN(II509), .A(n3099gat) );
  INV_X1 NOT_229( .ZN(n2730gat), .A(II509) );
  INV_X1 NOT_230( .ZN(II512), .A(n2730gat) );
  INV_X1 NOT_231( .ZN(n2729gat), .A(II512) );
  INV_X1 NOT_232( .ZN(n2470gat), .A(n2472gat) );
  INV_X1 NOT_233( .ZN(n2317gat), .A(n2319gat) );
  INV_X1 NOT_234( .ZN(n1819gat), .A(n1821gat) );
  INV_X1 NOT_235( .ZN(n1823gat), .A(n1825gat) );
  INV_X1 NOT_236( .ZN(n1816gat), .A(n1817gat) );
  INV_X1 NOT_237( .ZN(n2027gat), .A(n2029gat) );
  INV_X1 NOT_238( .ZN(II572), .A(n1829gat) );
  INV_X1 NOT_239( .ZN(n1828gat), .A(II572) );
  INV_X1 NOT_240( .ZN(II576), .A(n3100gat) );
  INV_X1 NOT_241( .ZN(n2851gat), .A(II576) );
  INV_X1 NOT_242( .ZN(II579), .A(n2851gat) );
  INV_X1 NOT_243( .ZN(n2850gat), .A(II579) );
  INV_X1 NOT_244( .ZN(II583), .A(n2786gat) );
  INV_X1 NOT_245( .ZN(n2785gat), .A(II583) );
  INV_X1 NOT_246( .ZN(n92gat), .A(n2785gat) );
  INV_X1 NOT_247( .ZN(n637gat), .A(n529gat) );
  INV_X1 NOT_248( .ZN(n293gat), .A(n361gat) );
  INV_X1 NOT_249( .ZN(II591), .A(n3094gat) );
  INV_X1 NOT_250( .ZN(n2722gat), .A(II591) );
  INV_X1 NOT_251( .ZN(II594), .A(n2722gat) );
  INV_X1 NOT_252( .ZN(n2721gat), .A(II594) );
  INV_X1 NOT_253( .ZN(n297gat), .A(n2721gat) );
  INV_X1 NOT_254( .ZN(II606), .A(n283gat) );
  INV_X1 NOT_255( .ZN(n282gat), .A(II606) );
  INV_X1 NOT_256( .ZN(II609), .A(n282gat) );
  INV_X1 NOT_257( .ZN(n172gat), .A(II609) );
  INV_X1 NOT_258( .ZN(II620), .A(n165gat) );
  INV_X1 NOT_259( .ZN(n164gat), .A(II620) );
  INV_X1 NOT_260( .ZN(II623), .A(n164gat) );
  INV_X1 NOT_261( .ZN(n173gat), .A(II623) );
  INV_X1 NOT_262( .ZN(II634), .A(n279gat) );
  INV_X1 NOT_263( .ZN(n278gat), .A(II634) );
  INV_X1 NOT_264( .ZN(II637), .A(n278gat) );
  INV_X1 NOT_265( .ZN(n174gat), .A(II637) );
  INV_X1 NOT_266( .ZN(n163gat), .A(n165gat) );
  INV_X1 NOT_267( .ZN(II642), .A(n163gat) );
  INV_X1 NOT_268( .ZN(n175gat), .A(II642) );
  INV_X1 NOT_269( .ZN(n277gat), .A(n279gat) );
  INV_X1 NOT_270( .ZN(II646), .A(n277gat) );
  INV_X1 NOT_271( .ZN(n176gat), .A(II646) );
  INV_X1 NOT_272( .ZN(n281gat), .A(n283gat) );
  INV_X1 NOT_273( .ZN(II651), .A(n281gat) );
  INV_X1 NOT_274( .ZN(n177gat), .A(II651) );
  INV_X1 NOT_275( .ZN(n54gat), .A(n167gat) );
  INV_X1 NOT_276( .ZN(II658), .A(n54gat) );
  INV_X1 NOT_277( .ZN(n60gat), .A(II658) );
  INV_X1 NOT_278( .ZN(II661), .A(n845gat) );
  INV_X1 NOT_279( .ZN(n911gat), .A(II661) );
  INV_X1 NOT_280( .ZN(II672), .A(n1026gat) );
  INV_X1 NOT_281( .ZN(n1025gat), .A(II672) );
  INV_X1 NOT_282( .ZN(II675), .A(n1025gat) );
  INV_X1 NOT_283( .ZN(n912gat), .A(II675) );
  INV_X8 NOT_284( .ZN(II678), .A(n918gat) );
  INV_X1 NOT_285( .ZN(n913gat), .A(II678) );
  INV_X1 NOT_286( .ZN(n1024gat), .A(n1026gat) );
  INV_X4 NOT_287( .ZN(II683), .A(n1024gat) );
  INV_X1 NOT_288( .ZN(n914gat), .A(II683) );
  INV_X1 NOT_289( .ZN(n917gat), .A(n919gat) );
  INV_X1 NOT_290( .ZN(II687), .A(n917gat) );
  INV_X1 NOT_291( .ZN(n915gat), .A(II687) );
  INV_X1 NOT_292( .ZN(n844gat), .A(n846gat) );
  INV_X1 NOT_293( .ZN(II692), .A(n844gat) );
  INV_X1 NOT_294( .ZN(n916gat), .A(II692) );
  INV_X1 NOT_295( .ZN(II698), .A(n906gat) );
  INV_X1 NOT_296( .ZN(n61gat), .A(II698) );
  INV_X1 NOT_297( .ZN(II709), .A(n275gat) );
  INV_X1 NOT_298( .ZN(n274gat), .A(II709) );
  INV_X1 NOT_299( .ZN(II712), .A(n274gat) );
  INV_X1 NOT_300( .ZN(n348gat), .A(II712) );
  INV_X1 NOT_301( .ZN(II715), .A(n401gat) );
  INV_X1 NOT_302( .ZN(n349gat), .A(II715) );
  INV_X1 NOT_303( .ZN(II718), .A(n398gat) );
  INV_X1 NOT_304( .ZN(n397gat), .A(II718) );
  INV_X1 NOT_305( .ZN(II721), .A(n397gat) );
  INV_X1 NOT_306( .ZN(n350gat), .A(II721) );
  INV_X1 NOT_307( .ZN(n400gat), .A(n402gat) );
  INV_X1 NOT_308( .ZN(II726), .A(n400gat) );
  INV_X1 NOT_309( .ZN(n351gat), .A(II726) );
  INV_X1 NOT_310( .ZN(II729), .A(n396gat) );
  INV_X1 NOT_311( .ZN(n352gat), .A(II729) );
  INV_X1 NOT_312( .ZN(n273gat), .A(n275gat) );
  INV_X1 NOT_313( .ZN(II734), .A(n273gat) );
  INV_X1 NOT_314( .ZN(n353gat), .A(II734) );
  INV_X1 NOT_315( .ZN(n178gat), .A(n343gat) );
  INV_X1 NOT_316( .ZN(II741), .A(n178gat) );
  INV_X1 NOT_317( .ZN(n62gat), .A(II741) );
  INV_X1 NOT_318( .ZN(n66gat), .A(n906gat) );
  INV_X1 NOT_319( .ZN(II746), .A(n66gat) );
  INV_X1 NOT_320( .ZN(n63gat), .A(II746) );
  INV_X1 NOT_321( .ZN(II749), .A(n343gat) );
  INV_X1 NOT_322( .ZN(n64gat), .A(II749) );
  INV_X1 NOT_323( .ZN(II753), .A(n167gat) );
  INV_X1 NOT_324( .ZN(n65gat), .A(II753) );
  INV_X1 NOT_325( .ZN(n2474gat), .A(n2476gat) );
  INV_X1 NOT_326( .ZN(II768), .A(n3090gat) );
  INV_X4 NOT_327( .ZN(n2832gat), .A(II768) );
  INV_X4 NOT_328( .ZN(II771), .A(n2832gat) );
  INV_X1 NOT_329( .ZN(n2831gat), .A(II771) );
  INV_X1 NOT_330( .ZN(n2731gat), .A(n2733gat) );
  INV_X1 NOT_331( .ZN(II776), .A(n3074gat) );
  INV_X1 NOT_332( .ZN(n2719gat), .A(II776) );
  INV_X1 NOT_333( .ZN(n2718gat), .A(n2719gat) );
  INV_X1 NOT_334( .ZN(II790), .A(n1068gat) );
  INV_X1 NOT_335( .ZN(n1067gat), .A(II790) );
  INV_X1 NOT_336( .ZN(II793), .A(n1067gat) );
  INV_X1 NOT_337( .ZN(n949gat), .A(II793) );
  INV_X1 NOT_338( .ZN(II796), .A(n3076gat) );
  INV_X1 NOT_339( .ZN(n2839gat), .A(II796) );
  INV_X1 NOT_340( .ZN(n2838gat), .A(n2839gat) );
  INV_X1 NOT_341( .ZN(n2775gat), .A(n2777gat) );
  INV_X1 NOT_342( .ZN(II812), .A(n957gat) );
  INV_X1 NOT_343( .ZN(n956gat), .A(II812) );
  INV_X1 NOT_344( .ZN(II815), .A(n956gat) );
  INV_X1 NOT_345( .ZN(n950gat), .A(II815) );
  INV_X1 NOT_346( .ZN(II818), .A(n3075gat) );
  INV_X1 NOT_347( .ZN(n2712gat), .A(II818) );
  INV_X1 NOT_348( .ZN(n2711gat), .A(n2712gat) );
  INV_X1 NOT_349( .ZN(n2734gat), .A(n2736gat) );
  INV_X1 NOT_350( .ZN(II834), .A(n861gat) );
  INV_X1 NOT_351( .ZN(n860gat), .A(II834) );
  INV_X1 NOT_352( .ZN(II837), .A(n860gat) );
  INV_X1 NOT_353( .ZN(n951gat), .A(II837) );
  INV_X1 NOT_354( .ZN(n955gat), .A(n957gat) );
  INV_X1 NOT_355( .ZN(II842), .A(n955gat) );
  INV_X1 NOT_356( .ZN(n952gat), .A(II842) );
  INV_X1 NOT_357( .ZN(n859gat), .A(n861gat) );
  INV_X1 NOT_358( .ZN(II846), .A(n859gat) );
  INV_X1 NOT_359( .ZN(n953gat), .A(II846) );
  INV_X1 NOT_360( .ZN(n1066gat), .A(n1068gat) );
  INV_X1 NOT_361( .ZN(II851), .A(n1066gat) );
  INV_X1 NOT_362( .ZN(n954gat), .A(II851) );
  INV_X1 NOT_363( .ZN(n857gat), .A(n944gat) );
  INV_X1 NOT_364( .ZN(II858), .A(n857gat) );
  INV_X1 NOT_365( .ZN(n938gat), .A(II858) );
  INV_X1 NOT_366( .ZN(n2792gat), .A(n2794gat) );
  INV_X1 NOT_367( .ZN(II863), .A(n3080gat) );
  INV_X1 NOT_368( .ZN(n2847gat), .A(II863) );
  INV_X1 NOT_369( .ZN(n2846gat), .A(n2847gat) );
  INV_X1 NOT_370( .ZN(II877), .A(n1294gat) );
  INV_X1 NOT_371( .ZN(n1293gat), .A(II877) );
  INV_X1 NOT_372( .ZN(II880), .A(n1293gat) );
  INV_X1 NOT_373( .ZN(n1233gat), .A(II880) );
  INV_X1 NOT_374( .ZN(n2672gat), .A(n2674gat) );
  INV_X1 NOT_375( .ZN(II885), .A(n3082gat) );
  INV_X1 NOT_376( .ZN(n2853gat), .A(II885) );
  INV_X1 NOT_377( .ZN(n2852gat), .A(n2853gat) );
  INV_X1 NOT_378( .ZN(II899), .A(n1241gat) );
  INV_X1 NOT_379( .ZN(n1240gat), .A(II899) );
  INV_X1 NOT_380( .ZN(II902), .A(n1240gat) );
  INV_X1 NOT_381( .ZN(n1234gat), .A(II902) );
  INV_X1 NOT_382( .ZN(II913), .A(n1298gat) );
  INV_X1 NOT_383( .ZN(n1297gat), .A(II913) );
  INV_X1 NOT_384( .ZN(II916), .A(n1297gat) );
  INV_X1 NOT_385( .ZN(n1235gat), .A(II916) );
  INV_X1 NOT_386( .ZN(n1239gat), .A(n1241gat) );
  INV_X1 NOT_387( .ZN(II921), .A(n1239gat) );
  INV_X1 NOT_388( .ZN(n1236gat), .A(II921) );
  INV_X1 NOT_389( .ZN(n1296gat), .A(n1298gat) );
  INV_X1 NOT_390( .ZN(II925), .A(n1296gat) );
  INV_X1 NOT_391( .ZN(n1237gat), .A(II925) );
  INV_X1 NOT_392( .ZN(n1292gat), .A(n1294gat) );
  INV_X1 NOT_393( .ZN(II930), .A(n1292gat) );
  INV_X1 NOT_394( .ZN(n1238gat), .A(II930) );
  INV_X1 NOT_395( .ZN(II936), .A(n1228gat) );
  INV_X1 NOT_396( .ZN(n939gat), .A(II936) );
  INV_X1 NOT_397( .ZN(n2778gat), .A(n2780gat) );
  INV_X1 NOT_398( .ZN(II941), .A(n3077gat) );
  INV_X2 NOT_399( .ZN(n2837gat), .A(II941) );
  INV_X2 NOT_400( .ZN(n2836gat), .A(n2837gat) );
  INV_X1 NOT_401( .ZN(II955), .A(n865gat) );
  INV_X1 NOT_402( .ZN(n864gat), .A(II955) );
  INV_X1 NOT_403( .ZN(II958), .A(n864gat) );
  INV_X1 NOT_404( .ZN(n1055gat), .A(II958) );
  INV_X1 NOT_405( .ZN(n2789gat), .A(n2791gat) );
  INV_X1 NOT_406( .ZN(II963), .A(n3079gat) );
  INV_X1 NOT_407( .ZN(n2841gat), .A(II963) );
  INV_X1 NOT_408( .ZN(n2840gat), .A(n2841gat) );
  INV_X1 NOT_409( .ZN(II977), .A(n1080gat) );
  INV_X1 NOT_410( .ZN(n1079gat), .A(II977) );
  INV_X1 NOT_411( .ZN(II980), .A(n1079gat) );
  INV_X1 NOT_412( .ZN(n1056gat), .A(II980) );
  INV_X1 NOT_413( .ZN(n2781gat), .A(n2783gat) );
  INV_X1 NOT_414( .ZN(II985), .A(n3078gat) );
  INV_X1 NOT_415( .ZN(n2843gat), .A(II985) );
  INV_X1 NOT_416( .ZN(n2842gat), .A(n2843gat) );
  INV_X1 NOT_417( .ZN(II999), .A(n1148gat) );
  INV_X1 NOT_418( .ZN(n1147gat), .A(II999) );
  INV_X1 NOT_419( .ZN(II1002), .A(n1147gat) );
  INV_X1 NOT_420( .ZN(n1057gat), .A(II1002) );
  INV_X1 NOT_421( .ZN(n1078gat), .A(n1080gat) );
  INV_X1 NOT_422( .ZN(II1007), .A(n1078gat) );
  INV_X1 NOT_423( .ZN(n1058gat), .A(II1007) );
  INV_X1 NOT_424( .ZN(n1146gat), .A(n1148gat) );
  INV_X1 NOT_425( .ZN(II1011), .A(n1146gat) );
  INV_X1 NOT_426( .ZN(n1059gat), .A(II1011) );
  INV_X1 NOT_427( .ZN(n863gat), .A(n865gat) );
  INV_X1 NOT_428( .ZN(II1016), .A(n863gat) );
  INV_X1 NOT_429( .ZN(n1060gat), .A(II1016) );
  INV_X1 NOT_430( .ZN(n928gat), .A(n1050gat) );
  INV_X1 NOT_431( .ZN(II1023), .A(n928gat) );
  INV_X1 NOT_432( .ZN(n940gat), .A(II1023) );
  INV_X1 NOT_433( .ZN(n858gat), .A(n1228gat) );
  INV_X1 NOT_434( .ZN(II1028), .A(n858gat) );
  INV_X1 NOT_435( .ZN(n941gat), .A(II1028) );
  INV_X1 NOT_436( .ZN(II1031), .A(n1050gat) );
  INV_X1 NOT_437( .ZN(n942gat), .A(II1031) );
  INV_X1 NOT_438( .ZN(II1035), .A(n944gat) );
  INV_X1 NOT_439( .ZN(n943gat), .A(II1035) );
  INV_X1 NOT_440( .ZN(n2466gat), .A(n2468gat) );
  INV_X1 NOT_441( .ZN(n2720gat), .A(n2722gat) );
  INV_X1 NOT_442( .ZN(n740gat), .A(n2667gat) );
  INV_X1 NOT_443( .ZN(n2784gat), .A(n2786gat) );
  INV_X1 NOT_444( .ZN(n743gat), .A(n746gat) );
  INV_X1 NOT_445( .ZN(n294gat), .A(n360gat) );
  INV_X1 NOT_446( .ZN(n374gat), .A(n2767gat) );
  INV_X1 NOT_447( .ZN(n616gat), .A(n618gat) );
  INV_X1 NOT_448( .ZN(II1067), .A(n616gat) );
  INV_X1 NOT_449( .ZN(n501gat), .A(II1067) );
  INV_X2 NOT_450( .ZN(n489gat), .A(n491gat) );
  INV_X1 NOT_451( .ZN(II1079), .A(n489gat) );
  INV_X1 NOT_452( .ZN(n502gat), .A(II1079) );
  INV_X1 NOT_453( .ZN(II1082), .A(n618gat) );
  INV_X1 NOT_454( .ZN(n617gat), .A(II1082) );
  INV_X1 NOT_455( .ZN(II1085), .A(n617gat) );
  INV_X1 NOT_456( .ZN(n499gat), .A(II1085) );
  INV_X1 NOT_457( .ZN(II1088), .A(n491gat) );
  INV_X1 NOT_458( .ZN(n490gat), .A(II1088) );
  INV_X1 NOT_459( .ZN(II1091), .A(n490gat) );
  INV_X1 NOT_460( .ZN(n500gat), .A(II1091) );
  INV_X1 NOT_461( .ZN(n620gat), .A(n622gat) );
  INV_X1 NOT_462( .ZN(II1103), .A(n620gat) );
  INV_X1 NOT_463( .ZN(n738gat), .A(II1103) );
  INV_X4 NOT_464( .ZN(n624gat), .A(n626gat) );
  INV_X1 NOT_465( .ZN(II1115), .A(n624gat) );
  INV_X1 NOT_466( .ZN(n737gat), .A(II1115) );
  INV_X1 NOT_467( .ZN(II1118), .A(n622gat) );
  INV_X1 NOT_468( .ZN(n621gat), .A(II1118) );
  INV_X1 NOT_469( .ZN(II1121), .A(n621gat) );
  INV_X1 NOT_470( .ZN(n733gat), .A(II1121) );
  INV_X1 NOT_471( .ZN(II1124), .A(n626gat) );
  INV_X1 NOT_472( .ZN(n625gat), .A(II1124) );
  INV_X1 NOT_473( .ZN(II1127), .A(n625gat) );
  INV_X1 NOT_474( .ZN(n735gat), .A(II1127) );
  INV_X1 NOT_475( .ZN(II1138), .A(n834gat) );
  INV_X1 NOT_476( .ZN(n833gat), .A(II1138) );
  INV_X1 NOT_477( .ZN(II1141), .A(n833gat) );
  INV_X1 NOT_478( .ZN(n714gat), .A(II1141) );
  INV_X1 NOT_479( .ZN(II1152), .A(n707gat) );
  INV_X1 NOT_480( .ZN(n706gat), .A(II1152) );
  INV_X1 NOT_481( .ZN(II1155), .A(n706gat) );
  INV_X1 NOT_482( .ZN(n715gat), .A(II1155) );
  INV_X2 NOT_483( .ZN(II1166), .A(n838gat) );
  INV_X1 NOT_484( .ZN(n837gat), .A(II1166) );
  INV_X1 NOT_485( .ZN(II1169), .A(n837gat) );
  INV_X1 NOT_486( .ZN(n716gat), .A(II1169) );
  INV_X1 NOT_487( .ZN(n705gat), .A(n707gat) );
  INV_X1 NOT_488( .ZN(II1174), .A(n705gat) );
  INV_X1 NOT_489( .ZN(n717gat), .A(II1174) );
  INV_X1 NOT_490( .ZN(n836gat), .A(n838gat) );
  INV_X1 NOT_491( .ZN(II1178), .A(n836gat) );
  INV_X1 NOT_492( .ZN(n718gat), .A(II1178) );
  INV_X1 NOT_493( .ZN(n832gat), .A(n834gat) );
  INV_X1 NOT_494( .ZN(II1183), .A(n832gat) );
  INV_X1 NOT_495( .ZN(n719gat), .A(II1183) );
  INV_X1 NOT_496( .ZN(n515gat), .A(n709gat) );
  INV_X1 NOT_497( .ZN(II1190), .A(n515gat) );
  INV_X1 NOT_498( .ZN(n509gat), .A(II1190) );
  INV_X1 NOT_499( .ZN(II1201), .A(n830gat) );
  INV_X1 NOT_500( .ZN(n829gat), .A(II1201) );
  INV_X1 NOT_501( .ZN(II1204), .A(n829gat) );
  INV_X1 NOT_502( .ZN(n734gat), .A(II1204) );
  INV_X1 NOT_503( .ZN(n828gat), .A(n830gat) );
  INV_X1 NOT_504( .ZN(II1209), .A(n828gat) );
  INV_X1 NOT_505( .ZN(n736gat), .A(II1209) );
  INV_X8 NOT_506( .ZN(II1216), .A(n728gat) );
  INV_X1 NOT_507( .ZN(n510gat), .A(II1216) );
  INV_X1 NOT_508( .ZN(II1227), .A(n614gat) );
  INV_X1 NOT_509( .ZN(n613gat), .A(II1227) );
  INV_X1 NOT_510( .ZN(II1230), .A(n613gat) );
  INV_X1 NOT_511( .ZN(n498gat), .A(II1230) );
  INV_X1 NOT_512( .ZN(n612gat), .A(n614gat) );
  INV_X1 NOT_513( .ZN(II1236), .A(n612gat) );
  INV_X1 NOT_514( .ZN(n503gat), .A(II1236) );
  INV_X1 NOT_515( .ZN(n404gat), .A(n493gat) );
  INV_X1 NOT_516( .ZN(II1243), .A(n404gat) );
  INV_X1 NOT_517( .ZN(n511gat), .A(II1243) );
  INV_X1 NOT_518( .ZN(n405gat), .A(n728gat) );
  INV_X1 NOT_519( .ZN(II1248), .A(n405gat) );
  INV_X1 NOT_520( .ZN(n512gat), .A(II1248) );
  INV_X1 NOT_521( .ZN(II1251), .A(n493gat) );
  INV_X1 NOT_522( .ZN(n513gat), .A(II1251) );
  INV_X1 NOT_523( .ZN(II1255), .A(n709gat) );
  INV_X1 NOT_524( .ZN(n514gat), .A(II1255) );
  INV_X1 NOT_525( .ZN(n2524gat), .A(n2526gat) );
  INV_X1 NOT_526( .ZN(n17gat), .A(n564gat) );
  INV_X1 NOT_527( .ZN(n79gat), .A(n86gat) );
  INV_X1 NOT_528( .ZN(n219gat), .A(n78gat) );
  INV_X1 NOT_529( .ZN(n563gat), .A(II1278) );
  INV_X1 NOT_530( .ZN(n289gat), .A(n563gat) );
  INV_X1 NOT_531( .ZN(n179gat), .A(n287gat) );
  INV_X1 NOT_532( .ZN(n188gat), .A(n288gat) );
  INV_X1 NOT_533( .ZN(n72gat), .A(n181gat) );
  INV_X1 NOT_534( .ZN(n111gat), .A(n182gat) );
  INV_X1 NOT_535( .ZN(II1302), .A(n680gat) );
  INV_X1 NOT_536( .ZN(n679gat), .A(II1302) );
  INV_X1 NOT_537( .ZN(II1305), .A(n679gat) );
  INV_X1 NOT_538( .ZN(n808gat), .A(II1305) );
  INV_X1 NOT_539( .ZN(II1319), .A(n816gat) );
  INV_X1 NOT_540( .ZN(n815gat), .A(II1319) );
  INV_X1 NOT_541( .ZN(II1322), .A(n815gat) );
  INV_X1 NOT_542( .ZN(n809gat), .A(II1322) );
  INV_X1 NOT_543( .ZN(II1336), .A(n580gat) );
  INV_X1 NOT_544( .ZN(n579gat), .A(II1336) );
  INV_X1 NOT_545( .ZN(II1339), .A(n579gat) );
  INV_X1 NOT_546( .ZN(n810gat), .A(II1339) );
  INV_X16 NOT_547( .ZN(n814gat), .A(n816gat) );
  INV_X1 NOT_548( .ZN(II1344), .A(n814gat) );
  INV_X1 NOT_549( .ZN(n811gat), .A(II1344) );
  INV_X1 NOT_550( .ZN(n578gat), .A(n580gat) );
  INV_X1 NOT_551( .ZN(II1348), .A(n578gat) );
  INV_X1 NOT_552( .ZN(n812gat), .A(II1348) );
  INV_X1 NOT_553( .ZN(n678gat), .A(n680gat) );
  INV_X1 NOT_554( .ZN(II1353), .A(n678gat) );
  INV_X1 NOT_555( .ZN(n813gat), .A(II1353) );
  INV_X1 NOT_556( .ZN(n677gat), .A(n803gat) );
  INV_X1 NOT_557( .ZN(II1360), .A(n677gat) );
  INV_X1 NOT_558( .ZN(n572gat), .A(II1360) );
  INV_X1 NOT_559( .ZN(II1371), .A(n824gat) );
  INV_X1 NOT_560( .ZN(n823gat), .A(II1371) );
  INV_X1 NOT_561( .ZN(II1374), .A(n823gat) );
  INV_X1 NOT_562( .ZN(n591gat), .A(II1374) );
  INV_X1 NOT_563( .ZN(II1385), .A(n820gat) );
  INV_X1 NOT_564( .ZN(n819gat), .A(II1385) );
  INV_X1 NOT_565( .ZN(II1388), .A(n819gat) );
  INV_X1 NOT_566( .ZN(n592gat), .A(II1388) );
  INV_X1 NOT_567( .ZN(II1399), .A(n883gat) );
  INV_X1 NOT_568( .ZN(n882gat), .A(II1399) );
  INV_X1 NOT_569( .ZN(II1402), .A(n882gat) );
  INV_X1 NOT_570( .ZN(n593gat), .A(II1402) );
  INV_X1 NOT_571( .ZN(n818gat), .A(n820gat) );
  INV_X16 NOT_572( .ZN(II1407), .A(n818gat) );
  INV_X1 NOT_573( .ZN(n594gat), .A(II1407) );
  INV_X1 NOT_574( .ZN(n881gat), .A(n883gat) );
  INV_X1 NOT_575( .ZN(II1411), .A(n881gat) );
  INV_X1 NOT_576( .ZN(n595gat), .A(II1411) );
  INV_X1 NOT_577( .ZN(n822gat), .A(n824gat) );
  INV_X1 NOT_578( .ZN(II1416), .A(n822gat) );
  INV_X1 NOT_579( .ZN(n596gat), .A(II1416) );
  INV_X1 NOT_580( .ZN(II1422), .A(n586gat) );
  INV_X1 NOT_581( .ZN(n573gat), .A(II1422) );
  INV_X1 NOT_582( .ZN(II1436), .A(n584gat) );
  INV_X1 NOT_583( .ZN(n583gat), .A(II1436) );
  INV_X1 NOT_584( .ZN(II1439), .A(n583gat) );
  INV_X1 NOT_585( .ZN(n691gat), .A(II1439) );
  INV_X1 NOT_586( .ZN(II1450), .A(n684gat) );
  INV_X1 NOT_587( .ZN(n683gat), .A(II1450) );
  INV_X1 NOT_588( .ZN(II1453), .A(n683gat) );
  INV_X1 NOT_589( .ZN(n692gat), .A(II1453) );
  INV_X1 NOT_590( .ZN(II1464), .A(n699gat) );
  INV_X1 NOT_591( .ZN(n698gat), .A(II1464) );
  INV_X1 NOT_592( .ZN(II1467), .A(n698gat) );
  INV_X1 NOT_593( .ZN(n693gat), .A(II1467) );
  INV_X1 NOT_594( .ZN(n682gat), .A(n684gat) );
  INV_X1 NOT_595( .ZN(II1472), .A(n682gat) );
  INV_X1 NOT_596( .ZN(n694gat), .A(II1472) );
  INV_X1 NOT_597( .ZN(n697gat), .A(n699gat) );
  INV_X1 NOT_598( .ZN(II1476), .A(n697gat) );
  INV_X1 NOT_599( .ZN(n695gat), .A(II1476) );
  INV_X1 NOT_600( .ZN(n582gat), .A(n584gat) );
  INV_X2 NOT_601( .ZN(II1481), .A(n582gat) );
  INV_X1 NOT_602( .ZN(n696gat), .A(II1481) );
  INV_X1 NOT_603( .ZN(n456gat), .A(n686gat) );
  INV_X1 NOT_604( .ZN(II1488), .A(n456gat) );
  INV_X1 NOT_605( .ZN(n574gat), .A(II1488) );
  INV_X1 NOT_606( .ZN(n565gat), .A(n586gat) );
  INV_X1 NOT_607( .ZN(II1493), .A(n565gat) );
  INV_X2 NOT_608( .ZN(n575gat), .A(II1493) );
  INV_X1 NOT_609( .ZN(II1496), .A(n686gat) );
  INV_X1 NOT_610( .ZN(n576gat), .A(II1496) );
  INV_X1 NOT_611( .ZN(II1500), .A(n803gat) );
  INV_X1 NOT_612( .ZN(n577gat), .A(II1500) );
  INV_X1 NOT_613( .ZN(n2462gat), .A(n2464gat) );
  INV_X1 NOT_614( .ZN(n2665gat), .A(II1516) );
  INV_X1 NOT_615( .ZN(n2596gat), .A(n2665gat) );
  INV_X1 NOT_616( .ZN(n189gat), .A(n286gat) );
  INV_X1 NOT_617( .ZN(n194gat), .A(n187gat) );
  INV_X1 NOT_618( .ZN(n21gat), .A(n15gat) );
  INV_X1 NOT_619( .ZN(II1538), .A(n2399gat) );
  INV_X1 NOT_620( .ZN(n2398gat), .A(II1538) );
  INV_X1 NOT_621( .ZN(n2353gat), .A(n2398gat) );
  INV_X1 NOT_622( .ZN(II1550), .A(n2343gat) );
  INV_X1 NOT_623( .ZN(n2342gat), .A(II1550) );
  INV_X1 NOT_624( .ZN(n2284gat), .A(n2342gat) );
  INV_X1 NOT_625( .ZN(n2201gat), .A(n2203gat) );
  INV_X1 NOT_626( .ZN(n2354gat), .A(n2201gat) );
  INV_X1 NOT_627( .ZN(n2560gat), .A(n2562gat) );
  INV_X1 NOT_628( .ZN(n2356gat), .A(n2560gat) );
  INV_X1 NOT_629( .ZN(n2205gat), .A(n2207gat) );
  INV_X1 NOT_630( .ZN(n2214gat), .A(n2205gat) );
  INV_X1 NOT_631( .ZN(n2286gat), .A(II1585) );
  INV_X1 NOT_632( .ZN(n2624gat), .A(n2626gat) );
  INV_X1 NOT_633( .ZN(II1606), .A(n2490gat) );
  INV_X1 NOT_634( .ZN(n2489gat), .A(II1606) );
  INV_X1 NOT_635( .ZN(II1617), .A(n2622gat) );
  INV_X1 NOT_636( .ZN(n2621gat), .A(II1617) );
  INV_X1 NOT_637( .ZN(n2533gat), .A(n2534gat) );
  INV_X1 NOT_638( .ZN(II1630), .A(n2630gat) );
  INV_X1 NOT_639( .ZN(n2629gat), .A(II1630) );
  INV_X1 NOT_640( .ZN(n2486gat), .A(n2629gat) );
  INV_X1 NOT_641( .ZN(n2541gat), .A(n2543gat) );
  INV_X1 NOT_642( .ZN(n2429gat), .A(n2541gat) );
  INV_X1 NOT_643( .ZN(n2432gat), .A(n2430gat) );
  INV_X1 NOT_644( .ZN(II1655), .A(n2102gat) );
  INV_X1 NOT_645( .ZN(n2101gat), .A(II1655) );
  INV_X1 NOT_646( .ZN(n1693gat), .A(n2101gat) );
  INV_X1 NOT_647( .ZN(II1667), .A(n1880gat) );
  INV_X1 NOT_648( .ZN(n1879gat), .A(II1667) );
  INV_X1 NOT_649( .ZN(n1698gat), .A(n1934gat) );
  INV_X1 NOT_650( .ZN(n1543gat), .A(n1606gat) );
  INV_X1 NOT_651( .ZN(II1683), .A(n1763gat) );
  INV_X1 NOT_652( .ZN(n1762gat), .A(II1683) );
  INV_X1 NOT_653( .ZN(n1673gat), .A(n2989gat) );
  INV_X1 NOT_654( .ZN(n1858gat), .A(n1673gat) );
  INV_X1 NOT_655( .ZN(II1698), .A(n2155gat) );
  INV_X1 NOT_656( .ZN(n2154gat), .A(II1698) );
  INV_X1 NOT_657( .ZN(n2488gat), .A(n2490gat) );
  INV_X1 NOT_658( .ZN(II1703), .A(n2626gat) );
  INV_X4 NOT_659( .ZN(n2625gat), .A(II1703) );
  INV_X1 NOT_660( .ZN(n2530gat), .A(n2531gat) );
  INV_X1 NOT_661( .ZN(II1708), .A(n2543gat) );
  INV_X1 NOT_662( .ZN(n2542gat), .A(II1708) );
  INV_X1 NOT_663( .ZN(n2482gat), .A(n2542gat) );
  INV_X1 NOT_664( .ZN(n2426gat), .A(n2480gat) );
  INV_X1 NOT_665( .ZN(n2153gat), .A(n2155gat) );
  INV_X1 NOT_666( .ZN(n2341gat), .A(n2343gat) );
  INV_X1 NOT_667( .ZN(n2355gat), .A(n2341gat) );
  INV_X1 NOT_668( .ZN(II1719), .A(n2562gat) );
  INV_X2 NOT_669( .ZN(n2561gat), .A(II1719) );
  INV_X1 NOT_670( .ZN(n2443gat), .A(n2561gat) );
  INV_X1 NOT_671( .ZN(n2289gat), .A(II1724) );
  INV_X1 NOT_672( .ZN(n2148gat), .A(II1734) );
  INV_X1 NOT_673( .ZN(n855gat), .A(n2148gat) );
  INV_X1 NOT_674( .ZN(n759gat), .A(n855gat) );
  INV_X1 NOT_675( .ZN(II1749), .A(n1035gat) );
  INV_X1 NOT_676( .ZN(n1034gat), .A(II1749) );
  INV_X1 NOT_677( .ZN(II1752), .A(n1034gat) );
  INV_X1 NOT_678( .ZN(n1189gat), .A(II1752) );
  INV_X1 NOT_679( .ZN(n1075gat), .A(n855gat) );
  INV_X1 NOT_680( .ZN(II1766), .A(n1121gat) );
  INV_X1 NOT_681( .ZN(n1120gat), .A(II1766) );
  INV_X1 NOT_682( .ZN(II1769), .A(n1120gat) );
  INV_X1 NOT_683( .ZN(n1190gat), .A(II1769) );
  INV_X1 NOT_684( .ZN(n760gat), .A(n855gat) );
  INV_X1 NOT_685( .ZN(II1783), .A(n1072gat) );
  INV_X1 NOT_686( .ZN(n1071gat), .A(II1783) );
  INV_X1 NOT_687( .ZN(II1786), .A(n1071gat) );
  INV_X1 NOT_688( .ZN(n1191gat), .A(II1786) );
  INV_X1 NOT_689( .ZN(n1119gat), .A(n1121gat) );
  INV_X1 NOT_690( .ZN(II1791), .A(n1119gat) );
  INV_X1 NOT_691( .ZN(n1192gat), .A(II1791) );
  INV_X1 NOT_692( .ZN(n1070gat), .A(n1072gat) );
  INV_X1 NOT_693( .ZN(II1795), .A(n1070gat) );
  INV_X1 NOT_694( .ZN(n1193gat), .A(II1795) );
  INV_X1 NOT_695( .ZN(n1033gat), .A(n1035gat) );
  INV_X1 NOT_696( .ZN(II1800), .A(n1033gat) );
  INV_X1 NOT_697( .ZN(n1194gat), .A(II1800) );
  INV_X1 NOT_698( .ZN(n1183gat), .A(n1184gat) );
  INV_X1 NOT_699( .ZN(II1807), .A(n1183gat) );
  INV_X1 NOT_700( .ZN(n1274gat), .A(II1807) );
  INV_X1 NOT_701( .ZN(n644gat), .A(n855gat) );
  INV_X1 NOT_702( .ZN(n1280gat), .A(n1282gat) );
  INV_X1 NOT_703( .ZN(n641gat), .A(n855gat) );
  INV_X1 NOT_704( .ZN(II1833), .A(n1226gat) );
  INV_X1 NOT_705( .ZN(n1225gat), .A(II1833) );
  INV_X1 NOT_706( .ZN(II1837), .A(n1282gat) );
  INV_X1 NOT_707( .ZN(n1281gat), .A(II1837) );
  INV_X1 NOT_708( .ZN(n1224gat), .A(n1226gat) );
  INV_X1 NOT_709( .ZN(II1843), .A(n2970gat) );
  INV_X1 NOT_710( .ZN(n1275gat), .A(II1843) );
  INV_X1 NOT_711( .ZN(n761gat), .A(n855gat) );
  INV_X1 NOT_712( .ZN(II1857), .A(n931gat) );
  INV_X1 NOT_713( .ZN(n930gat), .A(II1857) );
  INV_X1 NOT_714( .ZN(II1860), .A(n930gat) );
  INV_X1 NOT_715( .ZN(n1206gat), .A(II1860) );
  INV_X1 NOT_716( .ZN(n762gat), .A(n855gat) );
  INV_X1 NOT_717( .ZN(II1874), .A(n1135gat) );
  INV_X1 NOT_718( .ZN(n1134gat), .A(II1874) );
  INV_X1 NOT_719( .ZN(II1877), .A(n1134gat) );
  INV_X1 NOT_720( .ZN(n1207gat), .A(II1877) );
  INV_X1 NOT_721( .ZN(n643gat), .A(n855gat) );
  INV_X1 NOT_722( .ZN(II1891), .A(n1045gat) );
  INV_X1 NOT_723( .ZN(n1044gat), .A(II1891) );
  INV_X1 NOT_724( .ZN(II1894), .A(n1044gat) );
  INV_X2 NOT_725( .ZN(n1208gat), .A(II1894) );
  INV_X2 NOT_726( .ZN(n1133gat), .A(n1135gat) );
  INV_X1 NOT_727( .ZN(II1899), .A(n1133gat) );
  INV_X1 NOT_728( .ZN(n1209gat), .A(II1899) );
  INV_X1 NOT_729( .ZN(n1043gat), .A(n1045gat) );
  INV_X1 NOT_730( .ZN(II1903), .A(n1043gat) );
  INV_X1 NOT_731( .ZN(n1210gat), .A(II1903) );
  INV_X1 NOT_732( .ZN(n929gat), .A(n931gat) );
  INV_X1 NOT_733( .ZN(II1908), .A(n929gat) );
  INV_X1 NOT_734( .ZN(n1211gat), .A(II1908) );
  INV_X1 NOT_735( .ZN(n1268gat), .A(n1201gat) );
  INV_X1 NOT_736( .ZN(II1915), .A(n1268gat) );
  INV_X1 NOT_737( .ZN(n1276gat), .A(II1915) );
  INV_X1 NOT_738( .ZN(n1329gat), .A(n2970gat) );
  INV_X1 NOT_739( .ZN(II1920), .A(n1329gat) );
  INV_X1 NOT_740( .ZN(n1277gat), .A(II1920) );
  INV_X1 NOT_741( .ZN(II1923), .A(n1201gat) );
  INV_X1 NOT_742( .ZN(n1278gat), .A(II1923) );
  INV_X1 NOT_743( .ZN(II1927), .A(n1184gat) );
  INV_X1 NOT_744( .ZN(n1279gat), .A(II1927) );
  INV_X1 NOT_745( .ZN(n1284gat), .A(n1269gat) );
  INV_X1 NOT_746( .ZN(n642gat), .A(n855gat) );
  INV_X1 NOT_747( .ZN(n1195gat), .A(n1197gat) );
  INV_X1 NOT_748( .ZN(II1947), .A(n1197gat) );
  INV_X1 NOT_749( .ZN(n1196gat), .A(II1947) );
  INV_X1 NOT_750( .ZN(n2516gat), .A(n2518gat) );
  INV_X1 NOT_751( .ZN(II1961), .A(n2516gat) );
  INV_X1 NOT_752( .ZN(n3017gat), .A(II1961) );
  INV_X1 NOT_753( .ZN(n851gat), .A(n853gat) );
  INV_X1 NOT_754( .ZN(n1725gat), .A(n2148gat) );
  INV_X1 NOT_755( .ZN(n664gat), .A(n1725gat) );
  INV_X1 NOT_756( .ZN(n852gat), .A(n854gat) );
  INV_X1 NOT_757( .ZN(II1981), .A(n667gat) );
  INV_X1 NOT_758( .ZN(n666gat), .A(II1981) );
  INV_X1 NOT_759( .ZN(n368gat), .A(n1725gat) );
  INV_X1 NOT_760( .ZN(II1996), .A(n659gat) );
  INV_X1 NOT_761( .ZN(n658gat), .A(II1996) );
  INV_X1 NOT_762( .ZN(II1999), .A(n658gat) );
  INV_X1 NOT_763( .ZN(n784gat), .A(II1999) );
  INV_X1 NOT_764( .ZN(n662gat), .A(n1725gat) );
  INV_X1 NOT_765( .ZN(II2014), .A(n553gat) );
  INV_X1 NOT_766( .ZN(n552gat), .A(II2014) );
  INV_X1 NOT_767( .ZN(II2017), .A(n552gat) );
  INV_X1 NOT_768( .ZN(n785gat), .A(II2017) );
  INV_X1 NOT_769( .ZN(n661gat), .A(n1725gat) );
  INV_X1 NOT_770( .ZN(II2032), .A(n777gat) );
  INV_X1 NOT_771( .ZN(n776gat), .A(II2032) );
  INV_X1 NOT_772( .ZN(II2035), .A(n776gat) );
  INV_X1 NOT_773( .ZN(n786gat), .A(II2035) );
  INV_X1 NOT_774( .ZN(n551gat), .A(n553gat) );
  INV_X1 NOT_775( .ZN(II2040), .A(n551gat) );
  INV_X1 NOT_776( .ZN(n787gat), .A(II2040) );
  INV_X1 NOT_777( .ZN(n775gat), .A(n777gat) );
  INV_X2 NOT_778( .ZN(II2044), .A(n775gat) );
  INV_X2 NOT_779( .ZN(n788gat), .A(II2044) );
  INV_X2 NOT_780( .ZN(n657gat), .A(n659gat) );
  INV_X1 NOT_781( .ZN(II2049), .A(n657gat) );
  INV_X1 NOT_782( .ZN(n789gat), .A(II2049) );
  INV_X1 NOT_783( .ZN(n35gat), .A(n779gat) );
  INV_X1 NOT_784( .ZN(II2056), .A(n35gat) );
  INV_X1 NOT_785( .ZN(n125gat), .A(II2056) );
  INV_X1 NOT_786( .ZN(n558gat), .A(n1725gat) );
  INV_X1 NOT_787( .ZN(n559gat), .A(n561gat) );
  INV_X1 NOT_788( .ZN(n371gat), .A(n1725gat) );
  INV_X1 NOT_789( .ZN(II2084), .A(n366gat) );
  INV_X1 NOT_790( .ZN(n365gat), .A(II2084) );
  INV_X1 NOT_791( .ZN(II2088), .A(n561gat) );
  INV_X1 NOT_792( .ZN(n560gat), .A(II2088) );
  INV_X1 NOT_793( .ZN(n364gat), .A(n366gat) );
  INV_X1 NOT_794( .ZN(II2094), .A(n2876gat) );
  INV_X1 NOT_795( .ZN(n126gat), .A(II2094) );
  INV_X1 NOT_796( .ZN(n663gat), .A(n1725gat) );
  INV_X1 NOT_797( .ZN(II2109), .A(n322gat) );
  INV_X1 NOT_798( .ZN(n321gat), .A(II2109) );
  INV_X1 NOT_799( .ZN(II2112), .A(n321gat) );
  INV_X1 NOT_800( .ZN(n226gat), .A(II2112) );
  INV_X1 NOT_801( .ZN(n370gat), .A(n1725gat) );
  INV_X1 NOT_802( .ZN(II2127), .A(n318gat) );
  INV_X1 NOT_803( .ZN(n317gat), .A(II2127) );
  INV_X1 NOT_804( .ZN(II2130), .A(n317gat) );
  INV_X1 NOT_805( .ZN(n227gat), .A(II2130) );
  INV_X1 NOT_806( .ZN(n369gat), .A(n1725gat) );
  INV_X1 NOT_807( .ZN(II2145), .A(n314gat) );
  INV_X1 NOT_808( .ZN(n313gat), .A(II2145) );
  INV_X1 NOT_809( .ZN(II2148), .A(n313gat) );
  INV_X1 NOT_810( .ZN(n228gat), .A(II2148) );
  INV_X1 NOT_811( .ZN(n316gat), .A(n318gat) );
  INV_X1 NOT_812( .ZN(II2153), .A(n316gat) );
  INV_X1 NOT_813( .ZN(n229gat), .A(II2153) );
  INV_X1 NOT_814( .ZN(n312gat), .A(n314gat) );
  INV_X1 NOT_815( .ZN(II2157), .A(n312gat) );
  INV_X1 NOT_816( .ZN(n230gat), .A(II2157) );
  INV_X1 NOT_817( .ZN(n320gat), .A(n322gat) );
  INV_X1 NOT_818( .ZN(II2162), .A(n320gat) );
  INV_X1 NOT_819( .ZN(n231gat), .A(II2162) );
  INV_X1 NOT_820( .ZN(n34gat), .A(n221gat) );
  INV_X1 NOT_821( .ZN(II2169), .A(n34gat) );
  INV_X1 NOT_822( .ZN(n127gat), .A(II2169) );
  INV_X1 NOT_823( .ZN(n133gat), .A(n2876gat) );
  INV_X1 NOT_824( .ZN(II2174), .A(n133gat) );
  INV_X1 NOT_825( .ZN(n128gat), .A(II2174) );
  INV_X1 NOT_826( .ZN(II2177), .A(n221gat) );
  INV_X1 NOT_827( .ZN(n129gat), .A(II2177) );
  INV_X1 NOT_828( .ZN(II2181), .A(n779gat) );
  INV_X1 NOT_829( .ZN(n130gat), .A(II2181) );
  INV_X1 NOT_830( .ZN(n665gat), .A(n667gat) );
  INV_X1 NOT_831( .ZN(n1601gat), .A(n120gat) );
  INV_X1 NOT_832( .ZN(n2597gat), .A(n2599gat) );
  INV_X1 NOT_833( .ZN(n2595gat), .A(n2594gat) );
  INV_X1 NOT_834( .ZN(n2586gat), .A(n2588gat) );
  INV_X1 NOT_835( .ZN(II2213), .A(n2342gat) );
  INV_X1 NOT_836( .ZN(n2573gat), .A(II2213) );
  INV_X1 NOT_837( .ZN(n2638gat), .A(n2640gat) );
  INV_X4 NOT_838( .ZN(II2225), .A(n2638gat) );
  INV_X4 NOT_839( .ZN(n2574gat), .A(II2225) );
  INV_X4 NOT_840( .ZN(II2228), .A(n2561gat) );
  INV_X1 NOT_841( .ZN(n2575gat), .A(II2228) );
  INV_X1 NOT_842( .ZN(II2232), .A(n2640gat) );
  INV_X1 NOT_843( .ZN(n2639gat), .A(II2232) );
  INV_X1 NOT_844( .ZN(II2235), .A(n2639gat) );
  INV_X1 NOT_845( .ZN(n2576gat), .A(II2235) );
  INV_X1 NOT_846( .ZN(II2238), .A(n2560gat) );
  INV_X1 NOT_847( .ZN(n2577gat), .A(II2238) );
  INV_X1 NOT_848( .ZN(II2242), .A(n2341gat) );
  INV_X1 NOT_849( .ZN(n2578gat), .A(II2242) );
  INV_X1 NOT_850( .ZN(II2248), .A(n2568gat) );
  INV_X1 NOT_851( .ZN(n2582gat), .A(II2248) );
  INV_X1 NOT_852( .ZN(II2251), .A(n2207gat) );
  INV_X1 NOT_853( .ZN(n2206gat), .A(II2251) );
  INV_X1 NOT_854( .ZN(II2254), .A(n2206gat) );
  INV_X1 NOT_855( .ZN(n2414gat), .A(II2254) );
  INV_X1 NOT_856( .ZN(II2257), .A(n2398gat) );
  INV_X1 NOT_857( .ZN(n2415gat), .A(II2257) );
  INV_X1 NOT_858( .ZN(II2260), .A(n2203gat) );
  INV_X1 NOT_859( .ZN(n2202gat), .A(II2260) );
  INV_X1 NOT_860( .ZN(II2263), .A(n2202gat) );
  INV_X1 NOT_861( .ZN(n2416gat), .A(II2263) );
  INV_X1 NOT_862( .ZN(n2397gat), .A(n2399gat) );
  INV_X1 NOT_863( .ZN(II2268), .A(n2397gat) );
  INV_X1 NOT_864( .ZN(n2417gat), .A(II2268) );
  INV_X1 NOT_865( .ZN(II2271), .A(n2201gat) );
  INV_X1 NOT_866( .ZN(n2418gat), .A(II2271) );
  INV_X1 NOT_867( .ZN(II2275), .A(n2205gat) );
  INV_X1 NOT_868( .ZN(n2419gat), .A(II2275) );
  INV_X1 NOT_869( .ZN(II2281), .A(n2409gat) );
  INV_X1 NOT_870( .ZN(n2585gat), .A(II2281) );
  INV_X1 NOT_871( .ZN(n2656gat), .A(n2658gat) );
  INV_X1 NOT_872( .ZN(n2493gat), .A(n2495gat) );
  INV_X1 NOT_873( .ZN(n2388gat), .A(n2390gat) );
  INV_X1 NOT_874( .ZN(II2316), .A(n2390gat) );
  INV_X1 NOT_875( .ZN(n2389gat), .A(II2316) );
  INV_X1 NOT_876( .ZN(II2319), .A(n2495gat) );
  INV_X1 NOT_877( .ZN(n2494gat), .A(II2319) );
  INV_X1 NOT_878( .ZN(II2324), .A(n3014gat) );
  INV_X1 NOT_879( .ZN(n2649gat), .A(II2324) );
  INV_X1 NOT_880( .ZN(n2268gat), .A(n2270gat) );
  INV_X1 NOT_881( .ZN(II2344), .A(n2339gat) );
  INV_X1 NOT_882( .ZN(n2338gat), .A(II2344) );
  INV_X1 NOT_883( .ZN(n2337gat), .A(n2339gat) );
  INV_X1 NOT_884( .ZN(II2349), .A(n2270gat) );
  INV_X1 NOT_885( .ZN(n2269gat), .A(II2349) );
  INV_X1 NOT_886( .ZN(II2354), .A(n2880gat) );
  INV_X8 NOT_887( .ZN(n2652gat), .A(II2354) );
  INV_X8 NOT_888( .ZN(n2500gat), .A(n2502gat) );
  INV_X1 NOT_889( .ZN(n2620gat), .A(n2622gat) );
  INV_X1 NOT_890( .ZN(n2612gat), .A(n2620gat) );
  INV_X1 NOT_891( .ZN(II2372), .A(n2612gat) );
  INV_X1 NOT_892( .ZN(n2606gat), .A(II2372) );
  INV_X1 NOT_893( .ZN(n2532gat), .A(n2625gat) );
  INV_X1 NOT_894( .ZN(II2376), .A(n2532gat) );
  INV_X1 NOT_895( .ZN(n2607gat), .A(II2376) );
  INV_X1 NOT_896( .ZN(n2540gat), .A(n2488gat) );
  INV_X1 NOT_897( .ZN(II2380), .A(n2540gat) );
  INV_X1 NOT_898( .ZN(n2608gat), .A(II2380) );
  INV_X1 NOT_899( .ZN(n2536gat), .A(n2624gat) );
  INV_X1 NOT_900( .ZN(II2385), .A(n2536gat) );
  INV_X1 NOT_901( .ZN(n2609gat), .A(II2385) );
  INV_X1 NOT_902( .ZN(n2487gat), .A(n2489gat) );
  INV_X1 NOT_903( .ZN(II2389), .A(n2487gat) );
  INV_X1 NOT_904( .ZN(n2610gat), .A(II2389) );
  INV_X1 NOT_905( .ZN(n2557gat), .A(n2621gat) );
  INV_X1 NOT_906( .ZN(II2394), .A(n2557gat) );
  INV_X1 NOT_907( .ZN(n2611gat), .A(II2394) );
  INV_X1 NOT_908( .ZN(II2400), .A(n2601gat) );
  INV_X1 NOT_909( .ZN(n2616gat), .A(II2400) );
  INV_X1 NOT_910( .ZN(II2403), .A(n2629gat) );
  INV_X1 NOT_911( .ZN(n2550gat), .A(II2403) );
  INV_X1 NOT_912( .ZN(II2414), .A(n2634gat) );
  INV_X1 NOT_913( .ZN(n2633gat), .A(II2414) );
  INV_X1 NOT_914( .ZN(II2417), .A(n2633gat) );
  INV_X1 NOT_915( .ZN(n2551gat), .A(II2417) );
  INV_X1 NOT_916( .ZN(II2420), .A(n2542gat) );
  INV_X1 NOT_917( .ZN(n2552gat), .A(II2420) );
  INV_X1 NOT_918( .ZN(n2632gat), .A(n2634gat) );
  INV_X1 NOT_919( .ZN(II2425), .A(n2632gat) );
  INV_X1 NOT_920( .ZN(n2553gat), .A(II2425) );
  INV_X1 NOT_921( .ZN(II2428), .A(n2541gat) );
  INV_X1 NOT_922( .ZN(n2554gat), .A(II2428) );
  INV_X1 NOT_923( .ZN(n2628gat), .A(n2630gat) );
  INV_X1 NOT_924( .ZN(II2433), .A(n2628gat) );
  INV_X1 NOT_925( .ZN(n2555gat), .A(II2433) );
  INV_X1 NOT_926( .ZN(II2439), .A(n2545gat) );
  INV_X1 NOT_927( .ZN(n2619gat), .A(II2439) );
  INV_X1 NOT_928( .ZN(n2504gat), .A(n2506gat) );
  INV_X1 NOT_929( .ZN(n2660gat), .A(n2655gat) );
  INV_X1 NOT_930( .ZN(n1528gat), .A(n2293gat) );
  INV_X1 NOT_931( .ZN(n1523gat), .A(n2219gat) );
  INV_X1 NOT_932( .ZN(n1592gat), .A(n1529gat) );
  INV_X1 NOT_933( .ZN(n2666gat), .A(n1704gat) );
  INV_X1 NOT_934( .ZN(n2422gat), .A(n3013gat) );
  INV_X1 NOT_935( .ZN(n2290gat), .A(n2202gat) );
  INV_X1 NOT_936( .ZN(n2081gat), .A(n2218gat) );
  INV_X1 NOT_937( .ZN(n2285gat), .A(n2397gat) );
  INV_X1 NOT_938( .ZN(n2359gat), .A(n2358gat) );
  INV_X1 NOT_939( .ZN(n1414gat), .A(n1415gat) );
  INV_X1 NOT_940( .ZN(n566gat), .A(n364gat) );
  INV_X1 NOT_941( .ZN(n1480gat), .A(n2292gat) );
  INV_X1 NOT_942( .ZN(n1301gat), .A(n1416gat) );
  INV_X16 NOT_943( .ZN(n1150gat), .A(n312gat) );
  INV_X16 NOT_944( .ZN(n873gat), .A(n316gat) );
  INV_X1 NOT_945( .ZN(n2011gat), .A(n2306gat) );
  INV_X1 NOT_946( .ZN(n1478gat), .A(n1481gat) );
  INV_X1 NOT_947( .ZN(n875gat), .A(n559gat) );
  INV_X1 NOT_948( .ZN(n1410gat), .A(n2357gat) );
  INV_X1 NOT_949( .ZN(n876gat), .A(n1347gat) );
  INV_X1 NOT_950( .ZN(n1160gat), .A(n1484gat) );
  INV_X1 NOT_951( .ZN(n1084gat), .A(n657gat) );
  INV_X1 NOT_952( .ZN(n983gat), .A(n320gat) );
  INV_X1 NOT_953( .ZN(n1482gat), .A(n2363gat) );
  INV_X1 NOT_954( .ZN(n1157gat), .A(n1483gat) );
  INV_X1 NOT_955( .ZN(n985gat), .A(n775gat) );
  INV_X1 NOT_956( .ZN(n1530gat), .A(n2364gat) );
  INV_X1 NOT_957( .ZN(n1307gat), .A(n1308gat) );
  INV_X1 NOT_958( .ZN(n1085gat), .A(n551gat) );
  INV_X1 NOT_959( .ZN(n1479gat), .A(n2291gat) );
  INV_X1 NOT_960( .ZN(n1348gat), .A(n1349gat) );
  INV_X1 NOT_961( .ZN(n2217gat), .A(n2206gat) );
  INV_X1 NOT_962( .ZN(n1591gat), .A(n2223gat) );
  INV_X1 NOT_963( .ZN(n1437gat), .A(n1438gat) );
  INV_X1 NOT_964( .ZN(n1832gat), .A(n1834gat) );
  INV_X1 NOT_965( .ZN(n1765gat), .A(n1767gat) );
  INV_X1 NOT_966( .ZN(n1878gat), .A(n1880gat) );
  INV_X1 NOT_967( .ZN(n1442gat), .A(n1831gat) );
  INV_X1 NOT_968( .ZN(n1444gat), .A(n1442gat) );
  INV_X1 NOT_969( .ZN(n1378gat), .A(n2975gat) );
  INV_X1 NOT_970( .ZN(n1322gat), .A(n2974gat) );
  INV_X1 NOT_971( .ZN(n1439gat), .A(n1486gat) );
  INV_X1 NOT_972( .ZN(n1370gat), .A(n1426gat) );
  INV_X1 NOT_973( .ZN(n1369gat), .A(n2966gat) );
  INV_X1 NOT_974( .ZN(n1366gat), .A(n1365gat) );
  INV_X1 NOT_975( .ZN(n1374gat), .A(n2979gat) );
  INV_X1 NOT_976( .ZN(n2162gat), .A(n2220gat) );
  INV_X1 NOT_977( .ZN(n1450gat), .A(n1423gat) );
  INV_X1 NOT_978( .ZN(n1427gat), .A(n1608gat) );
  INV_X1 NOT_979( .ZN(n1603gat), .A(n1831gat) );
  INV_X1 NOT_980( .ZN(n2082gat), .A(n2084gat) );
  INV_X1 NOT_981( .ZN(n1449gat), .A(n1494gat) );
  INV_X1 NOT_982( .ZN(n1590gat), .A(n1603gat) );
  INV_X1 NOT_983( .ZN(n1248gat), .A(n2954gat) );
  INV_X1 NOT_984( .ZN(n1418gat), .A(n1417gat) );
  INV_X1 NOT_985( .ZN(n1306gat), .A(n2964gat) );
  INV_X1 NOT_986( .ZN(n1353gat), .A(n1419gat) );
  INV_X1 NOT_987( .ZN(n1247gat), .A(n2958gat) );
  INV_X1 NOT_988( .ZN(n1355gat), .A(n1422gat) );
  INV_X1 NOT_989( .ZN(n1300gat), .A(n2963gat) );
  INV_X1 NOT_990( .ZN(n1487gat), .A(n1485gat) );
  INV_X1 NOT_991( .ZN(n1164gat), .A(n2953gat) );
  INV_X1 NOT_992( .ZN(n1356gat), .A(n1354gat) );
  INV_X1 NOT_993( .ZN(n1436gat), .A(n1435gat) );
  INV_X1 NOT_994( .ZN(n1106gat), .A(n2949gat) );
  INV_X1 NOT_995( .ZN(n1425gat), .A(n1421gat) );
  INV_X1 NOT_996( .ZN(n1105gat), .A(n2934gat) );
  INV_X1 NOT_997( .ZN(n1424gat), .A(n1420gat) );
  INV_X1 NOT_998( .ZN(n1309gat), .A(n2959gat) );
  INV_X1 NOT_999( .ZN(II2672), .A(n2143gat) );
  INV_X1 NOT_1000( .ZN(n2142gat), .A(II2672) );
  INV_X1 NOT_1001( .ZN(n1788gat), .A(n2142gat) );
  INV_X1 NOT_1002( .ZN(II2684), .A(n2061gat) );
  INV_X32 NOT_1003( .ZN(n2060gat), .A(II2684) );
  INV_X1 NOT_1004( .ZN(n1786gat), .A(n2060gat) );
  INV_X1 NOT_1005( .ZN(II2696), .A(n2139gat) );
  INV_X1 NOT_1006( .ZN(n2138gat), .A(II2696) );
  INV_X1 NOT_1007( .ZN(n1839gat), .A(n2138gat) );
  INV_X1 NOT_1008( .ZN(n1897gat), .A(n1899gat) );
  INV_X1 NOT_1009( .ZN(n1884gat), .A(n1897gat) );
  INV_X1 NOT_1010( .ZN(n1848gat), .A(n1850gat) );
  INV_X1 NOT_1011( .ZN(n1783gat), .A(n1848gat) );
  INV_X1 NOT_1012( .ZN(n1548gat), .A(II2721) );
  INV_X16 NOT_1013( .ZN(n1719gat), .A(n1548gat) );
  INV_X1 NOT_1014( .ZN(n2137gat), .A(n2139gat) );
  INV_X1 NOT_1015( .ZN(n1633gat), .A(n2137gat) );
  INV_X1 NOT_1016( .ZN(n2059gat), .A(n2061gat) );
  INV_X1 NOT_1017( .ZN(n1785gat), .A(n2059gat) );
  INV_X1 NOT_1018( .ZN(II2731), .A(n1850gat) );
  INV_X1 NOT_1019( .ZN(n1849gat), .A(II2731) );
  INV_X1 NOT_1020( .ZN(n1784gat), .A(n1849gat) );
  INV_X1 NOT_1021( .ZN(n1716gat), .A(II2736) );
  INV_X1 NOT_1022( .ZN(n1635gat), .A(n1716gat) );
  INV_X1 NOT_1023( .ZN(n2401gat), .A(n2403gat) );
  INV_X1 NOT_1024( .ZN(n1989gat), .A(n2401gat) );
  INV_X1 NOT_1025( .ZN(n2392gat), .A(n2394gat) );
  INV_X1 NOT_1026( .ZN(n1918gat), .A(n2392gat) );
  INV_X1 NOT_1027( .ZN(II2771), .A(n2440gat) );
  INV_X1 NOT_1028( .ZN(n2439gat), .A(II2771) );
  INV_X1 NOT_1029( .ZN(n1986gat), .A(n2439gat) );
  INV_X1 NOT_1030( .ZN(n1866gat), .A(n1865gat) );
  INV_X1 NOT_1031( .ZN(II2785), .A(n2407gat) );
  INV_X1 NOT_1032( .ZN(n2406gat), .A(II2785) );
  INV_X1 NOT_1033( .ZN(n2216gat), .A(n2406gat) );
  INV_X1 NOT_1034( .ZN(n2345gat), .A(n2347gat) );
  INV_X1 NOT_1035( .ZN(n1988gat), .A(n2345gat) );
  INV_X1 NOT_1036( .ZN(n1735gat), .A(n1861gat) );
  INV_X1 NOT_1037( .ZN(n1387gat), .A(n1389gat) );
  INV_X1 NOT_1038( .ZN(n1694gat), .A(II2813) );
  INV_X1 NOT_1039( .ZN(n1777gat), .A(n1694gat) );
  INV_X1 NOT_1040( .ZN(n1781gat), .A(n1780gat) );
  INV_X1 NOT_1041( .ZN(n2019gat), .A(n2021gat) );
  INV_X1 NOT_1042( .ZN(n1549gat), .A(II2832) );
  INV_X1 NOT_1043( .ZN(n1551gat), .A(n1549gat) );
  INV_X1 NOT_1044( .ZN(II2837), .A(n2347gat) );
  INV_X1 NOT_1045( .ZN(n2346gat), .A(II2837) );
  INV_X1 NOT_1046( .ZN(n2152gat), .A(n2346gat) );
  INV_X1 NOT_1047( .ZN(n2405gat), .A(n2407gat) );
  INV_X1 NOT_1048( .ZN(n2351gat), .A(n2405gat) );
  INV_X1 NOT_1049( .ZN(II2843), .A(n2403gat) );
  INV_X1 NOT_1050( .ZN(n2402gat), .A(II2843) );
  INV_X1 NOT_1051( .ZN(n2212gat), .A(n2402gat) );
  INV_X1 NOT_1052( .ZN(II2847), .A(n2394gat) );
  INV_X1 NOT_1053( .ZN(n2393gat), .A(II2847) );
  INV_X2 NOT_1054( .ZN(n1991gat), .A(n2393gat) );
  INV_X2 NOT_1055( .ZN(n1665gat), .A(n1666gat) );
  INV_X2 NOT_1056( .ZN(n1517gat), .A(n1578gat) );
  INV_X1 NOT_1057( .ZN(n1392gat), .A(n1394gat) );
  INV_X1 NOT_1058( .ZN(II2873), .A(n1496gat) );
  INV_X1 NOT_1059( .ZN(n1495gat), .A(II2873) );
  INV_X1 NOT_1060( .ZN(n1685gat), .A(n1604gat) );
  INV_X1 NOT_1061( .ZN(II2885), .A(n2091gat) );
  INV_X1 NOT_1062( .ZN(n2090gat), .A(II2885) );
  INV_X1 NOT_1063( .ZN(n1550gat), .A(II2890) );
  INV_X1 NOT_1064( .ZN(n1552gat), .A(n1550gat) );
  INV_X1 NOT_1065( .ZN(n1330gat), .A(n1332gat) );
  INV_X1 NOT_1066( .ZN(n1738gat), .A(n1740gat) );
  INV_X1 NOT_1067( .ZN(II2915), .A(n1740gat) );
  INV_X1 NOT_1068( .ZN(n1739gat), .A(II2915) );
  INV_X1 NOT_1069( .ZN(n1925gat), .A(n1920gat) );
  INV_X1 NOT_1070( .ZN(n1917gat), .A(n1921gat) );
  INV_X1 NOT_1071( .ZN(n2141gat), .A(n2143gat) );
  INV_X1 NOT_1072( .ZN(n1787gat), .A(n2141gat) );
  INV_X1 NOT_1073( .ZN(n1717gat), .A(II2926) );
  INV_X1 NOT_1074( .ZN(n1859gat), .A(n1717gat) );
  INV_X1 NOT_1075( .ZN(n1922gat), .A(n1798gat) );
  INV_X1 NOT_1076( .ZN(n1713gat), .A(II2935) );
  INV_X1 NOT_1077( .ZN(n1743gat), .A(n1713gat) );
  INV_X1 NOT_1078( .ZN(n1923gat), .A(n1864gat) );
  INV_X1 NOT_1079( .ZN(n1945gat), .A(n1690gat) );
  INV_X1 NOT_1080( .ZN(II2953), .A(n2179gat) );
  INV_X1 NOT_1081( .ZN(n2178gat), .A(II2953) );
  INV_X1 NOT_1082( .ZN(n1661gat), .A(n1660gat) );
  INV_X1 NOT_1083( .ZN(n1572gat), .A(n1576gat) );
  INV_X1 NOT_1084( .ZN(n2438gat), .A(n2440gat) );
  INV_X1 NOT_1085( .ZN(n2283gat), .A(n2438gat) );
  INV_X1 NOT_1086( .ZN(n1520gat), .A(n1582gat) );
  INV_X1 NOT_1087( .ZN(n1580gat), .A(n1577gat) );
  INV_X1 NOT_1088( .ZN(n1990gat), .A(n2988gat) );
  INV_X1 NOT_1089( .ZN(II2978), .A(n2190gat) );
  INV_X1 NOT_1090( .ZN(n2189gat), .A(II2978) );
  INV_X1 NOT_1091( .ZN(II2989), .A(n2135gat) );
  INV_X1 NOT_1092( .ZN(n2134gat), .A(II2989) );
  INV_X1 NOT_1093( .ZN(II3000), .A(n2262gat) );
  INV_X1 NOT_1094( .ZN(n2261gat), .A(II3000) );
  INV_X1 NOT_1095( .ZN(n2128gat), .A(n2129gat) );
  INV_X1 NOT_1096( .ZN(n1836gat), .A(n1695gat) );
  INV_X1 NOT_1097( .ZN(II3016), .A(n2182gat) );
  INV_X1 NOT_1098( .ZN(n2181gat), .A(II3016) );
  INV_X1 NOT_1099( .ZN(n1431gat), .A(n1433gat) );
  INV_X1 NOT_1100( .ZN(n1314gat), .A(n1316gat) );
  INV_X1 NOT_1101( .ZN(n1361gat), .A(n1363gat) );
  INV_X1 NOT_1102( .ZN(II3056), .A(n1312gat) );
  INV_X1 NOT_1103( .ZN(n1311gat), .A(II3056) );
  INV_X1 NOT_1104( .ZN(n1707gat), .A(n1626gat) );
  INV_X1 NOT_1105( .ZN(n1773gat), .A(n1775gat) );
  INV_X1 NOT_1106( .ZN(n1659gat), .A(n2987gat) );
  INV_X1 NOT_1107( .ZN(n1515gat), .A(n1521gat) );
  INV_X1 NOT_1108( .ZN(n1736gat), .A(n1737gat) );
  INV_X1 NOT_1109( .ZN(n1658gat), .A(n2216gat) );
  INV_X1 NOT_1110( .ZN(n1724gat), .A(n1732gat) );
  INV_X1 NOT_1111( .ZN(n1662gat), .A(n1663gat) );
  INV_X4 NOT_1112( .ZN(n1656gat), .A(n1655gat) );
  INV_X4 NOT_1113( .ZN(n1670gat), .A(n1667gat) );
  INV_X4 NOT_1114( .ZN(n1569gat), .A(n1570gat) );
  INV_X1 NOT_1115( .ZN(n1568gat), .A(n1575gat) );
  INV_X1 NOT_1116( .ZN(n1727gat), .A(n1728gat) );
  INV_X1 NOT_1117( .ZN(n1797gat), .A(n1801gat) );
  INV_X1 NOT_1118( .ZN(n1730gat), .A(n1731gat) );
  INV_X1 NOT_1119( .ZN(n1561gat), .A(n1571gat) );
  INV_X1 NOT_1120( .ZN(n1668gat), .A(n1734gat) );
  INV_X1 NOT_1121( .ZN(n1742gat), .A(n2216gat) );
  INV_X1 NOT_1122( .ZN(n1671gat), .A(n1669gat) );
  INV_X1 NOT_1123( .ZN(n1652gat), .A(n1657gat) );
  INV_X1 NOT_1124( .ZN(n1648gat), .A(n1729gat) );
  INV_X1 NOT_1125( .ZN(n1790gat), .A(n1726gat) );
  INV_X1 NOT_1126( .ZN(n2004gat), .A(n1929gat) );
  INV_X1 NOT_1127( .ZN(n1869gat), .A(n1871gat) );
  INV_X1 NOT_1128( .ZN(II3143), .A(n2592gat) );
  INV_X1 NOT_1129( .ZN(n2591gat), .A(II3143) );
  INV_X1 NOT_1130( .ZN(n1584gat), .A(n2989gat) );
  INV_X1 NOT_1131( .ZN(n1714gat), .A(II3149) );
  INV_X1 NOT_1132( .ZN(n1718gat), .A(n1714gat) );
  INV_X1 NOT_1133( .ZN(II3163), .A(n1508gat) );
  INV_X1 NOT_1134( .ZN(n1507gat), .A(II3163) );
  INV_X1 NOT_1135( .ZN(n1396gat), .A(n1401gat) );
  INV_X1 NOT_1136( .ZN(II3168), .A(n1394gat) );
  INV_X1 NOT_1137( .ZN(n1393gat), .A(II3168) );
  INV_X1 NOT_1138( .ZN(n1409gat), .A(n1476gat) );
  INV_X1 NOT_1139( .ZN(II3174), .A(n1899gat) );
  INV_X1 NOT_1140( .ZN(n1898gat), .A(II3174) );
  INV_X1 NOT_1141( .ZN(n1838gat), .A(n1898gat) );
  INV_X1 NOT_1142( .ZN(n1712gat), .A(II3179) );
  INV_X1 NOT_1143( .ZN(II3191), .A(n1678gat) );
  INV_X1 NOT_1144( .ZN(n1677gat), .A(II3191) );
  INV_X1 NOT_1145( .ZN(n2000gat), .A(n1412gat) );
  INV_X1 NOT_1146( .ZN(n2001gat), .A(n1412gat) );
  INV_X1 NOT_1147( .ZN(n1999gat), .A(n2001gat) );
  INV_X1 NOT_1148( .ZN(n2307gat), .A(n2309gat) );
  INV_X1 NOT_1149( .ZN(II3211), .A(n2663gat) );
  INV_X1 NOT_1150( .ZN(n3018gat), .A(II3211) );
  INV_X1 NOT_1151( .ZN(n2448gat), .A(n2450gat) );
  INV_X1 NOT_1152( .ZN(n2661gat), .A(n2662gat) );
  INV_X1 NOT_1153( .ZN(n2444gat), .A(n2446gat) );
  INV_X1 NOT_1154( .ZN(II3235), .A(n2238gat) );
  INV_X1 NOT_1155( .ZN(n3019gat), .A(II3235) );
  INV_X1 NOT_1156( .ZN(n1310gat), .A(n1312gat) );
  INV_X1 NOT_1157( .ZN(n199gat), .A(n87gat) );
  INV_X1 NOT_1158( .ZN(n195gat), .A(n184gat) );
  INV_X1 NOT_1159( .ZN(n827gat), .A(n204gat) );
  INV_X1 NOT_1160( .ZN(n2093gat), .A(n2095gat) );
  INV_X1 NOT_1161( .ZN(n2174gat), .A(n2176gat) );
  INV_X1 NOT_1162( .ZN(II3273), .A(n2169gat) );
  INV_X1 NOT_1163( .ZN(n2168gat), .A(II3273) );
  INV_X1 NOT_1164( .ZN(n2452gat), .A(n2454gat) );
  INV_X1 NOT_1165( .ZN(n1691gat), .A(n2452gat) );
  INV_X1 NOT_1166( .ZN(II3287), .A(n1691gat) );
  INV_X1 NOT_1167( .ZN(n3020gat), .A(II3287) );
  INV_X1 NOT_1168( .ZN(II3290), .A(n1691gat) );
  INV_X1 NOT_1169( .ZN(n3021gat), .A(II3290) );
  INV_X2 NOT_1170( .ZN(II3293), .A(n1691gat) );
  INV_X2 NOT_1171( .ZN(n3022gat), .A(II3293) );
  INV_X1 NOT_1172( .ZN(n1699gat), .A(n2452gat) );
  INV_X1 NOT_1173( .ZN(II3297), .A(n1699gat) );
  INV_X1 NOT_1174( .ZN(n3023gat), .A(II3297) );
  INV_X1 NOT_1175( .ZN(II3300), .A(n1699gat) );
  INV_X1 NOT_1176( .ZN(n3024gat), .A(II3300) );
  INV_X1 NOT_1177( .ZN(II3303), .A(n1691gat) );
  INV_X1 NOT_1178( .ZN(n3025gat), .A(II3303) );
  INV_X1 NOT_1179( .ZN(II3306), .A(n1699gat) );
  INV_X1 NOT_1180( .ZN(n3026gat), .A(II3306) );
  INV_X1 NOT_1181( .ZN(II3309), .A(n1699gat) );
  INV_X1 NOT_1182( .ZN(n3027gat), .A(II3309) );
  INV_X1 NOT_1183( .ZN(II3312), .A(n1699gat) );
  INV_X1 NOT_1184( .ZN(n3028gat), .A(II3312) );
  INV_X1 NOT_1185( .ZN(II3315), .A(n1869gat) );
  INV_X1 NOT_1186( .ZN(n3029gat), .A(II3315) );
  INV_X1 NOT_1187( .ZN(II3318), .A(n1869gat) );
  INV_X1 NOT_1188( .ZN(n3030gat), .A(II3318) );
  INV_X1 NOT_1189( .ZN(n2260gat), .A(n2262gat) );
  INV_X1 NOT_1190( .ZN(n2257gat), .A(n2189gat) );
  INV_X1 NOT_1191( .ZN(n2188gat), .A(n2190gat) );
  INV_X1 NOT_1192( .ZN(n2187gat), .A(n3004gat) );
  INV_X1 NOT_1193( .ZN(II3336), .A(n2040gat) );
  INV_X1 NOT_1194( .ZN(n2039gat), .A(II3336) );
  INV_X1 NOT_1195( .ZN(II3339), .A(n1775gat) );
  INV_X1 NOT_1196( .ZN(n1774gat), .A(II3339) );
  INV_X1 NOT_1197( .ZN(II3342), .A(n1316gat) );
  INV_X1 NOT_1198( .ZN(n1315gat), .A(II3342) );
  INV_X1 NOT_1199( .ZN(n2042gat), .A(n2044gat) );
  INV_X1 NOT_1200( .ZN(n2035gat), .A(n2037gat) );
  INV_X1 NOT_1201( .ZN(n2023gat), .A(n2025gat) );
  INV_X1 NOT_1202( .ZN(n2097gat), .A(n2099gat) );
  INV_X1 NOT_1203( .ZN(n1855gat), .A(n2014gat) );
  INV_X1 NOT_1204( .ZN(II3387), .A(n2194gat) );
  INV_X1 NOT_1205( .ZN(n3031gat), .A(II3387) );
  INV_X1 NOT_1206( .ZN(II3390), .A(n2261gat) );
  INV_X1 NOT_1207( .ZN(n3032gat), .A(II3390) );
  INV_X1 NOT_1208( .ZN(n2256gat), .A(n3032gat) );
  INV_X1 NOT_1209( .ZN(II3394), .A(n2260gat) );
  INV_X1 NOT_1210( .ZN(n3033gat), .A(II3394) );
  INV_X1 NOT_1211( .ZN(n2251gat), .A(n3033gat) );
  INV_X1 NOT_1212( .ZN(n2184gat), .A(n3003gat) );
  INV_X1 NOT_1213( .ZN(II3401), .A(n2192gat) );
  INV_X1 NOT_1214( .ZN(n3034gat), .A(II3401) );
  INV_X1 NOT_1215( .ZN(n2133gat), .A(n2135gat) );
  INV_X1 NOT_1216( .ZN(n2131gat), .A(n2185gat) );
  INV_X1 NOT_1217( .ZN(n2049gat), .A(n3001gat) );
  INV_X1 NOT_1218( .ZN(II3412), .A(n2057gat) );
  INV_X1 NOT_1219( .ZN(n3035gat), .A(II3412) );
  INV_X1 NOT_1220( .ZN(n2253gat), .A(n2189gat) );
  INV_X1 NOT_1221( .ZN(n2252gat), .A(n2260gat) );
  INV_X1 NOT_1222( .ZN(n2248gat), .A(n3006gat) );
  INV_X1 NOT_1223( .ZN(n2264gat), .A(n2266gat) );
  INV_X2 NOT_1224( .ZN(II3429), .A(n2266gat) );
  INV_X2 NOT_1225( .ZN(n2265gat), .A(II3429) );
  INV_X1 NOT_1226( .ZN(n2492gat), .A(n2329gat) );
  INV_X1 NOT_1227( .ZN(II3436), .A(n2492gat) );
  INV_X1 NOT_1228( .ZN(n3036gat), .A(II3436) );
  INV_X1 NOT_1229( .ZN(n1709gat), .A(n1849gat) );
  INV_X1 NOT_1230( .ZN(n1845gat), .A(n2141gat) );
  INV_X1 NOT_1231( .ZN(n1891gat), .A(n2059gat) );
  INV_X1 NOT_1232( .ZN(n1963gat), .A(n2137gat) );
  INV_X1 NOT_1233( .ZN(n1886gat), .A(n1897gat) );
  INV_X1 NOT_1234( .ZN(n1968gat), .A(n1958gat) );
  INV_X1 NOT_1235( .ZN(n1629gat), .A(n1895gat) );
  INV_X1 NOT_1236( .ZN(n1631gat), .A(n1848gat) );
  INV_X1 NOT_1237( .ZN(n1711gat), .A(n2990gat) );
  INV_X1 NOT_1238( .ZN(n2200gat), .A(n2078gat) );
  INV_X1 NOT_1239( .ZN(n2437gat), .A(n2195gat) );
  INV_X1 NOT_1240( .ZN(II3457), .A(n2556gat) );
  INV_X1 NOT_1241( .ZN(n3037gat), .A(II3457) );
  INV_X1 NOT_1242( .ZN(n1956gat), .A(n1898gat) );
  INV_X1 NOT_1243( .ZN(II3461), .A(n1956gat) );
  INV_X1 NOT_1244( .ZN(n3038gat), .A(II3461) );
  INV_X1 NOT_1245( .ZN(n1954gat), .A(n3038gat) );
  INV_X1 NOT_1246( .ZN(II3465), .A(n1886gat) );
  INV_X1 NOT_1247( .ZN(n3039gat), .A(II3465) );
  INV_X1 NOT_1248( .ZN(n1888gat), .A(n3039gat) );
  INV_X1 NOT_1249( .ZN(n2048gat), .A(n2994gat) );
  INV_X1 NOT_1250( .ZN(II3472), .A(n2539gat) );
  INV_X1 NOT_1251( .ZN(n3040gat), .A(II3472) );
  INV_X1 NOT_1252( .ZN(n1969gat), .A(n2142gat) );
  INV_X1 NOT_1253( .ZN(n1893gat), .A(n2060gat) );
  INV_X1 NOT_1254( .ZN(n1892gat), .A(n2993gat) );
  INV_X1 NOT_1255( .ZN(II3483), .A(n2436gat) );
  INV_X1 NOT_1256( .ZN(n3041gat), .A(II3483) );
  INV_X1 NOT_1257( .ZN(n2056gat), .A(n2998gat) );
  INV_X1 NOT_1258( .ZN(II3491), .A(n2387gat) );
  INV_X1 NOT_1259( .ZN(n3042gat), .A(II3491) );
  INV_X1 NOT_1260( .ZN(II3494), .A(n1963gat) );
  INV_X1 NOT_1261( .ZN(n3043gat), .A(II3494) );
  INV_X1 NOT_1262( .ZN(n1960gat), .A(n3043gat) );
  INV_X1 NOT_1263( .ZN(n1887gat), .A(n2138gat) );
  INV_X1 NOT_1264( .ZN(n1961gat), .A(n2996gat) );
  INV_X1 NOT_1265( .ZN(II3504), .A(n2330gat) );
  INV_X1 NOT_1266( .ZN(n3044gat), .A(II3504) );
  INV_X1 NOT_1267( .ZN(n2199gat), .A(n2147gat) );
  INV_X1 NOT_1268( .ZN(II3509), .A(n2438gat) );
  INV_X1 NOT_1269( .ZN(n3045gat), .A(II3509) );
  INV_X1 NOT_1270( .ZN(n2332gat), .A(n3045gat) );
  INV_X1 NOT_1271( .ZN(II3513), .A(n2439gat) );
  INV_X1 NOT_1272( .ZN(n3046gat), .A(II3513) );
  INV_X1 NOT_1273( .ZN(n2259gat), .A(n3046gat) );
  INV_X1 NOT_1274( .ZN(n2328gat), .A(n3008gat) );
  INV_X1 NOT_1275( .ZN(II3520), .A(n2498gat) );
  INV_X1 NOT_1276( .ZN(n3047gat), .A(II3520) );
  INV_X2 NOT_1277( .ZN(n2151gat), .A(n2193gat) );
  INV_X2 NOT_1278( .ZN(n2209gat), .A(n3005gat) );
  INV_X1 NOT_1279( .ZN(II3530), .A(n2396gat) );
  INV_X1 NOT_1280( .ZN(n3048gat), .A(II3530) );
  INV_X1 NOT_1281( .ZN(n2052gat), .A(n2393gat) );
  INV_X1 NOT_1282( .ZN(n2058gat), .A(n2997gat) );
  INV_X1 NOT_1283( .ZN(II3539), .A(n2198gat) );
  INV_X1 NOT_1284( .ZN(n3049gat), .A(II3539) );
  INV_X1 NOT_1285( .ZN(n2349gat), .A(n2215gat) );
  INV_X1 NOT_1286( .ZN(n2281gat), .A(n3009gat) );
  INV_X1 NOT_1287( .ZN(II3549), .A(n2197gat) );
  INV_X1 NOT_1288( .ZN(n3050gat), .A(II3549) );
  INV_X1 NOT_1289( .ZN(n2146gat), .A(n3002gat) );
  INV_X1 NOT_1290( .ZN(II3558), .A(n2196gat) );
  INV_X1 NOT_1291( .ZN(n3051gat), .A(II3558) );
  INV_X1 NOT_1292( .ZN(n2031gat), .A(n2033gat) );
  INV_X1 NOT_1293( .ZN(n2108gat), .A(n2110gat) );
  INV_X1 NOT_1294( .ZN(II3587), .A(n2125gat) );
  INV_X1 NOT_1295( .ZN(n2124gat), .A(II3587) );
  INV_X1 NOT_1296( .ZN(n2123gat), .A(n2125gat) );
  INV_X1 NOT_1297( .ZN(n2119gat), .A(n2121gat) );
  INV_X1 NOT_1298( .ZN(n2115gat), .A(n2117gat) );
  INV_X1 NOT_1299( .ZN(II3610), .A(n1882gat) );
  INV_X1 NOT_1300( .ZN(n3052gat), .A(II3610) );
  INV_X1 NOT_1301( .ZN(II3621), .A(n1975gat) );
  INV_X1 NOT_1302( .ZN(n1974gat), .A(II3621) );
  INV_X1 NOT_1303( .ZN(n1955gat), .A(n1956gat) );
  INV_X1 NOT_1304( .ZN(n1970gat), .A(n1896gat) );
  INV_X1 NOT_1305( .ZN(n1973gat), .A(n1975gat) );
  INV_X1 NOT_1306( .ZN(n2558gat), .A(n2559gat) );
  INV_X1 NOT_1307( .ZN(II3635), .A(n2558gat) );
  INV_X1 NOT_1308( .ZN(n3053gat), .A(II3635) );
  INV_X1 NOT_1309( .ZN(II3646), .A(n2644gat) );
  INV_X1 NOT_1310( .ZN(n2643gat), .A(II3646) );
  INV_X1 NOT_1311( .ZN(n2333gat), .A(n2438gat) );
  INV_X1 NOT_1312( .ZN(n2564gat), .A(n2352gat) );
  INV_X1 NOT_1313( .ZN(n2642gat), .A(n2644gat) );
  INV_X1 NOT_1314( .ZN(n2636gat), .A(n2637gat) );
  INV_X1 NOT_1315( .ZN(II3660), .A(n2636gat) );
  INV_X1 NOT_1316( .ZN(n3054gat), .A(II3660) );
  INV_X1 NOT_1317( .ZN(n88gat), .A(n84gat) );
  INV_X1 NOT_1318( .ZN(n375gat), .A(n110gat) );
  INV_X1 NOT_1319( .ZN(II3677), .A(n156gat) );
  INV_X1 NOT_1320( .ZN(n155gat), .A(II3677) );
  INV_X1 NOT_1321( .ZN(n253gat), .A(n1702gat) );
  INV_X1 NOT_1322( .ZN(n150gat), .A(n152gat) );
  INV_X1 NOT_1323( .ZN(II3691), .A(n152gat) );
  INV_X1 NOT_1324( .ZN(n151gat), .A(II3691) );
  INV_X1 NOT_1325( .ZN(n243gat), .A(n1702gat) );
  INV_X1 NOT_1326( .ZN(n233gat), .A(n243gat) );
  INV_X1 NOT_1327( .ZN(n154gat), .A(n156gat) );
  INV_X1 NOT_1328( .ZN(n800gat), .A(n2874gat) );
  INV_X1 NOT_1329( .ZN(II3703), .A(n2917gat) );
  INV_X1 NOT_1330( .ZN(n3055gat), .A(II3703) );
  INV_X1 NOT_1331( .ZN(n235gat), .A(n2878gat) );
  INV_X1 NOT_1332( .ZN(II3713), .A(n2892gat) );
  INV_X1 NOT_1333( .ZN(n3056gat), .A(II3713) );
  INV_X4 NOT_1334( .ZN(n372gat), .A(n212gat) );
  INV_X4 NOT_1335( .ZN(n329gat), .A(n331gat) );
  INV_X1 NOT_1336( .ZN(II3736), .A(n388gat) );
  INV_X1 NOT_1337( .ZN(n387gat), .A(II3736) );
  INV_X1 NOT_1338( .ZN(n334gat), .A(n1700gat) );
  INV_X1 NOT_1339( .ZN(n386gat), .A(n388gat) );
  INV_X1 NOT_1340( .ZN(II3742), .A(n331gat) );
  INV_X1 NOT_1341( .ZN(n330gat), .A(II3742) );
  INV_X1 NOT_1342( .ZN(n1430gat), .A(n1700gat) );
  INV_X1 NOT_1343( .ZN(n1490gat), .A(n1430gat) );
  INV_X1 NOT_1344( .ZN(n452gat), .A(n2885gat) );
  INV_X1 NOT_1345( .ZN(II3754), .A(n2900gat) );
  INV_X1 NOT_1346( .ZN(n3057gat), .A(II3754) );
  INV_X1 NOT_1347( .ZN(n333gat), .A(n2883gat) );
  INV_X1 NOT_1348( .ZN(II3765), .A(n2929gat) );
  INV_X1 NOT_1349( .ZN(n3058gat), .A(II3765) );
  INV_X1 NOT_1350( .ZN(II3777), .A(n463gat) );
  INV_X1 NOT_1351( .ZN(n462gat), .A(II3777) );
  INV_X1 NOT_1352( .ZN(n325gat), .A(n327gat) );
  INV_X1 NOT_1353( .ZN(n457gat), .A(n2884gat) );
  INV_X1 NOT_1354( .ZN(n461gat), .A(n463gat) );
  INV_X1 NOT_1355( .ZN(n458gat), .A(n2902gat) );
  INV_X1 NOT_1356( .ZN(II3801), .A(n2925gat) );
  INV_X1 NOT_1357( .ZN(n3059gat), .A(II3801) );
  INV_X1 NOT_1358( .ZN(n144gat), .A(n247gat) );
  INV_X1 NOT_1359( .ZN(II3808), .A(n327gat) );
  INV_X1 NOT_1360( .ZN(n326gat), .A(II3808) );
  INV_X1 NOT_1361( .ZN(n878gat), .A(n2879gat) );
  INV_X1 NOT_1362( .ZN(II3817), .A(n2916gat) );
  INV_X1 NOT_1363( .ZN(n3060gat), .A(II3817) );
  INV_X1 NOT_1364( .ZN(n382gat), .A(n384gat) );
  INV_X1 NOT_1365( .ZN(II3831), .A(n384gat) );
  INV_X1 NOT_1366( .ZN(n383gat), .A(II3831) );
  INV_X1 NOT_1367( .ZN(n134gat), .A(n2875gat) );
  INV_X1 NOT_1368( .ZN(II3841), .A(n2899gat) );
  INV_X1 NOT_1369( .ZN(n3061gat), .A(II3841) );
  INV_X1 NOT_1370( .ZN(n254gat), .A(n256gat) );
  INV_X1 NOT_1371( .ZN(n252gat), .A(n2877gat) );
  INV_X1 NOT_1372( .ZN(n468gat), .A(n470gat) );
  INV_X1 NOT_1373( .ZN(II3867), .A(n470gat) );
  INV_X1 NOT_1374( .ZN(n469gat), .A(II3867) );
  INV_X1 NOT_1375( .ZN(n381gat), .A(n2893gat) );
  INV_X1 NOT_1376( .ZN(II3876), .A(n2926gat) );
  INV_X1 NOT_1377( .ZN(n3062gat), .A(II3876) );
  INV_X1 NOT_1378( .ZN(n241gat), .A(n140gat) );
  INV_X1 NOT_1379( .ZN(II3882), .A(n256gat) );
  INV_X1 NOT_1380( .ZN(n255gat), .A(II3882) );
  INV_X1 NOT_1381( .ZN(n802gat), .A(n2882gat) );
  INV_X1 NOT_1382( .ZN(II3891), .A(n2924gat) );
  INV_X1 NOT_1383( .ZN(n3063gat), .A(II3891) );
  INV_X1 NOT_1384( .ZN(n146gat), .A(n148gat) );
  INV_X1 NOT_1385( .ZN(II3904), .A(n148gat) );
  INV_X1 NOT_1386( .ZN(n147gat), .A(II3904) );
  INV_X1 NOT_1387( .ZN(n380gat), .A(n2881gat) );
  INV_X1 NOT_1388( .ZN(II3914), .A(n2923gat) );
  INV_X1 NOT_1389( .ZN(n3064gat), .A(II3914) );
  INV_X4 NOT_1390( .ZN(n69gat), .A(n68gat) );
  INV_X4 NOT_1391( .ZN(n1885gat), .A(n2048gat) );
  INV_X1 NOT_1392( .ZN(II3923), .A(n2710gat) );
  INV_X1 NOT_1393( .ZN(n2707gat), .A(II3923) );
  INV_X1 NOT_1394( .ZN(n16gat), .A(n564gat) );
  INV_X1 NOT_1395( .ZN(n295gat), .A(n357gat) );
  INV_X1 NOT_1396( .ZN(n11gat), .A(n12gat) );
  INV_X1 NOT_1397( .ZN(n1889gat), .A(n1961gat) );
  INV_X1 NOT_1398( .ZN(II3935), .A(n2704gat) );
  INV_X1 NOT_1399( .ZN(n2700gat), .A(II3935) );
  INV_X1 NOT_1400( .ZN(n2051gat), .A(n2056gat) );
  INV_X1 NOT_1401( .ZN(II3941), .A(n2684gat) );
  INV_X1 NOT_1402( .ZN(n2680gat), .A(II3941) );
  INV_X1 NOT_1403( .ZN(n1350gat), .A(n1831gat) );
  INV_X1 NOT_1404( .ZN(II3945), .A(n1350gat) );
  INV_X1 NOT_1405( .ZN(n2696gat), .A(II3945) );
  INV_X1 NOT_1406( .ZN(II3948), .A(n2696gat) );
  INV_X1 NOT_1407( .ZN(n2692gat), .A(II3948) );
  INV_X1 NOT_1408( .ZN(II3951), .A(n2448gat) );
  INV_X1 NOT_1409( .ZN(n2683gat), .A(II3951) );
  INV_X1 NOT_1410( .ZN(II3954), .A(n2683gat) );
  INV_X1 NOT_1411( .ZN(n2679gat), .A(II3954) );
  INV_X1 NOT_1412( .ZN(II3957), .A(n2450gat) );
  INV_X1 NOT_1413( .ZN(n2449gat), .A(II3957) );
  INV_X1 NOT_1414( .ZN(n1754gat), .A(n2449gat) );
  INV_X1 NOT_1415( .ZN(II3962), .A(n2830gat) );
  INV_X1 NOT_1416( .ZN(n2827gat), .A(II3962) );
  INV_X1 NOT_1417( .ZN(n2590gat), .A(n2592gat) );
  INV_X1 NOT_1418( .ZN(n2456gat), .A(n2458gat) );
  INV_X1 NOT_1419( .ZN(n2512gat), .A(n2514gat) );
  INV_X1 NOT_1420( .ZN(n1544gat), .A(n1625gat) );
  INV_X1 NOT_1421( .ZN(n1769gat), .A(n1771gat) );
  INV_X1 NOT_1422( .ZN(n1683gat), .A(n1756gat) );
  INV_X1 NOT_1423( .ZN(n2167gat), .A(n2169gat) );
  INV_X1 NOT_1424( .ZN(n2013gat), .A(II4000) );
  INV_X1 NOT_1425( .ZN(n1791gat), .A(n2013gat) );
  INV_X1 NOT_1426( .ZN(n2691gat), .A(n2695gat) );
  INV_X1 NOT_1427( .ZN(n1518gat), .A(n1694gat) );
  INV_X1 NOT_1428( .ZN(n2699gat), .A(n2703gat) );
  INV_X1 NOT_1429( .ZN(n2159gat), .A(n1412gat) );
  INV_X1 NOT_1430( .ZN(n2478gat), .A(n2579gat) );
  INV_X1 NOT_1431( .ZN(II4014), .A(n2744gat) );
  INV_X1 NOT_1432( .ZN(n2740gat), .A(II4014) );
  INV_X1 NOT_1433( .ZN(n2158gat), .A(n1412gat) );
  INV_X1 NOT_1434( .ZN(n2186gat), .A(n2613gat) );
  INV_X1 NOT_1435( .ZN(II4020), .A(n2800gat) );
  INV_X1 NOT_1436( .ZN(n2797gat), .A(II4020) );
  INV_X1 NOT_1437( .ZN(n2288gat), .A(II4024) );
  INV_X1 NOT_1438( .ZN(n1513gat), .A(n2288gat) );
  INV_X1 NOT_1439( .ZN(n2537gat), .A(n2538gat) );
  INV_X1 NOT_1440( .ZN(n2442gat), .A(n2483gat) );
  INV_X1 NOT_1441( .ZN(n1334gat), .A(n1336gat) );
  INV_X1 NOT_1442( .ZN(II4055), .A(n1748gat) );
  INV_X1 NOT_1443( .ZN(n1747gat), .A(II4055) );
  INV_X1 NOT_1444( .ZN(II4067), .A(n1675gat) );
  INV_X1 NOT_1445( .ZN(n1674gat), .A(II4067) );
  INV_X1 NOT_1446( .ZN(n1403gat), .A(n1402gat) );
  INV_X8 NOT_1447( .ZN(II4081), .A(n1807gat) );
  INV_X8 NOT_1448( .ZN(n1806gat), .A(II4081) );
  INV_X8 NOT_1449( .ZN(n1634gat), .A(n1712gat) );
  INV_X1 NOT_1450( .ZN(n1338gat), .A(n1340gat) );
  INV_X1 NOT_1451( .ZN(II4105), .A(n1456gat) );
  INV_X1 NOT_1452( .ZN(n1455gat), .A(II4105) );
  INV_X1 NOT_1453( .ZN(II4108), .A(n1340gat) );
  INV_X1 NOT_1454( .ZN(n1339gat), .A(II4108) );
  INV_X1 NOT_1455( .ZN(n1505gat), .A(n2980gat) );
  INV_X1 NOT_1456( .ZN(II4117), .A(n1505gat) );
  INV_X1 NOT_1457( .ZN(n2758gat), .A(II4117) );
  INV_X1 NOT_1458( .ZN(n2755gat), .A(n2758gat) );
  INV_X1 NOT_1459( .ZN(n1546gat), .A(n2980gat) );
  INV_X1 NOT_1460( .ZN(II4122), .A(n1546gat) );
  INV_X1 NOT_1461( .ZN(n2752gat), .A(II4122) );
  INV_X1 NOT_1462( .ZN(n2748gat), .A(n2752gat) );
  INV_X1 NOT_1463( .ZN(n2012gat), .A(n2016gat) );
  INV_X1 NOT_1464( .ZN(n2002gat), .A(n2008gat) );
  INV_X1 NOT_1465( .ZN(II4129), .A(n3097gat) );
  INV_X1 NOT_1466( .ZN(n2858gat), .A(II4129) );
  INV_X1 NOT_1467( .ZN(n2857gat), .A(n2858gat) );
  INV_X1 NOT_1468( .ZN(II4135), .A(n3098gat) );
  INV_X1 NOT_1469( .ZN(n2766gat), .A(II4135) );
  INV_X1 NOT_1470( .ZN(II4138), .A(n2766gat) );
  INV_X1 NOT_1471( .ZN(n2765gat), .A(II4138) );
  INV_X1 NOT_1472( .ZN(n1684gat), .A(n1759gat) );
  INV_X1 NOT_1473( .ZN(n1632gat), .A(II4145) );
  INV_X1 NOT_1474( .ZN(II4157), .A(n1525gat) );
  INV_X1 NOT_1475( .ZN(n1524gat), .A(II4157) );
  INV_X1 NOT_1476( .ZN(n1862gat), .A(n1863gat) );
  INV_X1 NOT_1477( .ZN(n1919gat), .A(n1860gat) );
  INV_X1 NOT_1478( .ZN(n1460gat), .A(n1462gat) );
  INV_X1 NOT_1479( .ZN(II4185), .A(n1596gat) );
  INV_X1 NOT_1480( .ZN(n1595gat), .A(II4185) );
  INV_X1 NOT_1481( .ZN(n1454gat), .A(n1469gat) );
  INV_X1 NOT_1482( .ZN(n1468gat), .A(n1519gat) );
  INV_X1 NOT_1483( .ZN(II4194), .A(n1462gat) );
  INV_X1 NOT_1484( .ZN(n1461gat), .A(II4194) );
  INV_X1 NOT_1485( .ZN(n1477gat), .A(n2984gat) );
  INV_X1 NOT_1486( .ZN(n1594gat), .A(n1596gat) );
  INV_X1 NOT_1487( .ZN(II4212), .A(n1588gat) );
  INV_X1 NOT_1488( .ZN(n1587gat), .A(II4212) );
  INV_X1 NOT_1489( .ZN(n1681gat), .A(II4217) );
  INV_X1 NOT_1490( .ZN(II4222), .A(n1761gat) );
  INV_X1 NOT_1491( .ZN(n2751gat), .A(II4222) );
  INV_X1 NOT_1492( .ZN(n2747gat), .A(n2751gat) );
  INV_X1 NOT_1493( .ZN(II4227), .A(n1760gat) );
  INV_X1 NOT_1494( .ZN(n2743gat), .A(II4227) );
  INV_X1 NOT_1495( .ZN(n2739gat), .A(n2743gat) );
  INV_X1 NOT_1496( .ZN(n1978gat), .A(n2286gat) );
  INV_X1 NOT_1497( .ZN(II4233), .A(n1721gat) );
  INV_X1 NOT_1498( .ZN(n2808gat), .A(II4233) );
  INV_X1 NOT_1499( .ZN(II4236), .A(n2808gat) );
  INV_X8 NOT_1500( .ZN(n2804gat), .A(II4236) );
  INV_X8 NOT_1501( .ZN(n517gat), .A(n518gat) );
  INV_X1 NOT_1502( .ZN(n417gat), .A(n418gat) );
  INV_X1 NOT_1503( .ZN(n413gat), .A(n411gat) );
  INV_X1 NOT_1504( .ZN(n412gat), .A(n522gat) );
  INV_X1 NOT_1505( .ZN(n406gat), .A(n516gat) );
  INV_X1 NOT_1506( .ZN(n407gat), .A(n355gat) );
  INV_X1 NOT_1507( .ZN(n290gat), .A(n525gat) );
  INV_X1 NOT_1508( .ZN(n527gat), .A(n356gat) );
  INV_X1 NOT_1509( .ZN(n416gat), .A(n415gat) );
  INV_X1 NOT_1510( .ZN(n528gat), .A(n521gat) );
  INV_X1 NOT_1511( .ZN(n358gat), .A(n532gat) );
  INV_X1 NOT_1512( .ZN(n639gat), .A(n523gat) );
  INV_X1 NOT_1513( .ZN(n1111gat), .A(n635gat) );
  INV_X1 NOT_1514( .ZN(n524gat), .A(n414gat) );
  INV_X1 NOT_1515( .ZN(n1112gat), .A(n630gat) );
  INV_X1 NOT_1516( .ZN(n741gat), .A(n629gat) );
  INV_X1 NOT_1517( .ZN(n633gat), .A(n634gat) );
  INV_X1 NOT_1518( .ZN(n926gat), .A(n632gat) );
  INV_X1 NOT_1519( .ZN(n670gat), .A(n636gat) );
  INV_X1 NOT_1520( .ZN(n1123gat), .A(n632gat) );
  INV_X1 NOT_1521( .ZN(n1007gat), .A(n635gat) );
  INV_X1 NOT_1522( .ZN(n1006gat), .A(n630gat) );
  INV_X1 NOT_1523( .ZN(II4309), .A(n2941gat) );
  INV_X1 NOT_1524( .ZN(n2814gat), .A(II4309) );
  INV_X1 NOT_1525( .ZN(II4312), .A(n2814gat) );
  INV_X1 NOT_1526( .ZN(n2811gat), .A(II4312) );
  INV_X1 NOT_1527( .ZN(n1002gat), .A(n2946gat) );
  INV_X1 NOT_1528( .ZN(II4329), .A(n2950gat) );
  INV_X1 NOT_1529( .ZN(n2813gat), .A(II4329) );
  INV_X1 NOT_1530( .ZN(II4332), .A(n2813gat) );
  INV_X1 NOT_1531( .ZN(n2810gat), .A(II4332) );
  INV_X1 NOT_1532( .ZN(n888gat), .A(n2933gat) );
  INV_X1 NOT_1533( .ZN(II4349), .A(n2935gat) );
  INV_X1 NOT_1534( .ZN(n2818gat), .A(II4349) );
  INV_X1 NOT_1535( .ZN(II4352), .A(n2818gat) );
  INV_X1 NOT_1536( .ZN(n2816gat), .A(II4352) );
  INV_X1 NOT_1537( .ZN(n898gat), .A(n2940gat) );
  INV_X1 NOT_1538( .ZN(II4369), .A(n2937gat) );
  INV_X1 NOT_1539( .ZN(n2817gat), .A(II4369) );
  INV_X1 NOT_1540( .ZN(II4372), .A(n2817gat) );
  INV_X1 NOT_1541( .ZN(n2815gat), .A(II4372) );
  INV_X1 NOT_1542( .ZN(n1179gat), .A(n2947gat) );
  INV_X1 NOT_1543( .ZN(II4389), .A(n2956gat) );
  INV_X1 NOT_1544( .ZN(n2824gat), .A(II4389) );
  INV_X1 NOT_1545( .ZN(II4392), .A(n2824gat) );
  INV_X1 NOT_1546( .ZN(n2821gat), .A(II4392) );
  INV_X1 NOT_1547( .ZN(n897gat), .A(n2939gat) );
  INV_X1 NOT_1548( .ZN(II4409), .A(n2938gat) );
  INV_X1 NOT_1549( .ZN(n2823gat), .A(II4409) );
  INV_X1 NOT_1550( .ZN(II4412), .A(n2823gat) );
  INV_X1 NOT_1551( .ZN(n2820gat), .A(II4412) );
  INV_X1 NOT_1552( .ZN(n894gat), .A(n2932gat) );
  INV_X1 NOT_1553( .ZN(II4429), .A(n2936gat) );
  INV_X1 NOT_1554( .ZN(n2829gat), .A(II4429) );
  INV_X1 NOT_1555( .ZN(II4432), .A(n2829gat) );
  INV_X1 NOT_1556( .ZN(n2826gat), .A(II4432) );
  INV_X8 NOT_1557( .ZN(n1180gat), .A(n2948gat) );
  INV_X8 NOT_1558( .ZN(II4449), .A(n2955gat) );
  INV_X1 NOT_1559( .ZN(n2828gat), .A(II4449) );
  INV_X1 NOT_1560( .ZN(II4452), .A(n2828gat) );
  INV_X1 NOT_1561( .ZN(n2825gat), .A(II4452) );
  INV_X1 NOT_1562( .ZN(n671gat), .A(n673gat) );
  INV_X1 NOT_1563( .ZN(n628gat), .A(n631gat) );
  INV_X1 NOT_1564( .ZN(n976gat), .A(n628gat) );
  INV_X1 NOT_1565( .ZN(II4475), .A(n2951gat) );
  INV_X1 NOT_1566( .ZN(n2807gat), .A(II4475) );
  INV_X1 NOT_1567( .ZN(II4478), .A(n2807gat) );
  INV_X1 NOT_1568( .ZN(n2803gat), .A(II4478) );
  INV_X1 NOT_1569( .ZN(n2127gat), .A(n2389gat) );
  INV_X1 NOT_1570( .ZN(II4482), .A(n2127gat) );
  INV_X1 NOT_1571( .ZN(n2682gat), .A(II4482) );
  INV_X1 NOT_1572( .ZN(II4485), .A(n2682gat) );
  INV_X1 NOT_1573( .ZN(n2678gat), .A(II4485) );
  INV_X1 NOT_1574( .ZN(n2046gat), .A(n2269gat) );
  INV_X1 NOT_1575( .ZN(II4489), .A(n2046gat) );
  INV_X1 NOT_1576( .ZN(n2681gat), .A(II4489) );
  INV_X1 NOT_1577( .ZN(II4492), .A(n2681gat) );
  INV_X1 NOT_1578( .ZN(n2677gat), .A(II4492) );
  INV_X1 NOT_1579( .ZN(n1708gat), .A(n2338gat) );
  INV_X1 NOT_1580( .ZN(II4496), .A(n1708gat) );
  INV_X1 NOT_1581( .ZN(n2688gat), .A(II4496) );
  INV_X1 NOT_1582( .ZN(II4499), .A(n2688gat) );
  INV_X1 NOT_1583( .ZN(n2686gat), .A(II4499) );
  INV_X1 NOT_1584( .ZN(n455gat), .A(n291gat) );
  INV_X1 NOT_1585( .ZN(n2237gat), .A(n2646gat) );
  INV_X1 NOT_1586( .ZN(II4506), .A(n2764gat) );
  INV_X1 NOT_1587( .ZN(n2763gat), .A(II4506) );
  INV_X1 NOT_1588( .ZN(n1782gat), .A(n2971gat) );
  INV_X1 NOT_1589( .ZN(II4512), .A(n2762gat) );
  INV_X1 NOT_1590( .ZN(n2760gat), .A(II4512) );
  INV_X1 NOT_1591( .ZN(n2325gat), .A(n3010gat) );
  INV_X1 NOT_1592( .ZN(II4518), .A(n2761gat) );
  INV_X1 NOT_1593( .ZN(n2759gat), .A(II4518) );
  INV_X1 NOT_1594( .ZN(n2245gat), .A(n504gat) );
  INV_X1 NOT_1595( .ZN(II4524), .A(n2757gat) );
  INV_X1 NOT_1596( .ZN(n2754gat), .A(II4524) );
  INV_X1 NOT_1597( .ZN(n2244gat), .A(n567gat) );
  INV_X1 NOT_1598( .ZN(II4530), .A(n2756gat) );
  INV_X1 NOT_1599( .ZN(n2753gat), .A(II4530) );
  INV_X1 NOT_1600( .ZN(n2243gat), .A(n55gat) );
  INV_X1 NOT_1601( .ZN(II4536), .A(n2750gat) );
  INV_X1 NOT_1602( .ZN(n2746gat), .A(II4536) );
  INV_X1 NOT_1603( .ZN(n2246gat), .A(n933gat) );
  INV_X1 NOT_1604( .ZN(II4542), .A(n2749gat) );
  INV_X1 NOT_1605( .ZN(n2745gat), .A(II4542) );
  INV_X1 NOT_1606( .ZN(n2384gat), .A(n43gat) );
  INV_X1 NOT_1607( .ZN(II4548), .A(n2742gat) );
  INV_X1 NOT_1608( .ZN(n2738gat), .A(II4548) );
  INV_X1 NOT_1609( .ZN(n2385gat), .A(n748gat) );
  INV_X16 NOT_1610( .ZN(II4554), .A(n2741gat) );
  INV_X16 NOT_1611( .ZN(n2737gat), .A(II4554) );
  INV_X16 NOT_1612( .ZN(n1286gat), .A(n1269gat) );
  INV_X1 NOT_1613( .ZN(II4558), .A(n1286gat) );
  INV_X1 NOT_1614( .ZN(n2687gat), .A(II4558) );
  INV_X1 NOT_1615( .ZN(n2685gat), .A(n2687gat) );
  INV_X1 NOT_1616( .ZN(n1328gat), .A(n1224gat) );
  INV_X1 NOT_1617( .ZN(n1381gat), .A(n1328gat) );
  INV_X1 NOT_1618( .ZN(n1384gat), .A(n2184gat) );
  INV_X1 NOT_1619( .ZN(II4566), .A(n2694gat) );
  INV_X1 NOT_1620( .ZN(n2690gat), .A(II4566) );
  INV_X1 NOT_1621( .ZN(n1382gat), .A(n1280gat) );
  INV_X1 NOT_1622( .ZN(n1451gat), .A(n1382gat) );
  INV_X1 NOT_1623( .ZN(n1453gat), .A(n2187gat) );
  INV_X1 NOT_1624( .ZN(II4573), .A(n2693gat) );
  INV_X1 NOT_1625( .ZN(n2689gat), .A(II4573) );
  INV_X1 NOT_1626( .ZN(n927gat), .A(n1133gat) );
  INV_X1 NOT_1627( .ZN(n925gat), .A(n927gat) );
  INV_X1 NOT_1628( .ZN(n1452gat), .A(n2049gat) );
  INV_X1 NOT_1629( .ZN(II4580), .A(n2702gat) );
  INV_X1 NOT_1630( .ZN(n2698gat), .A(II4580) );
  INV_X1 NOT_1631( .ZN(n923gat), .A(n1043gat) );
  INV_X1 NOT_1632( .ZN(n921gat), .A(n923gat) );
  INV_X1 NOT_1633( .ZN(n1890gat), .A(n2328gat) );
  INV_X1 NOT_1634( .ZN(II4587), .A(n2701gat) );
  INV_X1 NOT_1635( .ZN(n2697gat), .A(II4587) );
  INV_X1 NOT_1636( .ZN(n850gat), .A(n929gat) );
  INV_X1 NOT_1637( .ZN(n739gat), .A(n850gat) );
  INV_X1 NOT_1638( .ZN(n1841gat), .A(n2058gat) );
  INV_X1 NOT_1639( .ZN(II4594), .A(n2709gat) );
  INV_X1 NOT_1640( .ZN(n2706gat), .A(II4594) );
  INV_X1 NOT_1641( .ZN(n922gat), .A(n1119gat) );
  INV_X1 NOT_1642( .ZN(n848gat), .A(n922gat) );
  INV_X1 NOT_1643( .ZN(n2047gat), .A(n2209gat) );
  INV_X1 NOT_1644( .ZN(II4601), .A(n2708gat) );
  INV_X1 NOT_1645( .ZN(n2705gat), .A(II4601) );
  INV_X1 NOT_1646( .ZN(n924gat), .A(n1070gat) );
  INV_X1 NOT_1647( .ZN(n849gat), .A(n924gat) );
  INV_X1 NOT_1648( .ZN(n2050gat), .A(n2146gat) );
  INV_X1 NOT_1649( .ZN(II4608), .A(n2799gat) );
  INV_X1 NOT_1650( .ZN(n2796gat), .A(II4608) );
  INV_X1 NOT_1651( .ZN(n1118gat), .A(n1033gat) );
  INV_X1 NOT_1652( .ZN(n1032gat), .A(n1118gat) );
  INV_X1 NOT_1653( .ZN(n2054gat), .A(n2281gat) );
  INV_X1 NOT_1654( .ZN(II4615), .A(n2798gat) );
  INV_X1 NOT_1655( .ZN(n2795gat), .A(II4615) );
  INV_X1 NOT_1656( .ZN(II4620), .A(n1745gat) );
  INV_X1 NOT_1657( .ZN(n2806gat), .A(II4620) );
  INV_X1 NOT_1658( .ZN(II4623), .A(n2806gat) );
  INV_X1 NOT_1659( .ZN(n2802gat), .A(II4623) );
  INV_X1 NOT_1660( .ZN(II4626), .A(n1871gat) );
  INV_X1 NOT_1661( .ZN(n1870gat), .A(II4626) );
  INV_X1 NOT_1662( .ZN(n1086gat), .A(n1870gat) );
  INV_X1 NOT_1663( .ZN(II4630), .A(n1086gat) );
  INV_X1 NOT_1664( .ZN(n2805gat), .A(II4630) );
  INV_X1 NOT_1665( .ZN(II4633), .A(n2805gat) );
  INV_X1 NOT_1666( .ZN(n2801gat), .A(II4633) );
  INV_X1 NOT_1667( .ZN(n67gat), .A(n85gat) );
  INV_X1 NOT_1668( .ZN(n71gat), .A(n180gat) );
  INV_X1 NOT_1669( .ZN(n1840gat), .A(n1892gat) );
  INV_X16 NOT_1670( .ZN(II4642), .A(n2812gat) );
  INV_X32 NOT_1671( .ZN(n2809gat), .A(II4642) );
  INV_X1 NOT_1672( .ZN(n76gat), .A(n82gat) );
  INV_X1 NOT_1673( .ZN(n14gat), .A(n186gat) );
  INV_X1 NOT_1674( .ZN(n1842gat), .A(n1711gat) );
  INV_X1 NOT_1675( .ZN(II4651), .A(n2822gat) );
  INV_X1 NOT_1676( .ZN(n2819gat), .A(II4651) );
  INV_X1 NOT_1677( .ZN(II4654), .A(n2819gat) );
  INV_X1 NOT_1678( .ZN(n3104gat), .A(II4654) );
  INV_X1 NOT_1679( .ZN(II4657), .A(n2809gat) );
  INV_X1 NOT_1680( .ZN(n3105gat), .A(II4657) );
  INV_X1 NOT_1681( .ZN(II4660), .A(n2801gat) );
  INV_X1 NOT_1682( .ZN(n3106gat), .A(II4660) );
  INV_X1 NOT_1683( .ZN(II4663), .A(n2802gat) );
  INV_X1 NOT_1684( .ZN(n3107gat), .A(II4663) );
  INV_X1 NOT_1685( .ZN(II4666), .A(n2795gat) );
  INV_X1 NOT_1686( .ZN(n3108gat), .A(II4666) );
  INV_X1 NOT_1687( .ZN(II4669), .A(n2796gat) );
  INV_X1 NOT_1688( .ZN(n3109gat), .A(II4669) );
  INV_X1 NOT_1689( .ZN(II4672), .A(n2705gat) );
  INV_X1 NOT_1690( .ZN(n3110gat), .A(II4672) );
  INV_X1 NOT_1691( .ZN(II4675), .A(n2706gat) );
  INV_X1 NOT_1692( .ZN(n3111gat), .A(II4675) );
  INV_X1 NOT_1693( .ZN(II4678), .A(n2697gat) );
  INV_X1 NOT_1694( .ZN(n3112gat), .A(II4678) );
  INV_X1 NOT_1695( .ZN(II4681), .A(n2698gat) );
  INV_X1 NOT_1696( .ZN(n3113gat), .A(II4681) );
  INV_X1 NOT_1697( .ZN(II4684), .A(n2689gat) );
  INV_X1 NOT_1698( .ZN(n3114gat), .A(II4684) );
  INV_X1 NOT_1699( .ZN(II4687), .A(n2690gat) );
  INV_X1 NOT_1700( .ZN(n3115gat), .A(II4687) );
  INV_X1 NOT_1701( .ZN(II4690), .A(n2685gat) );
  INV_X1 NOT_1702( .ZN(n3116gat), .A(II4690) );
  INV_X1 NOT_1703( .ZN(II4693), .A(n2737gat) );
  INV_X1 NOT_1704( .ZN(n3117gat), .A(II4693) );
  INV_X1 NOT_1705( .ZN(II4696), .A(n2738gat) );
  INV_X1 NOT_1706( .ZN(n3118gat), .A(II4696) );
  INV_X1 NOT_1707( .ZN(II4699), .A(n2745gat) );
  INV_X1 NOT_1708( .ZN(n3119gat), .A(II4699) );
  INV_X1 NOT_1709( .ZN(II4702), .A(n2746gat) );
  INV_X1 NOT_1710( .ZN(n3120gat), .A(II4702) );
  INV_X1 NOT_1711( .ZN(II4705), .A(n2753gat) );
  INV_X1 NOT_1712( .ZN(n3121gat), .A(II4705) );
  INV_X1 NOT_1713( .ZN(II4708), .A(n2754gat) );
  INV_X1 NOT_1714( .ZN(n3122gat), .A(II4708) );
  INV_X1 NOT_1715( .ZN(II4711), .A(n2759gat) );
  INV_X1 NOT_1716( .ZN(n3123gat), .A(II4711) );
  INV_X1 NOT_1717( .ZN(II4714), .A(n2760gat) );
  INV_X1 NOT_1718( .ZN(n3124gat), .A(II4714) );
  INV_X1 NOT_1719( .ZN(II4717), .A(n2763gat) );
  INV_X1 NOT_1720( .ZN(n3125gat), .A(II4717) );
  INV_X1 NOT_1721( .ZN(II4720), .A(n2686gat) );
  INV_X1 NOT_1722( .ZN(n3126gat), .A(II4720) );
  INV_X1 NOT_1723( .ZN(II4723), .A(n2677gat) );
  INV_X1 NOT_1724( .ZN(n3127gat), .A(II4723) );
  INV_X32 NOT_1725( .ZN(II4726), .A(n2678gat) );
  INV_X32 NOT_1726( .ZN(n3128gat), .A(II4726) );
  INV_X32 NOT_1727( .ZN(II4729), .A(n2803gat) );
  INV_X1 NOT_1728( .ZN(n3129gat), .A(II4729) );
  INV_X1 NOT_1729( .ZN(II4732), .A(n2825gat) );
  INV_X1 NOT_1730( .ZN(n3130gat), .A(II4732) );
  INV_X1 NOT_1731( .ZN(II4735), .A(n2826gat) );
  INV_X1 NOT_1732( .ZN(n3131gat), .A(II4735) );
  INV_X1 NOT_1733( .ZN(II4738), .A(n2820gat) );
  INV_X1 NOT_1734( .ZN(n3132gat), .A(II4738) );
  INV_X1 NOT_1735( .ZN(II4741), .A(n2821gat) );
  INV_X1 NOT_1736( .ZN(n3133gat), .A(II4741) );
  INV_X1 NOT_1737( .ZN(II4744), .A(n2815gat) );
  INV_X1 NOT_1738( .ZN(n3134gat), .A(II4744) );
  INV_X1 NOT_1739( .ZN(II4747), .A(n2816gat) );
  INV_X1 NOT_1740( .ZN(n3135gat), .A(II4747) );
  INV_X1 NOT_1741( .ZN(II4750), .A(n2810gat) );
  INV_X1 NOT_1742( .ZN(n3136gat), .A(II4750) );
  INV_X1 NOT_1743( .ZN(II4753), .A(n2811gat) );
  INV_X1 NOT_1744( .ZN(n3137gat), .A(II4753) );
  INV_X1 NOT_1745( .ZN(II4756), .A(n2804gat) );
  INV_X1 NOT_1746( .ZN(n3138gat), .A(II4756) );
  INV_X1 NOT_1747( .ZN(II4759), .A(n2739gat) );
  INV_X1 NOT_1748( .ZN(n3139gat), .A(II4759) );
  INV_X1 NOT_1749( .ZN(II4762), .A(n2747gat) );
  INV_X1 NOT_1750( .ZN(n3140gat), .A(II4762) );
  INV_X1 NOT_1751( .ZN(II4765), .A(n2748gat) );
  INV_X1 NOT_1752( .ZN(n3141gat), .A(II4765) );
  INV_X1 NOT_1753( .ZN(II4768), .A(n2755gat) );
  INV_X1 NOT_1754( .ZN(n3142gat), .A(II4768) );
  INV_X1 NOT_1755( .ZN(II4771), .A(n2797gat) );
  INV_X1 NOT_1756( .ZN(n3143gat), .A(II4771) );
  INV_X1 NOT_1757( .ZN(II4774), .A(n2740gat) );
  INV_X1 NOT_1758( .ZN(n3144gat), .A(II4774) );
  INV_X1 NOT_1759( .ZN(II4777), .A(n2699gat) );
  INV_X1 NOT_1760( .ZN(n3145gat), .A(II4777) );
  INV_X1 NOT_1761( .ZN(II4780), .A(n2691gat) );
  INV_X1 NOT_1762( .ZN(n3146gat), .A(II4780) );
  INV_X1 NOT_1763( .ZN(II4783), .A(n2827gat) );
  INV_X1 NOT_1764( .ZN(n3147gat), .A(II4783) );
  INV_X1 NOT_1765( .ZN(II4786), .A(n2679gat) );
  INV_X1 NOT_1766( .ZN(n3148gat), .A(II4786) );
  INV_X1 NOT_1767( .ZN(II4789), .A(n2692gat) );
  INV_X1 NOT_1768( .ZN(n3149gat), .A(II4789) );
  INV_X1 NOT_1769( .ZN(II4792), .A(n2680gat) );
  INV_X1 NOT_1770( .ZN(n3150gat), .A(II4792) );
  INV_X1 NOT_1771( .ZN(II4795), .A(n2700gat) );
  INV_X1 NOT_1772( .ZN(n3151gat), .A(II4795) );
  INV_X1 NOT_1773( .ZN(II4798), .A(n2707gat) );
  INV_X1 NOT_1774( .ZN(n3152gat), .A(II4798) );
  OR2_X1 OR2_0( .ZN(n2897gat), .A1(n648gat), .A2(n442gat) );
  OR4_X2 OR4_0( .ZN(n1213gat), .A1(n1214gat), .A2(n1215gat), .A3(n1216gat), .A4(n1217gat) );
  OR2_X2 OR2_1( .ZN(n2906gat), .A1(n745gat), .A2(n638gat) );
  OR2_X2 OR2_2( .ZN(n2889gat), .A1(n423gat), .A2(n362gat) );
  OR4_X2 OR4_1( .ZN(n748gat), .A1(n749gat), .A2(n750gat), .A3(n751gat), .A4(n752gat) );
  OR4_X1 OR4_2( .ZN(n258gat), .A1(n259gat), .A2(n260gat), .A3(n261gat), .A4(n262gat) );
  OR4_X1 OR4_3( .ZN(n1013gat), .A1(n1014gat), .A2(n1015gat), .A3(n1016gat), .A4(n1017gat) );
  OR4_X1 OR4_4( .ZN(n475gat), .A1(n476gat), .A2(n477gat), .A3(n478gat), .A4(n479gat) );
  OR4_X1 OR4_5( .ZN(n43gat), .A1(n44gat), .A2(n45gat), .A3(n46gat), .A4(n47gat) );
  OR2_X1 OR2_3( .ZN(n2786gat), .A1(n3091gat), .A2(n3092gat) );
  OR4_X1 OR4_6( .ZN(n167gat), .A1(n168gat), .A2(n169gat), .A3(n170gat), .A4(n171gat) );
  OR4_X1 OR4_7( .ZN(n906gat), .A1(n907gat), .A2(n908gat), .A3(n909gat), .A4(n910gat) );
  OR4_X1 OR4_8( .ZN(n343gat), .A1(n344gat), .A2(n345gat), .A3(n346gat), .A4(n347gat) );
  OR4_X1 OR4_9( .ZN(n55gat), .A1(n56gat), .A2(n57gat), .A3(n58gat), .A4(n59gat) );
  OR2_X1 OR2_4( .ZN(n2914gat), .A1(n768gat), .A2(n655gat) );
  OR2_X1 OR2_5( .ZN(n2928gat), .A1(n963gat), .A2(n868gat) );
  OR2_X1 OR2_6( .ZN(n2927gat), .A1(n962gat), .A2(n959gat) );
  OR4_X1 OR4_10( .ZN(n944gat), .A1(n945gat), .A2(n946gat), .A3(n947gat), .A4(n948gat) );
  OR2_X1 OR2_7( .ZN(n2896gat), .A1(n647gat), .A2(n441gat) );
  OR2_X1 OR2_8( .ZN(n2922gat), .A1(n967gat), .A2(n792gat) );
  OR4_X1 OR4_11( .ZN(n1228gat), .A1(n1229gat), .A2(n1230gat), .A3(n1231gat), .A4(n1232gat) );
  OR2_X1 OR2_9( .ZN(n2894gat), .A1(n443gat), .A2(n439gat) );
  OR2_X1 OR2_10( .ZN(n2921gat), .A1(n966gat), .A2(n790gat) );
  OR2_X1 OR2_11( .ZN(n2895gat), .A1(n444gat), .A2(n440gat) );
  OR4_X1 OR4_12( .ZN(n1050gat), .A1(n1051gat), .A2(n1052gat), .A3(n1053gat), .A4(n1054gat) );
  OR4_X1 OR4_13( .ZN(n933gat), .A1(n934gat), .A2(n935gat), .A3(n936gat), .A4(n937gat) );
  OR4_X1 OR4_14( .ZN(n709gat), .A1(n710gat), .A2(n711gat), .A3(n712gat), .A4(n713gat) );
  OR4_X1 OR4_15( .ZN(n728gat), .A1(n729gat), .A2(n730gat), .A3(n731gat), .A4(n732gat) );
  OR4_X1 OR4_16( .ZN(n493gat), .A1(n494gat), .A2(n495gat), .A3(n496gat), .A4(n497gat) );
  OR4_X1 OR4_17( .ZN(n504gat), .A1(n505gat), .A2(n506gat), .A3(n507gat), .A4(n508gat) );
  OR3_X1 OR3_0( .ZN(II1277), .A1(n2860gat), .A2(n2855gat), .A3(n2863gat) );
  OR3_X1 OR3_1( .ZN(II1278), .A1(n740gat), .A2(n3030gat), .A3(II1277) );
  OR2_X1 OR2_12( .ZN(n2913gat), .A1(n767gat), .A2(n653gat) );
  OR2_X1 OR2_13( .ZN(n2920gat), .A1(n867gat), .A2(n771gat) );
  OR2_X1 OR2_14( .ZN(n2905gat), .A1(n964gat), .A2(n961gat) );
  OR4_X1 OR4_18( .ZN(n803gat), .A1(n804gat), .A2(n805gat), .A3(n806gat), .A4(n807gat) );
  OR4_X1 OR4_19( .ZN(n586gat), .A1(n587gat), .A2(n588gat), .A3(n589gat), .A4(n590gat) );
  OR2_X1 OR2_15( .ZN(n2898gat), .A1(n447gat), .A2(n445gat) );
  OR4_X1 OR4_20( .ZN(n686gat), .A1(n687gat), .A2(n688gat), .A3(n689gat), .A4(n690gat) );
  OR4_X1 OR4_21( .ZN(n567gat), .A1(n568gat), .A2(n569gat), .A3(n570gat), .A4(n571gat) );
  OR3_X1 OR3_2( .ZN(II1515), .A1(n2474gat), .A2(n2524gat), .A3(n2831gat) );
  OR3_X1 OR3_3( .ZN(II1516), .A1(n2466gat), .A2(n2462gat), .A3(II1515) );
  OR3_X1 OR3_4( .ZN(II1584), .A1(n2353gat), .A2(n2284gat), .A3(n2354gat) );
  OR3_X1 OR3_5( .ZN(II1585), .A1(n2356gat), .A2(n2214gat), .A3(II1584) );
  OR2_X1 OR2_16( .ZN(n2989gat), .A1(n1693gat), .A2(n1692gat) );
  OR3_X1 OR3_6( .ZN(II1723), .A1(n2354gat), .A2(n2353gat), .A3(n2214gat) );
  OR3_X1 OR3_7( .ZN(II1724), .A1(n2355gat), .A2(n2443gat), .A3(II1723) );
  OR3_X1 OR3_8( .ZN(II1733), .A1(n2286gat), .A2(n2428gat), .A3(n2289gat) );
  OR3_X1 OR3_9( .ZN(II1734), .A1(n1604gat), .A2(n2214gat), .A3(II1733) );
  OR2_X1 OR2_17( .ZN(n2918gat), .A1(n769gat), .A2(n759gat) );
  OR2_X1 OR2_18( .ZN(n2952gat), .A1(n1076gat), .A2(n1075gat) );
  OR2_X1 OR2_19( .ZN(n2919gat), .A1(n766gat), .A2(n760gat) );
  OR4_X1 OR4_22( .ZN(n1184gat), .A1(n1185gat), .A2(n1186gat), .A3(n1187gat), .A4(n1188gat) );
  OR2_X1 OR2_20( .ZN(n2910gat), .A1(n645gat), .A2(n644gat) );
  OR2_X1 OR2_21( .ZN(n2907gat), .A1(n646gat), .A2(n641gat) );
  OR2_X1 OR2_22( .ZN(n2970gat), .A1(n1383gat), .A2(n1327gat) );
  OR2_X1 OR2_23( .ZN(n2911gat), .A1(n761gat), .A2(n651gat) );
  OR2_X1 OR2_24( .ZN(n2912gat), .A1(n762gat), .A2(n652gat) );
  OR2_X1 OR2_25( .ZN(n2909gat), .A1(n765gat), .A2(n643gat) );
  OR4_X1 OR4_23( .ZN(n1201gat), .A1(n1202gat), .A2(n1203gat), .A3(n1204gat), .A4(n1205gat) );
  OR4_X1 OR4_24( .ZN(n1269gat), .A1(n1270gat), .A2(n1271gat), .A3(n1272gat), .A4(n1273gat) );
  OR2_X1 OR2_26( .ZN(n2908gat), .A1(n763gat), .A2(n642gat) );
  OR2_X1 OR2_27( .ZN(n2971gat), .A1(n1287gat), .A2(n1285gat) );
  OR3_X1 OR3_10( .ZN(n2904gat), .A1(n793gat), .A2(n664gat), .A3(n556gat) );
  OR3_X1 OR3_11( .ZN(n2891gat), .A1(n795gat), .A2(n656gat), .A3(n368gat) );
  OR3_X1 OR3_12( .ZN(n2903gat), .A1(n794gat), .A2(n773gat), .A3(n662gat) );
  OR3_X1 OR3_13( .ZN(n2915gat), .A1(n965gat), .A2(n960gat), .A3(n661gat) );
  OR4_X1 OR4_25( .ZN(n779gat), .A1(n780gat), .A2(n781gat), .A3(n782gat), .A4(n783gat) );
  OR3_X1 OR3_14( .ZN(n2901gat), .A1(n558gat), .A2(n555gat), .A3(n450gat) );
  OR3_X1 OR3_15( .ZN(n2890gat), .A1(n654gat), .A2(n557gat), .A3(n371gat) );
  OR2_X1 OR2_28( .ZN(n2876gat), .A1(n874gat), .A2(n132gat) );
  OR3_X1 OR3_16( .ZN(n2888gat), .A1(n663gat), .A2(n649gat), .A3(n449gat) );
  OR3_X1 OR3_17( .ZN(n2887gat), .A1(n791gat), .A2(n650gat), .A3(n370gat) );
  OR3_X2 OR3_18( .ZN(n2886gat), .A1(n774gat), .A2(n764gat), .A3(n369gat) );
  OR4_X2 OR4_26( .ZN(n221gat), .A1(n222gat), .A2(n223gat), .A3(n224gat), .A4(n225gat) );
  OR4_X2 OR4_27( .ZN(n120gat), .A1(n121gat), .A2(n122gat), .A3(n123gat), .A4(n124gat) );
  OR2_X1 OR2_29( .ZN(n3010gat), .A1(n2460gat), .A2(n2423gat) );
  OR2_X1 OR2_30( .ZN(n3016gat), .A1(n2596gat), .A2(n2595gat) );
  OR4_X1 OR4_28( .ZN(n2568gat), .A1(n2569gat), .A2(n2570gat), .A3(n2571gat), .A4(n2572gat) );
  OR4_X1 OR4_29( .ZN(n2409gat), .A1(n2410gat), .A2(n2411gat), .A3(n2412gat), .A4(n2413gat) );
  OR2_X1 OR2_31( .ZN(n2579gat), .A1(n2580gat), .A2(n2581gat) );
  OR2_X1 OR2_32( .ZN(n3014gat), .A1(n2567gat), .A2(n2499gat) );
  OR2_X1 OR2_33( .ZN(n2880gat), .A1(n299gat), .A2(n207gat) );
  OR2_X1 OR2_34( .ZN(n2646gat), .A1(n2647gat), .A2(n2648gat) );
  OR4_X1 OR4_30( .ZN(n2601gat), .A1(n2602gat), .A2(n2603gat), .A3(n2604gat), .A4(n2605gat) );
  OR4_X1 OR4_31( .ZN(n2545gat), .A1(n2546gat), .A2(n2547gat), .A3(n2548gat), .A4(n2549gat) );
  OR2_X1 OR2_35( .ZN(n2613gat), .A1(n2614gat), .A2(n2615gat) );
  OR2_X1 OR2_36( .ZN(n3013gat), .A1(n2461gat), .A2(n2421gat) );
  OR4_X1 OR4_32( .ZN(n2930gat), .A1(n1153gat), .A2(n1151gat), .A3(n982gat), .A4(n877gat) );
  OR4_X1 OR4_33( .ZN(n2957gat), .A1(n1159gat), .A2(n1158gat), .A3(n1156gat), .A4(n1155gat) );
  OR2_X1 OR2_37( .ZN(n2975gat), .A1(n1443gat), .A2(n1325gat) );
  OR2_X1 OR2_38( .ZN(n2974gat), .A1(n1321gat), .A2(n1320gat) );
  OR2_X1 OR2_39( .ZN(n2966gat), .A1(n1368gat), .A2(n1258gat) );
  OR2_X1 OR2_40( .ZN(n2979gat), .A1(n1373gat), .A2(n1372gat) );
  OR4_X1 OR4_34( .ZN(n2978gat), .A1(n1441gat), .A2(n1440gat), .A3(n1371gat), .A4(n1367gat) );
  OR2_X1 OR2_41( .ZN(n2982gat), .A1(n1504gat), .A2(n1502gat) );
  OR2_X1 OR2_42( .ZN(n2954gat), .A1(n1250gat), .A2(n1103gat) );
  OR2_X1 OR2_43( .ZN(n2964gat), .A1(n1304gat), .A2(n1249gat) );
  OR2_X1 OR2_44( .ZN(n2958gat), .A1(n1246gat), .A2(n1161gat) );
  OR2_X1 OR2_45( .ZN(n2963gat), .A1(n1291gat), .A2(n1245gat) );
  OR4_X1 OR4_35( .ZN(n2973gat), .A1(n1352gat), .A2(n1351gat), .A3(n1303gat), .A4(n1302gat) );
  OR2_X1 OR2_46( .ZN(n2953gat), .A1(n1163gat), .A2(n1102gat) );
  OR2_X1 OR2_47( .ZN(n2949gat), .A1(n1101gat), .A2(n996gat) );
  OR2_X1 OR2_48( .ZN(n2934gat), .A1(n1104gat), .A2(n887gat) );
  OR2_X1 OR2_49( .ZN(n2959gat), .A1(n1305gat), .A2(n1162gat) );
  OR4_X1 OR4_36( .ZN(n2977gat), .A1(n1360gat), .A2(n1359gat), .A3(n1358gat), .A4(n1357gat) );
  OR3_X1 OR3_19( .ZN(II2720), .A1(n1788gat), .A2(n1786gat), .A3(n1839gat) );
  OR3_X1 OR3_20( .ZN(II2721), .A1(n1884gat), .A2(n1783gat), .A3(II2720) );
  OR3_X1 OR3_21( .ZN(II2735), .A1(n1788gat), .A2(n1884gat), .A3(n1633gat) );
  OR3_X1 OR3_22( .ZN(II2736), .A1(n1785gat), .A2(n1784gat), .A3(II2735) );
  OR3_X1 OR3_23( .ZN(II2812), .A1(n1703gat), .A2(n1704gat), .A3(n1778gat) );
  OR4_X1 OR4_37( .ZN(II2813), .A1(n1609gat), .A2(n1702gat), .A3(n1700gat), .A4(II2812) );
  OR3_X1 OR3_24( .ZN(II2831), .A1(n1839gat), .A2(n1786gat), .A3(n1788gat) );
  OR3_X1 OR3_25( .ZN(II2832), .A1(n1884gat), .A2(n1784gat), .A3(II2831) );
  OR3_X1 OR3_26( .ZN(II2889), .A1(n1784gat), .A2(n1633gat), .A3(n1884gat) );
  OR3_X1 OR3_27( .ZN(II2890), .A1(n1788gat), .A2(n1786gat), .A3(II2889) );
  OR3_X1 OR3_28( .ZN(II2925), .A1(n1784gat), .A2(n1785gat), .A3(n1633gat) );
  OR3_X1 OR3_29( .ZN(II2926), .A1(n1884gat), .A2(n1787gat), .A3(II2925) );
  OR3_X1 OR3_30( .ZN(II2934), .A1(n1784gat), .A2(n1839gat), .A3(n1788gat) );
  OR3_X1 OR3_31( .ZN(II2935), .A1(n1785gat), .A2(n1884gat), .A3(II2934) );
  OR2_X1 OR2_50( .ZN(n2988gat), .A1(n1733gat), .A2(n1581gat) );
  OR2_X1 OR2_51( .ZN(n2983gat), .A1(n2079gat), .A2(n2073gat) );
  OR2_X1 OR2_52( .ZN(n2987gat), .A1(n1574gat), .A2(n1573gat) );
  OR3_X1 OR3_32( .ZN(n2992gat), .A1(n1723gat), .A2(n1647gat), .A3(n1646gat) );
  OR3_X1 OR3_33( .ZN(n2986gat), .A1(n1650gat), .A2(n1649gat), .A3(n1563gat) );
  OR3_X2 OR3_34( .ZN(n2991gat), .A1(n1654gat), .A2(n1653gat), .A3(n1644gat) );
  OR3_X2 OR3_35( .ZN(II3148), .A1(n1839gat), .A2(n1884gat), .A3(n1784gat) );
  OR3_X1 OR3_36( .ZN(II3149), .A1(n1786gat), .A2(n1787gat), .A3(II3148) );
  OR3_X1 OR3_37( .ZN(II3178), .A1(n1838gat), .A2(n1785gat), .A3(n1788gat) );
  OR3_X1 OR3_38( .ZN(II3179), .A1(n1839gat), .A2(n1784gat), .A3(II3178) );
  OR3_X1 OR3_39( .ZN(n2981gat), .A1(n1413gat), .A2(n1408gat), .A3(n1407gat) );
  OR2_X1 OR2_53( .ZN(n3000gat), .A1(n2000gat), .A2(n1999gat) );
  OR3_X1 OR3_40( .ZN(n3004gat), .A1(n2258gat), .A2(n2257gat), .A3(n2255gat) );
  OR2_X1 OR2_54( .ZN(n3003gat), .A1(n2256gat), .A2(n2251gat) );
  OR2_X1 OR2_55( .ZN(n3001gat), .A1(n2132gat), .A2(n2130gat) );
  OR2_X1 OR2_56( .ZN(n3006gat), .A1(n2253gat), .A2(n2252gat) );
  OR2_X1 OR2_57( .ZN(n3007gat), .A1(n2250gat), .A2(n2249gat) );
  OR2_X1 OR2_58( .ZN(n2990gat), .A1(n1710gat), .A2(n1630gat) );
  OR2_X1 OR2_59( .ZN(n2994gat), .A1(n1954gat), .A2(n1888gat) );
  OR3_X1 OR3_41( .ZN(n2993gat), .A1(n1894gat), .A2(n1847gat), .A3(n1846gat) );
  OR2_X1 OR2_60( .ZN(n2998gat), .A1(n2055gat), .A2(n1967gat) );
  OR3_X1 OR3_42( .ZN(n2996gat), .A1(n1960gat), .A2(n1959gat), .A3(n1957gat) );
  OR2_X1 OR2_61( .ZN(n3008gat), .A1(n2332gat), .A2(n2259gat) );
  OR2_X1 OR2_62( .ZN(n3005gat), .A1(n2211gat), .A2(n2210gat) );
  OR3_X1 OR3_43( .ZN(n2997gat), .A1(n2053gat), .A2(n2052gat), .A3(n1964gat) );
  OR2_X1 OR2_63( .ZN(n3009gat), .A1(n2350gat), .A2(n2282gat) );
  OR3_X1 OR3_44( .ZN(n3002gat), .A1(n2213gat), .A2(n2150gat), .A3(n2149gat) );
  OR2_X1 OR2_64( .ZN(n2995gat), .A1(n1962gat), .A2(n1955gat) );
  OR2_X1 OR2_65( .ZN(n2999gat), .A1(n1972gat), .A2(n1971gat) );
  OR2_X1 OR2_66( .ZN(n3011gat), .A1(n2333gat), .A2(n2331gat) );
  OR2_X1 OR2_67( .ZN(n3015gat), .A1(n2566gat), .A2(n2565gat) );
  OR3_X1 OR3_45( .ZN(n2874gat), .A1(n141gat), .A2(n38gat), .A3(n37gat) );
  OR2_X1 OR2_68( .ZN(n2917gat), .A1(n1074gat), .A2(n872gat) );
  OR2_X1 OR2_69( .ZN(n2878gat), .A1(n234gat), .A2(n137gat) );
  OR2_X1 OR2_70( .ZN(n2892gat), .A1(n378gat), .A2(n377gat) );
  OR3_X1 OR3_46( .ZN(n2885gat), .A1(n250gat), .A2(n249gat), .A3(n248gat) );
  OR3_X1 OR3_47( .ZN(n2900gat), .A1(n869gat), .A2(n453gat), .A3(n448gat) );
  OR2_X1 OR2_71( .ZN(n2883gat), .A1(n251gat), .A2(n244gat) );
  OR3_X1 OR3_48( .ZN(n2929gat), .A1(n974gat), .A2(n973gat), .A3(n870gat) );
  OR2_X1 OR2_72( .ZN(n2884gat), .A1(n246gat), .A2(n245gat) );
  OR2_X1 OR2_73( .ZN(n2902gat), .A1(n460gat), .A2(n459gat) );
  OR3_X1 OR3_49( .ZN(n2925gat), .A1(n975gat), .A2(n972gat), .A3(n969gat) );
  OR2_X1 OR2_74( .ZN(n2879gat), .A1(n145gat), .A2(n143gat) );
  OR3_X1 OR3_50( .ZN(n2916gat), .A1(n971gat), .A2(n970gat), .A3(n968gat) );
  OR3_X1 OR3_51( .ZN(n2875gat), .A1(n142gat), .A2(n40gat), .A3(n39gat) );
  OR3_X1 OR3_52( .ZN(n2899gat), .A1(n772gat), .A2(n451gat), .A3(n446gat) );
  OR2_X1 OR2_75( .ZN(n2877gat), .A1(n139gat), .A2(n136gat) );
  OR2_X1 OR2_76( .ZN(n2893gat), .A1(n391gat), .A2(n390gat) );
  OR2_X1 OR2_77( .ZN(n2926gat), .A1(n1083gat), .A2(n1077gat) );
  OR2_X1 OR2_78( .ZN(n2882gat), .A1(n242gat), .A2(n240gat) );
  OR2_X1 OR2_79( .ZN(n2924gat), .A1(n871gat), .A2(n797gat) );
  OR3_X1 OR3_53( .ZN(n2881gat), .A1(n324gat), .A2(n238gat), .A3(n237gat) );
  OR2_X1 OR2_80( .ZN(n2923gat), .A1(n1082gat), .A2(n796gat) );
  OR2_X1 OR2_81( .ZN(n2710gat), .A1(n69gat), .A2(n1885gat) );
  OR2_X1 OR2_82( .ZN(n2704gat), .A1(n11gat), .A2(n1889gat) );
  OR2_X1 OR2_83( .ZN(n2684gat), .A1(n1599gat), .A2(n2051gat) );
  OR2_X1 OR2_84( .ZN(n2830gat), .A1(n2444gat), .A2(n1754gat) );
  OR3_X1 OR3_54( .ZN(II3999), .A1(n2167gat), .A2(n2031gat), .A3(n2174gat) );
  OR4_X1 OR4_38( .ZN(II4000), .A1(n2108gat), .A2(n2093gat), .A3(n2035gat), .A4(II3999) );
  OR2_X1 OR2_85( .ZN(n2695gat), .A1(n1586gat), .A2(n1791gat) );
  OR2_X1 OR2_86( .ZN(n2703gat), .A1(n1755gat), .A2(n1518gat) );
  OR2_X1 OR2_87( .ZN(n2744gat), .A1(n2159gat), .A2(n2478gat) );
  OR2_X1 OR2_88( .ZN(n2800gat), .A1(n2158gat), .A2(n2186gat) );
  OR3_X1 OR3_55( .ZN(II4023), .A1(n2443gat), .A2(n2290gat), .A3(n2214gat) );
  OR3_X1 OR3_56( .ZN(II4024), .A1(n2353gat), .A2(n2284gat), .A3(II4023) );
  OR4_X2 OR4_39( .ZN(n2980gat), .A1(n1470gat), .A2(n1400gat), .A3(n1399gat), .A4(n1398gat) );
  OR3_X1 OR3_57( .ZN(II4144), .A1(n1633gat), .A2(n1838gat), .A3(n1786gat) );
  OR3_X1 OR3_58( .ZN(II4145), .A1(n1788gat), .A2(n1784gat), .A3(II4144) );
  OR2_X1 OR2_89( .ZN(n2984gat), .A1(n1467gat), .A2(n1466gat) );
  OR4_X1 OR4_40( .ZN(n2985gat), .A1(n1686gat), .A2(n1533gat), .A3(n1532gat), .A4(n1531gat) );
  OR3_X1 OR3_59( .ZN(II4216), .A1(n1427gat), .A2(n1595gat), .A3(n1677gat) );
  OR3_X1 OR3_60( .ZN(II4217), .A1(n1392gat), .A2(n2989gat), .A3(II4216) );
  OR4_X1 OR4_41( .ZN(n2931gat), .A1(n1100gat), .A2(n994gat), .A3(n989gat), .A4(n880gat) );
  OR2_X1 OR2_90( .ZN(n2943gat), .A1(n1012gat), .A2(n905gat) );
  OR2_X1 OR2_91( .ZN(n2941gat), .A1(n1003gat), .A2(n902gat) );
  OR4_X1 OR4_42( .ZN(n2946gat), .A1(n1099gat), .A2(n998gat), .A3(n995gat), .A4(n980gat) );
  OR2_X1 OR2_92( .ZN(n2960gat), .A1(n1175gat), .A2(n1174gat) );
  OR2_X1 OR2_93( .ZN(n2950gat), .A1(n1001gat), .A2(n999gat) );
  OR2_X1 OR2_94( .ZN(n2969gat), .A1(n1323gat), .A2(n1264gat) );
  OR4_X1 OR4_43( .ZN(n2933gat), .A1(n981gat), .A2(n890gat), .A3(n889gat), .A4(n886gat) );
  OR2_X1 OR2_95( .ZN(n2935gat), .A1(n892gat), .A2(n891gat) );
  OR2_X2 OR2_96( .ZN(n2942gat), .A1(n904gat), .A2(n903gat) );
  OR4_X1 OR4_44( .ZN(n2940gat), .A1(n1152gat), .A2(n1092gat), .A3(n997gat), .A4(n993gat) );
  OR2_X1 OR2_97( .ZN(n2937gat), .A1(n900gat), .A2(n895gat) );
  OR4_X1 OR4_45( .ZN(n2947gat), .A1(n1094gat), .A2(n1093gat), .A3(n988gat), .A4(n984gat) );
  OR2_X1 OR2_98( .ZN(n2965gat), .A1(n1267gat), .A2(n1257gat) );
  OR2_X1 OR2_99( .ZN(n2956gat), .A1(n1178gat), .A2(n1116gat) );
  OR2_X1 OR2_100( .ZN(n2961gat), .A1(n1375gat), .A2(n1324gat) );
  OR4_X1 OR4_46( .ZN(n2939gat), .A1(n1091gat), .A2(n1088gat), .A3(n992gat), .A4(n987gat) );
  OR2_X1 OR2_101( .ZN(n2938gat), .A1(n899gat), .A2(n896gat) );
  OR2_X1 OR2_102( .ZN(n2967gat), .A1(n1262gat), .A2(n1260gat) );
  OR4_X1 OR4_47( .ZN(n2932gat), .A1(n1098gat), .A2(n1090gat), .A3(n986gat), .A4(n885gat) );
  OR2_X1 OR2_103( .ZN(n2936gat), .A1(n901gat), .A2(n893gat) );
  OR4_X1 OR4_48( .ZN(n2948gat), .A1(n1097gat), .A2(n1089gat), .A3(n1087gat), .A4(n991gat) );
  OR2_X1 OR2_104( .ZN(n2968gat), .A1(n1326gat), .A2(n1261gat) );
  OR2_X1 OR2_105( .ZN(n2955gat), .A1(n1177gat), .A2(n1115gat) );
  OR2_X1 OR2_106( .ZN(n2944gat), .A1(n977gat), .A2(n976gat) );
  OR4_X1 OR4_49( .ZN(n2945gat), .A1(n1096gat), .A2(n1095gat), .A3(n990gat), .A4(n979gat) );
  OR2_X1 OR2_107( .ZN(n2962gat), .A1(n1176gat), .A2(n1173gat) );
  OR2_X1 OR2_108( .ZN(n2951gat), .A1(n1004gat), .A2(n1000gat) );
  OR2_X1 OR2_109( .ZN(n2764gat), .A1(n1029gat), .A2(n2237gat) );
  OR2_X1 OR2_110( .ZN(n2762gat), .A1(n1028gat), .A2(n1782gat) );
  OR2_X1 OR2_111( .ZN(n2761gat), .A1(n1031gat), .A2(n2325gat) );
  OR2_X1 OR2_112( .ZN(n2757gat), .A1(n1030gat), .A2(n2245gat) );
  OR2_X1 OR2_113( .ZN(n2756gat), .A1(n1011gat), .A2(n2244gat) );
  OR2_X1 OR2_114( .ZN(n2750gat), .A1(n1181gat), .A2(n2243gat) );
  OR2_X1 OR2_115( .ZN(n2749gat), .A1(n1010gat), .A2(n2246gat) );
  OR2_X1 OR2_116( .ZN(n2742gat), .A1(n1005gat), .A2(n2384gat) );
  OR2_X1 OR2_117( .ZN(n2741gat), .A1(n1182gat), .A2(n2385gat) );
  OR2_X1 OR2_118( .ZN(n2694gat), .A1(n1381gat), .A2(n1384gat) );
  OR2_X1 OR2_119( .ZN(n2693gat), .A1(n1451gat), .A2(n1453gat) );
  OR2_X1 OR2_120( .ZN(n2702gat), .A1(n925gat), .A2(n1452gat) );
  OR2_X1 OR2_121( .ZN(n2701gat), .A1(n921gat), .A2(n1890gat) );
  OR2_X1 OR2_122( .ZN(n2709gat), .A1(n739gat), .A2(n1841gat) );
  OR2_X1 OR2_123( .ZN(n2708gat), .A1(n848gat), .A2(n2047gat) );
  OR2_X2 OR2_124( .ZN(n2799gat), .A1(n849gat), .A2(n2050gat) );
  OR2_X1 OR2_125( .ZN(n2798gat), .A1(n1032gat), .A2(n2054gat) );
  OR3_X1 OR3_61( .ZN(n2812gat), .A1(n73gat), .A2(n70gat), .A3(n1840gat) );
  OR3_X1 OR3_62( .ZN(n2822gat), .A1(n77gat), .A2(n13gat), .A3(n1842gat) );
  NOR2_X1 NOR2_0( .ZN(n421gat), .A1(n2715gat), .A2(n2723gat) );
  NOR2_X1 NOR2_1( .ZN(n648gat), .A1(n373gat), .A2(n2669gat) );
  NOR2_X1 NOR2_2( .ZN(n442gat), .A1(n2844gat), .A2(n856gat) );
  NOR2_X1 NOR2_3( .ZN(n1499gat), .A1(n396gat), .A2(n401gat) );
  NOR2_X1 NOR2_4( .ZN(n1616gat), .A1(n918gat), .A2(n396gat) );
  NOR2_X2 NOR2_5( .ZN(n1614gat), .A1(n396gat), .A2(n845gat) );
  NOR3_X1 NOR3_0( .ZN(n1641gat), .A1(n1645gat), .A2(n1553gat), .A3(n1559gat) );
  NOR3_X1 NOR3_1( .ZN(n1642gat), .A1(n1559gat), .A2(n1616gat), .A3(n1645gat) );
  NOR3_X1 NOR3_2( .ZN(n1556gat), .A1(n1614gat), .A2(n1645gat), .A3(n1616gat) );
  NOR3_X1 NOR3_3( .ZN(n1557gat), .A1(n1553gat), .A2(n1645gat), .A3(n1614gat) );
  NOR3_X1 NOR3_4( .ZN(n1639gat), .A1(n1499gat), .A2(n1559gat), .A3(n1553gat) );
  NOR3_X1 NOR4_0_A( .ZN(extra0), .A1(n1614gat), .A2(n1616gat), .A3(n1499gat) );
  NOR2_X1 NOR4_0( .ZN(n1605gat), .A1(extra0), .A2(n396gat) );
  NOR3_X1 NOR3_5( .ZN(n1555gat), .A1(n1616gat), .A2(n1559gat), .A3(n1499gat) );
  NOR3_X1 NOR3_6( .ZN(n1558gat), .A1(n1614gat), .A2(n1553gat), .A3(n1499gat) );
  NOR2_X1 NOR2_6( .ZN(n1256gat), .A1(n392gat), .A2(n702gat) );
  NOR2_X1 NOR2_7( .ZN(n1117gat), .A1(n720gat), .A2(n725gat) );
  NOR2_X1 NOR2_8( .ZN(n1618gat), .A1(n1319gat), .A2(n1447gat) );
  NOR2_X1 NOR2_9( .ZN(n1114gat), .A1(n725gat), .A2(n721gat) );
  NOR2_X2 NOR2_10( .ZN(n1621gat), .A1(n1319gat), .A2(n1380gat) );
  NOR2_X1 NOR2_11( .ZN(n1318gat), .A1(n392gat), .A2(n701gat) );
  NOR2_X1 NOR2_12( .ZN(n1619gat), .A1(n1447gat), .A2(n1446gat) );
  NOR2_X1 NOR2_13( .ZN(n1622gat), .A1(n1380gat), .A2(n1446gat) );
  NOR3_X1 NOR3_7( .ZN(n1214gat), .A1(n1218gat), .A2(n1219gat), .A3(n1220gat) );
  NOR3_X1 NOR3_8( .ZN(n1215gat), .A1(n1218gat), .A2(n1221gat), .A3(n1222gat) );
  NOR3_X1 NOR3_9( .ZN(n1216gat), .A1(n1223gat), .A2(n1219gat), .A3(n1222gat) );
  NOR3_X1 NOR3_10( .ZN(n1217gat), .A1(n1223gat), .A2(n1221gat), .A3(n1220gat) );
  NOR2_X1 NOR2_14( .ZN(n745gat), .A1(n2716gat), .A2(n2867gat) );
  NOR2_X1 NOR2_15( .ZN(n638gat), .A1(n2715gat), .A2(n2868gat) );
  NOR2_X1 NOR2_16( .ZN(n423gat), .A1(n2724gat), .A2(n2726gat) );
  NOR2_X1 NOR2_17( .ZN(n362gat), .A1(n2723gat), .A2(n2727gat) );
  NOR3_X1 NOR3_11( .ZN(n749gat), .A1(n753gat), .A2(n754gat), .A3(n755gat) );
  NOR3_X1 NOR3_12( .ZN(n750gat), .A1(n753gat), .A2(n756gat), .A3(n757gat) );
  NOR3_X1 NOR3_13( .ZN(n751gat), .A1(n758gat), .A2(n754gat), .A3(n757gat) );
  NOR3_X1 NOR3_14( .ZN(n752gat), .A1(n758gat), .A2(n756gat), .A3(n755gat) );
  NOR3_X1 NOR3_15( .ZN(n259gat), .A1(n263gat), .A2(n264gat), .A3(n265gat) );
  NOR3_X2 NOR3_16( .ZN(n260gat), .A1(n263gat), .A2(n266gat), .A3(n267gat) );
  NOR3_X1 NOR3_17( .ZN(n261gat), .A1(n268gat), .A2(n264gat), .A3(n267gat) );
  NOR3_X1 NOR3_18( .ZN(n262gat), .A1(n268gat), .A2(n266gat), .A3(n265gat) );
  NOR3_X1 NOR3_19( .ZN(n1014gat), .A1(n1018gat), .A2(n1019gat), .A3(n1020gat) );
  NOR3_X1 NOR3_20( .ZN(n1015gat), .A1(n1018gat), .A2(n1021gat), .A3(n1022gat) );
  NOR3_X1 NOR3_21( .ZN(n1016gat), .A1(n1023gat), .A2(n1019gat), .A3(n1022gat) );
  NOR3_X1 NOR3_22( .ZN(n1017gat), .A1(n1023gat), .A2(n1021gat), .A3(n1020gat) );
  NOR3_X1 NOR3_23( .ZN(n476gat), .A1(n480gat), .A2(n481gat), .A3(n482gat) );
  NOR3_X1 NOR3_24( .ZN(n477gat), .A1(n480gat), .A2(n483gat), .A3(n484gat) );
  NOR3_X1 NOR3_25( .ZN(n478gat), .A1(n485gat), .A2(n481gat), .A3(n484gat) );
  NOR3_X1 NOR3_26( .ZN(n479gat), .A1(n485gat), .A2(n483gat), .A3(n482gat) );
  NOR3_X1 NOR3_27( .ZN(n44gat), .A1(n48gat), .A2(n49gat), .A3(n50gat) );
  NOR3_X1 NOR3_28( .ZN(n45gat), .A1(n48gat), .A2(n51gat), .A3(n52gat) );
  NOR3_X1 NOR3_29( .ZN(n46gat), .A1(n53gat), .A2(n49gat), .A3(n52gat) );
  NOR3_X2 NOR3_30( .ZN(n47gat), .A1(n53gat), .A2(n51gat), .A3(n50gat) );
  NOR2_X1 NOR2_18( .ZN(n1376gat), .A1(n724gat), .A2(n720gat) );
  NOR2_X1 NOR2_19( .ZN(n1617gat), .A1(n1319gat), .A2(n1448gat) );
  NOR2_X1 NOR2_20( .ZN(n1377gat), .A1(n724gat), .A2(n721gat) );
  NOR2_X1 NOR2_21( .ZN(n1624gat), .A1(n1319gat), .A2(n1379gat) );
  NOR2_X1 NOR2_22( .ZN(n1113gat), .A1(n393gat), .A2(n701gat) );
  NOR2_X1 NOR2_23( .ZN(n1501gat), .A1(n1448gat), .A2(n1500gat) );
  NOR2_X1 NOR2_24( .ZN(n1623gat), .A1(n1379gat), .A2(n1446gat) );
  NOR2_X1 NOR2_25( .ZN(n1620gat), .A1(n1448gat), .A2(n1446gat) );
  NOR2_X1 NOR2_26( .ZN(n1827gat), .A1(n2729gat), .A2(n2317gat) );
  NOR2_X1 NOR2_27( .ZN(n1817gat), .A1(n1819gat), .A2(n1823gat) );
  NOR2_X1 NOR2_28( .ZN(n1935gat), .A1(n1816gat), .A2(n1828gat) );
  NOR2_X1 NOR2_29( .ZN(n529gat), .A1(n2724gat), .A2(n2715gat) );
  NOR2_X1 NOR2_30( .ZN(n361gat), .A1(n2859gat), .A2(n2726gat) );
  NOR3_X1 NOR3_31( .ZN(n168gat), .A1(n172gat), .A2(n173gat), .A3(n174gat) );
  NOR3_X1 NOR3_32( .ZN(n169gat), .A1(n172gat), .A2(n175gat), .A3(n176gat) );
  NOR3_X1 NOR3_33( .ZN(n170gat), .A1(n177gat), .A2(n173gat), .A3(n176gat) );
  NOR3_X1 NOR3_34( .ZN(n171gat), .A1(n177gat), .A2(n175gat), .A3(n174gat) );
  NOR3_X1 NOR3_35( .ZN(n907gat), .A1(n911gat), .A2(n912gat), .A3(n913gat) );
  NOR3_X2 NOR3_36( .ZN(n908gat), .A1(n911gat), .A2(n914gat), .A3(n915gat) );
  NOR3_X1 NOR3_37( .ZN(n909gat), .A1(n916gat), .A2(n912gat), .A3(n915gat) );
  NOR3_X1 NOR3_38( .ZN(n910gat), .A1(n916gat), .A2(n914gat), .A3(n913gat) );
  NOR3_X1 NOR3_39( .ZN(n344gat), .A1(n348gat), .A2(n349gat), .A3(n350gat) );
  NOR3_X1 NOR3_40( .ZN(n345gat), .A1(n348gat), .A2(n351gat), .A3(n352gat) );
  NOR3_X1 NOR3_41( .ZN(n346gat), .A1(n353gat), .A2(n349gat), .A3(n352gat) );
  NOR3_X1 NOR3_42( .ZN(n347gat), .A1(n353gat), .A2(n351gat), .A3(n350gat) );
  NOR3_X1 NOR3_43( .ZN(n56gat), .A1(n60gat), .A2(n61gat), .A3(n62gat) );
  NOR3_X1 NOR3_44( .ZN(n57gat), .A1(n60gat), .A2(n63gat), .A3(n64gat) );
  NOR3_X1 NOR3_45( .ZN(n58gat), .A1(n65gat), .A2(n61gat), .A3(n64gat) );
  NOR3_X1 NOR3_46( .ZN(n59gat), .A1(n65gat), .A2(n63gat), .A3(n62gat) );
  NOR2_X1 NOR2_31( .ZN(n768gat), .A1(n373gat), .A2(n2731gat) );
  NOR2_X1 NOR2_32( .ZN(n655gat), .A1(n856gat), .A2(n2718gat) );
  NOR2_X1 NOR2_33( .ZN(n963gat), .A1(n856gat), .A2(n2838gat) );
  NOR2_X1 NOR2_34( .ZN(n868gat), .A1(n2775gat), .A2(n373gat) );
  NOR2_X1 NOR2_35( .ZN(n962gat), .A1(n856gat), .A2(n2711gat) );
  NOR2_X1 NOR2_36( .ZN(n959gat), .A1(n373gat), .A2(n2734gat) );
  NOR3_X2 NOR3_47( .ZN(n945gat), .A1(n949gat), .A2(n950gat), .A3(n951gat) );
  NOR3_X1 NOR3_48( .ZN(n946gat), .A1(n949gat), .A2(n952gat), .A3(n953gat) );
  NOR3_X1 NOR3_49( .ZN(n947gat), .A1(n954gat), .A2(n950gat), .A3(n953gat) );
  NOR3_X1 NOR3_50( .ZN(n948gat), .A1(n954gat), .A2(n952gat), .A3(n951gat) );
  NOR2_X1 NOR2_37( .ZN(n647gat), .A1(n2792gat), .A2(n373gat) );
  NOR2_X1 NOR2_38( .ZN(n441gat), .A1(n856gat), .A2(n2846gat) );
  NOR2_X1 NOR2_39( .ZN(n967gat), .A1(n373gat), .A2(n2672gat) );
  NOR2_X1 NOR2_40( .ZN(n792gat), .A1(n2852gat), .A2(n856gat) );
  NOR3_X1 NOR3_51( .ZN(n1229gat), .A1(n1233gat), .A2(n1234gat), .A3(n1235gat) );
  NOR3_X1 NOR3_52( .ZN(n1230gat), .A1(n1233gat), .A2(n1236gat), .A3(n1237gat) );
  NOR3_X1 NOR3_53( .ZN(n1231gat), .A1(n1238gat), .A2(n1234gat), .A3(n1237gat) );
  NOR3_X1 NOR3_54( .ZN(n1232gat), .A1(n1238gat), .A2(n1236gat), .A3(n1235gat) );
  NOR2_X1 NOR2_41( .ZN(n443gat), .A1(n2778gat), .A2(n373gat) );
  NOR2_X1 NOR2_42( .ZN(n439gat), .A1(n856gat), .A2(n2836gat) );
  NOR2_X1 NOR2_43( .ZN(n966gat), .A1(n2789gat), .A2(n373gat) );
  NOR2_X1 NOR2_44( .ZN(n790gat), .A1(n856gat), .A2(n2840gat) );
  NOR2_X1 NOR2_45( .ZN(n444gat), .A1(n373gat), .A2(n2781gat) );
  NOR2_X2 NOR2_46( .ZN(n440gat), .A1(n856gat), .A2(n2842gat) );
  NOR3_X1 NOR3_55( .ZN(n1051gat), .A1(n1055gat), .A2(n1056gat), .A3(n1057gat) );
  NOR3_X1 NOR3_56( .ZN(n1052gat), .A1(n1055gat), .A2(n1058gat), .A3(n1059gat) );
  NOR3_X1 NOR3_57( .ZN(n1053gat), .A1(n1060gat), .A2(n1056gat), .A3(n1059gat) );
  NOR3_X1 NOR3_58( .ZN(n1054gat), .A1(n1060gat), .A2(n1058gat), .A3(n1057gat) );
  NOR3_X1 NOR3_59( .ZN(n934gat), .A1(n938gat), .A2(n939gat), .A3(n940gat) );
  NOR3_X1 NOR3_60( .ZN(n935gat), .A1(n938gat), .A2(n941gat), .A3(n942gat) );
  NOR3_X1 NOR3_61( .ZN(n936gat), .A1(n943gat), .A2(n939gat), .A3(n942gat) );
  NOR3_X1 NOR3_62( .ZN(n937gat), .A1(n943gat), .A2(n941gat), .A3(n940gat) );
  NOR2_X1 NOR2_47( .ZN(n746gat), .A1(n2716gat), .A2(n2723gat) );
  NOR2_X1 NOR2_48( .ZN(n360gat), .A1(n2859gat), .A2(n2727gat) );
  NOR3_X1 NOR3_63( .ZN(n710gat), .A1(n714gat), .A2(n715gat), .A3(n716gat) );
  NOR3_X1 NOR3_64( .ZN(n711gat), .A1(n714gat), .A2(n717gat), .A3(n718gat) );
  NOR3_X1 NOR3_65( .ZN(n712gat), .A1(n719gat), .A2(n715gat), .A3(n718gat) );
  NOR3_X1 NOR3_66( .ZN(n713gat), .A1(n719gat), .A2(n717gat), .A3(n716gat) );
  NOR3_X1 NOR3_67( .ZN(n729gat), .A1(n733gat), .A2(n734gat), .A3(n735gat) );
  NOR3_X1 NOR3_68( .ZN(n730gat), .A1(n733gat), .A2(n736gat), .A3(n737gat) );
  NOR3_X1 NOR3_69( .ZN(n731gat), .A1(n738gat), .A2(n734gat), .A3(n737gat) );
  NOR3_X1 NOR3_70( .ZN(n732gat), .A1(n738gat), .A2(n736gat), .A3(n735gat) );
  NOR3_X1 NOR3_71( .ZN(n494gat), .A1(n498gat), .A2(n499gat), .A3(n500gat) );
  NOR3_X1 NOR3_72( .ZN(n495gat), .A1(n498gat), .A2(n501gat), .A3(n502gat) );
  NOR3_X1 NOR3_73( .ZN(n496gat), .A1(n503gat), .A2(n499gat), .A3(n502gat) );
  NOR3_X1 NOR3_74( .ZN(n497gat), .A1(n503gat), .A2(n501gat), .A3(n500gat) );
  NOR3_X1 NOR3_75( .ZN(n505gat), .A1(n509gat), .A2(n510gat), .A3(n511gat) );
  NOR3_X1 NOR3_76( .ZN(n506gat), .A1(n509gat), .A2(n512gat), .A3(n513gat) );
  NOR3_X1 NOR3_77( .ZN(n507gat), .A1(n514gat), .A2(n510gat), .A3(n513gat) );
  NOR3_X1 NOR3_78( .ZN(n508gat), .A1(n514gat), .A2(n512gat), .A3(n511gat) );
  NOR3_X1 NOR4_1_A( .ZN(extra1), .A1(n3029gat), .A2(n2863gat), .A3(n2855gat) );
  NOR2_X1 NOR4_1( .ZN(n564gat), .A1(extra1), .A2(n374gat) );
  NOR3_X2 NOR3_79( .ZN(n86gat), .A1(n743gat), .A2(n294gat), .A3(n17gat) );
  NOR2_X1 NOR2_49( .ZN(n78gat), .A1(n2784gat), .A2(n79gat) );
  NOR2_X1 NOR2_50( .ZN(n767gat), .A1(n219gat), .A2(n2731gat) );
  NOR2_X1 NOR2_51( .ZN(n286gat), .A1(n289gat), .A2(n2723gat) );
  NOR2_X1 NOR2_52( .ZN(n287gat), .A1(n289gat), .A2(n2715gat) );
  NOR2_X1 NOR2_53( .ZN(n288gat), .A1(n289gat), .A2(n2726gat) );
  NOR3_X1 NOR3_80( .ZN(n181gat), .A1(n286gat), .A2(n179gat), .A3(n188gat) );
  NOR2_X1 NOR2_54( .ZN(n182gat), .A1(n72gat), .A2(n2720gat) );
  NOR2_X1 NOR2_55( .ZN(n653gat), .A1(n2718gat), .A2(n111gat) );
  NOR2_X1 NOR2_56( .ZN(n867gat), .A1(n219gat), .A2(n2775gat) );
  NOR2_X2 NOR2_57( .ZN(n771gat), .A1(n2838gat), .A2(n111gat) );
  NOR2_X1 NOR2_58( .ZN(n964gat), .A1(n111gat), .A2(n2711gat) );
  NOR2_X1 NOR2_59( .ZN(n961gat), .A1(n219gat), .A2(n2734gat) );
  NOR3_X1 NOR3_81( .ZN(n804gat), .A1(n808gat), .A2(n809gat), .A3(n810gat) );
  NOR3_X1 NOR3_82( .ZN(n805gat), .A1(n808gat), .A2(n811gat), .A3(n812gat) );
  NOR3_X1 NOR3_83( .ZN(n806gat), .A1(n813gat), .A2(n809gat), .A3(n812gat) );
  NOR3_X1 NOR3_84( .ZN(n807gat), .A1(n813gat), .A2(n811gat), .A3(n810gat) );
  NOR3_X1 NOR3_85( .ZN(n587gat), .A1(n591gat), .A2(n592gat), .A3(n593gat) );
  NOR3_X1 NOR3_86( .ZN(n588gat), .A1(n591gat), .A2(n594gat), .A3(n595gat) );
  NOR3_X1 NOR3_87( .ZN(n589gat), .A1(n596gat), .A2(n592gat), .A3(n595gat) );
  NOR3_X1 NOR3_88( .ZN(n590gat), .A1(n596gat), .A2(n594gat), .A3(n593gat) );
  NOR2_X1 NOR2_60( .ZN(n447gat), .A1(n2836gat), .A2(n111gat) );
  NOR2_X1 NOR2_61( .ZN(n445gat), .A1(n2778gat), .A2(n219gat) );
  NOR3_X1 NOR3_89( .ZN(n687gat), .A1(n691gat), .A2(n692gat), .A3(n693gat) );
  NOR3_X1 NOR3_90( .ZN(n688gat), .A1(n691gat), .A2(n694gat), .A3(n695gat) );
  NOR3_X1 NOR3_91( .ZN(n689gat), .A1(n696gat), .A2(n692gat), .A3(n695gat) );
  NOR3_X1 NOR3_92( .ZN(n690gat), .A1(n696gat), .A2(n694gat), .A3(n693gat) );
  NOR3_X1 NOR3_93( .ZN(n568gat), .A1(n572gat), .A2(n573gat), .A3(n574gat) );
  NOR3_X1 NOR3_94( .ZN(n569gat), .A1(n572gat), .A2(n575gat), .A3(n576gat) );
  NOR3_X1 NOR3_95( .ZN(n570gat), .A1(n577gat), .A2(n573gat), .A3(n576gat) );
  NOR3_X1 NOR3_96( .ZN(n571gat), .A1(n577gat), .A2(n575gat), .A3(n574gat) );
  NOR3_X1 NOR3_97( .ZN(n187gat), .A1(n189gat), .A2(n287gat), .A3(n188gat) );
  NOR2_X1 NOR2_62( .ZN(n197gat), .A1(n194gat), .A2(n297gat) );
  NOR3_X1 NOR3_98( .ZN(n15gat), .A1(n637gat), .A2(n17gat), .A3(n293gat) );
  NOR2_X2 NOR2_63( .ZN(n22gat), .A1(n92gat), .A2(n21gat) );
  NOR2_X1 NOR2_64( .ZN(n93gat), .A1(n197gat), .A2(n22gat) );
  NOR2_X1 NOR2_65( .ZN(n769gat), .A1(n93gat), .A2(n2731gat) );
  NOR3_X1 NOR3_99( .ZN(n2534gat), .A1(n2624gat), .A2(n2489gat), .A3(n2621gat) );
  NOR3_X1 NOR3_100( .ZN(n2430gat), .A1(n2533gat), .A2(n2486gat), .A3(n2429gat) );
  NOR2_X1 NOR2_66( .ZN(n1606gat), .A1(n3020gat), .A2(n270gat) );
  NOR2_X1 NOR2_67( .ZN(n2239gat), .A1(n2850gat), .A2(n3019gat) );
  NOR3_X1 NOR3_101( .ZN(n1934gat), .A1(n2470gat), .A2(n1935gat), .A3(n2239gat) );
  NOR2_X1 NOR2_68( .ZN(n1610gat), .A1(n1698gat), .A2(n1543gat) );
  NOR2_X1 NOR2_69( .ZN(n1692gat), .A1(n1879gat), .A2(n1762gat) );
  NOR2_X1 NOR2_70( .ZN(n2433gat), .A1(n2432gat), .A2(n2154gat) );
  NOR3_X1 NOR3_102( .ZN(n2531gat), .A1(n2488gat), .A2(n2625gat), .A3(n2621gat) );
  NOR3_X1 NOR3_103( .ZN(n2480gat), .A1(n2530gat), .A2(n2482gat), .A3(n2486gat) );
  NOR2_X1 NOR2_71( .ZN(n2427gat), .A1(n2426gat), .A2(n2153gat) );
  NOR2_X1 NOR2_72( .ZN(n2428gat), .A1(n2433gat), .A2(n2427gat) );
  NOR2_X1 NOR2_73( .ZN(n1778gat), .A1(n3026gat), .A2(n1779gat) );
  NOR2_X2 NOR2_74( .ZN(n1609gat), .A1(n1503gat), .A2(n3025gat) );
  NOR2_X1 NOR2_75( .ZN(n1702gat), .A1(n3024gat), .A2(n1615gat) );
  NOR2_X1 NOR2_76( .ZN(n1700gat), .A1(n1701gat), .A2(n3023gat) );
  NOR3_X1 NOR4_2_A( .ZN(extra2), .A1(n1778gat), .A2(n1609gat), .A3(n1702gat) );
  NOR2_X1 NOR4_2( .ZN(n1604gat), .A1(extra2), .A2(n1700gat) );
  NOR2_X1 NOR2_77( .ZN(n1076gat), .A1(n93gat), .A2(n2775gat) );
  NOR2_X1 NOR2_78( .ZN(n766gat), .A1(n93gat), .A2(n2734gat) );
  NOR3_X1 NOR3_104( .ZN(n1185gat), .A1(n1189gat), .A2(n1190gat), .A3(n1191gat) );
  NOR3_X1 NOR3_105( .ZN(n1186gat), .A1(n1189gat), .A2(n1192gat), .A3(n1193gat) );
  NOR3_X1 NOR3_106( .ZN(n1187gat), .A1(n1194gat), .A2(n1190gat), .A3(n1193gat) );
  NOR3_X1 NOR3_107( .ZN(n1188gat), .A1(n1194gat), .A2(n1192gat), .A3(n1191gat) );
  NOR2_X1 NOR2_79( .ZN(n645gat), .A1(n2792gat), .A2(n93gat) );
  NOR2_X1 NOR2_80( .ZN(n646gat), .A1(n93gat), .A2(n2669gat) );
  NOR2_X1 NOR2_81( .ZN(n1383gat), .A1(n1280gat), .A2(n1225gat) );
  NOR2_X1 NOR2_82( .ZN(n1327gat), .A1(n1281gat), .A2(n1224gat) );
  NOR2_X1 NOR2_83( .ZN(n651gat), .A1(n93gat), .A2(n2778gat) );
  NOR2_X1 NOR2_84( .ZN(n652gat), .A1(n2789gat), .A2(n93gat) );
  NOR2_X1 NOR2_85( .ZN(n765gat), .A1(n2781gat), .A2(n93gat) );
  NOR3_X1 NOR3_108( .ZN(n1202gat), .A1(n1206gat), .A2(n1207gat), .A3(n1208gat) );
  NOR3_X1 NOR3_109( .ZN(n1203gat), .A1(n1206gat), .A2(n1209gat), .A3(n1210gat) );
  NOR3_X1 NOR3_110( .ZN(n1204gat), .A1(n1211gat), .A2(n1207gat), .A3(n1210gat) );
  NOR3_X1 NOR3_111( .ZN(n1205gat), .A1(n1211gat), .A2(n1209gat), .A3(n1208gat) );
  NOR3_X1 NOR3_112( .ZN(n1270gat), .A1(n1274gat), .A2(n1275gat), .A3(n1276gat) );
  NOR3_X2 NOR3_113( .ZN(n1271gat), .A1(n1274gat), .A2(n1277gat), .A3(n1278gat) );
  NOR3_X1 NOR3_114( .ZN(n1272gat), .A1(n1279gat), .A2(n1275gat), .A3(n1278gat) );
  NOR3_X1 NOR3_115( .ZN(n1273gat), .A1(n1279gat), .A2(n1277gat), .A3(n1276gat) );
  NOR2_X1 NOR2_86( .ZN(n763gat), .A1(n2672gat), .A2(n93gat) );
  NOR2_X1 NOR2_87( .ZN(n1287gat), .A1(n1284gat), .A2(n1195gat) );
  NOR2_X1 NOR2_88( .ZN(n1285gat), .A1(n1196gat), .A2(n1269gat) );
  NOR2_X1 NOR2_89( .ZN(n853gat), .A1(n740gat), .A2(n2148gat) );
  NOR2_X1 NOR2_90( .ZN(n793gat), .A1(n2852gat), .A2(n851gat) );
  NOR2_X1 NOR2_91( .ZN(n854gat), .A1(n2148gat), .A2(n374gat) );
  NOR2_X1 NOR2_92( .ZN(n556gat), .A1(n2672gat), .A2(n852gat) );
  NOR2_X1 NOR2_93( .ZN(n795gat), .A1(n2731gat), .A2(n852gat) );
  NOR2_X1 NOR2_94( .ZN(n656gat), .A1(n851gat), .A2(n2718gat) );
  NOR2_X2 NOR2_95( .ZN(n794gat), .A1(n852gat), .A2(n2775gat) );
  NOR2_X1 NOR2_96( .ZN(n773gat), .A1(n851gat), .A2(n2838gat) );
  NOR2_X1 NOR2_97( .ZN(n965gat), .A1(n2711gat), .A2(n851gat) );
  NOR2_X1 NOR2_98( .ZN(n960gat), .A1(n2734gat), .A2(n852gat) );
  NOR3_X1 NOR3_116( .ZN(n780gat), .A1(n784gat), .A2(n785gat), .A3(n786gat) );
  NOR3_X1 NOR3_117( .ZN(n781gat), .A1(n784gat), .A2(n787gat), .A3(n788gat) );
  NOR3_X1 NOR3_118( .ZN(n782gat), .A1(n789gat), .A2(n785gat), .A3(n788gat) );
  NOR3_X1 NOR3_119( .ZN(n783gat), .A1(n789gat), .A2(n787gat), .A3(n786gat) );
  NOR2_X1 NOR2_99( .ZN(n555gat), .A1(n852gat), .A2(n2792gat) );
  NOR2_X1 NOR2_100( .ZN(n450gat), .A1(n851gat), .A2(n2846gat) );
  NOR2_X1 NOR2_101( .ZN(n654gat), .A1(n851gat), .A2(n2844gat) );
  NOR2_X1 NOR2_102( .ZN(n557gat), .A1(n2669gat), .A2(n852gat) );
  NOR2_X1 NOR2_103( .ZN(n874gat), .A1(n559gat), .A2(n365gat) );
  NOR2_X1 NOR2_104( .ZN(n132gat), .A1(n560gat), .A2(n364gat) );
  NOR2_X1 NOR2_105( .ZN(n649gat), .A1(n2778gat), .A2(n852gat) );
  NOR2_X1 NOR2_106( .ZN(n449gat), .A1(n2836gat), .A2(n851gat) );
  NOR2_X1 NOR2_107( .ZN(n791gat), .A1(n851gat), .A2(n2840gat) );
  NOR2_X1 NOR2_108( .ZN(n650gat), .A1(n852gat), .A2(n2789gat) );
  NOR2_X1 NOR2_109( .ZN(n774gat), .A1(n2842gat), .A2(n851gat) );
  NOR2_X1 NOR2_110( .ZN(n764gat), .A1(n852gat), .A2(n2781gat) );
  NOR3_X1 NOR3_120( .ZN(n222gat), .A1(n226gat), .A2(n227gat), .A3(n228gat) );
  NOR3_X2 NOR3_121( .ZN(n223gat), .A1(n226gat), .A2(n229gat), .A3(n230gat) );
  NOR3_X1 NOR3_122( .ZN(n224gat), .A1(n231gat), .A2(n227gat), .A3(n230gat) );
  NOR3_X1 NOR3_123( .ZN(n225gat), .A1(n231gat), .A2(n229gat), .A3(n228gat) );
  NOR3_X1 NOR3_124( .ZN(n121gat), .A1(n125gat), .A2(n126gat), .A3(n127gat) );
  NOR3_X1 NOR3_125( .ZN(n122gat), .A1(n125gat), .A2(n128gat), .A3(n129gat) );
  NOR3_X1 NOR3_126( .ZN(n123gat), .A1(n130gat), .A2(n126gat), .A3(n129gat) );
  NOR3_X1 NOR3_127( .ZN(n124gat), .A1(n130gat), .A2(n128gat), .A3(n127gat) );
  NOR2_X1 NOR2_111( .ZN(n2460gat), .A1(n666gat), .A2(n120gat) );
  NOR2_X1 NOR2_112( .ZN(n2423gat), .A1(n665gat), .A2(n1601gat) );
  NOR3_X1 NOR3_128( .ZN(n2594gat), .A1(n3017gat), .A2(n2520gat), .A3(n2597gat) );
  NOR3_X1 NOR3_129( .ZN(n2569gat), .A1(n2573gat), .A2(n2574gat), .A3(n2575gat) );
  NOR3_X1 NOR3_130( .ZN(n2570gat), .A1(n2573gat), .A2(n2576gat), .A3(n2577gat) );
  NOR3_X1 NOR3_131( .ZN(n2571gat), .A1(n2578gat), .A2(n2574gat), .A3(n2577gat) );
  NOR3_X1 NOR3_132( .ZN(n2572gat), .A1(n2578gat), .A2(n2576gat), .A3(n2575gat) );
  NOR3_X1 NOR3_133( .ZN(n2410gat), .A1(n2414gat), .A2(n2415gat), .A3(n2416gat) );
  NOR3_X1 NOR3_134( .ZN(n2411gat), .A1(n2414gat), .A2(n2417gat), .A3(n2418gat) );
  NOR3_X1 NOR3_135( .ZN(n2412gat), .A1(n2419gat), .A2(n2415gat), .A3(n2418gat) );
  NOR3_X1 NOR3_136( .ZN(n2413gat), .A1(n2419gat), .A2(n2417gat), .A3(n2416gat) );
  NOR2_X1 NOR2_113( .ZN(n2583gat), .A1(n2582gat), .A2(n2585gat) );
  NOR2_X1 NOR2_114( .ZN(n2580gat), .A1(n2582gat), .A2(n2583gat) );
  NOR2_X2 NOR2_115( .ZN(n2581gat), .A1(n2583gat), .A2(n2585gat) );
  NOR2_X1 NOR2_116( .ZN(n2567gat), .A1(n2493gat), .A2(n2388gat) );
  NOR2_X1 NOR2_117( .ZN(n2499gat), .A1(n2389gat), .A2(n2494gat) );
  NOR2_X1 NOR2_118( .ZN(n299gat), .A1(n2268gat), .A2(n2338gat) );
  NOR2_X1 NOR2_119( .ZN(n207gat), .A1(n2337gat), .A2(n2269gat) );
  NOR2_X1 NOR2_120( .ZN(n2650gat), .A1(n2649gat), .A2(n2652gat) );
  NOR2_X1 NOR2_121( .ZN(n2647gat), .A1(n2649gat), .A2(n2650gat) );
  NOR2_X1 NOR2_122( .ZN(n2648gat), .A1(n2650gat), .A2(n2652gat) );
  NOR3_X1 NOR3_137( .ZN(n2602gat), .A1(n2606gat), .A2(n2607gat), .A3(n2608gat) );
  NOR3_X1 NOR3_138( .ZN(n2603gat), .A1(n2606gat), .A2(n2609gat), .A3(n2610gat) );
  NOR3_X1 NOR3_139( .ZN(n2604gat), .A1(n2611gat), .A2(n2607gat), .A3(n2610gat) );
  NOR3_X1 NOR3_140( .ZN(n2605gat), .A1(n2611gat), .A2(n2609gat), .A3(n2608gat) );
  NOR3_X1 NOR3_141( .ZN(n2546gat), .A1(n2550gat), .A2(n2551gat), .A3(n2552gat) );
  NOR3_X1 NOR3_142( .ZN(n2547gat), .A1(n2550gat), .A2(n2553gat), .A3(n2554gat) );
  NOR3_X1 NOR3_143( .ZN(n2548gat), .A1(n2555gat), .A2(n2551gat), .A3(n2554gat) );
  NOR3_X1 NOR3_144( .ZN(n2549gat), .A1(n2555gat), .A2(n2553gat), .A3(n2552gat) );
  NOR2_X1 NOR2_123( .ZN(n2617gat), .A1(n2616gat), .A2(n2619gat) );
  NOR2_X1 NOR2_124( .ZN(n2614gat), .A1(n2616gat), .A2(n2617gat) );
  NOR2_X1 NOR2_125( .ZN(n2615gat), .A1(n2617gat), .A2(n2619gat) );
  NOR3_X2 NOR4_3_A( .ZN(extra3), .A1(n2508gat), .A2(n2656gat), .A3(n2500gat) );
  NOR2_X1 NOR4_3( .ZN(n2655gat), .A1(extra3), .A2(n2504gat) );
  NOR3_X1 NOR3_145( .ZN(n2293gat), .A1(n2353gat), .A2(n2284gat), .A3(n2443gat) );
  NOR2_X1 NOR2_126( .ZN(n2219gat), .A1(n2354gat), .A2(n2214gat) );
  NOR2_X1 NOR2_127( .ZN(n1529gat), .A1(n1528gat), .A2(n1523gat) );
  NOR2_X1 NOR2_128( .ZN(n1704gat), .A1(n3027gat), .A2(n1706gat) );
  NOR2_X1 NOR2_129( .ZN(n2461gat), .A1(n120gat), .A2(n2666gat) );
  NOR2_X1 NOR2_130( .ZN(n2421gat), .A1(n1601gat), .A2(n1704gat) );
  NOR2_X1 NOR2_131( .ZN(n1598gat), .A1(n1592gat), .A2(n2422gat) );
  NOR2_X1 NOR2_132( .ZN(n2218gat), .A1(n2214gat), .A2(n2290gat) );
  NOR3_X1 NOR3_146( .ZN(n2358gat), .A1(n2285gat), .A2(n2356gat), .A3(n2355gat) );
  NOR2_X1 NOR2_133( .ZN(n1415gat), .A1(n2081gat), .A2(n2359gat) );
  NOR2_X1 NOR2_134( .ZN(n1153gat), .A1(n1414gat), .A2(n566gat) );
  NOR3_X1 NOR3_147( .ZN(n2292gat), .A1(n2443gat), .A2(n2284gat), .A3(n2285gat) );
  NOR2_X1 NOR2_135( .ZN(n1416gat), .A1(n2081gat), .A2(n1480gat) );
  NOR2_X1 NOR2_136( .ZN(n1151gat), .A1(n1301gat), .A2(n1150gat) );
  NOR3_X1 NOR3_148( .ZN(n2306gat), .A1(n2356gat), .A2(n2284gat), .A3(n2285gat) );
  NOR2_X1 NOR2_137( .ZN(n1481gat), .A1(n2081gat), .A2(n2011gat) );
  NOR2_X1 NOR2_138( .ZN(n982gat), .A1(n873gat), .A2(n1478gat) );
  NOR3_X2 NOR3_149( .ZN(n2357gat), .A1(n2285gat), .A2(n2355gat), .A3(n2443gat) );
  NOR2_X1 NOR2_139( .ZN(n1347gat), .A1(n2081gat), .A2(n1410gat) );
  NOR2_X1 NOR2_140( .ZN(n877gat), .A1(n875gat), .A2(n876gat) );
  NOR2_X1 NOR2_141( .ZN(n1484gat), .A1(n2081gat), .A2(n1528gat) );
  NOR2_X1 NOR2_142( .ZN(n1159gat), .A1(n1160gat), .A2(n1084gat) );
  NOR3_X1 NOR3_150( .ZN(n2363gat), .A1(n2353gat), .A2(n2356gat), .A3(n2355gat) );
  NOR2_X1 NOR2_143( .ZN(n1483gat), .A1(n2081gat), .A2(n1482gat) );
  NOR2_X1 NOR2_144( .ZN(n1158gat), .A1(n983gat), .A2(n1157gat) );
  NOR3_X1 NOR3_151( .ZN(n2364gat), .A1(n2353gat), .A2(n2284gat), .A3(n2356gat) );
  NOR2_X1 NOR2_145( .ZN(n1308gat), .A1(n2081gat), .A2(n1530gat) );
  NOR2_X1 NOR2_146( .ZN(n1156gat), .A1(n985gat), .A2(n1307gat) );
  NOR3_X1 NOR3_152( .ZN(n2291gat), .A1(n2353gat), .A2(n2355gat), .A3(n2443gat) );
  NOR2_X1 NOR2_147( .ZN(n1349gat), .A1(n1479gat), .A2(n2081gat) );
  NOR2_X1 NOR2_148( .ZN(n1155gat), .A1(n1085gat), .A2(n1348gat) );
  NOR3_X1 NOR3_153( .ZN(n1154gat), .A1(n1598gat), .A2(n2930gat), .A3(n2957gat) );
  NOR2_X1 NOR2_149( .ZN(n1703gat), .A1(n1705gat), .A2(n3028gat) );
  NOR2_X1 NOR2_150( .ZN(n1608gat), .A1(n1704gat), .A2(n1703gat) );
  NOR2_X1 NOR2_151( .ZN(n1411gat), .A1(n1154gat), .A2(n1608gat) );
  NOR2_X2 NOR2_152( .ZN(n2223gat), .A1(n2354gat), .A2(n2217gat) );
  NOR2_X1 NOR2_153( .ZN(n1438gat), .A1(n1591gat), .A2(n1480gat) );
  NOR2_X1 NOR2_154( .ZN(n1625gat), .A1(n3021gat), .A2(n1628gat) );
  NOR2_X1 NOR2_155( .ZN(n1626gat), .A1(n1627gat), .A2(n3022gat) );
  NOR3_X1 NOR3_154( .ZN(n1831gat), .A1(n1832gat), .A2(n1765gat), .A3(n1878gat) );
  NOR2_X1 NOR2_156( .ZN(n1443gat), .A1(n1442gat), .A2(n706gat) );
  NOR2_X1 NOR2_157( .ZN(n1325gat), .A1(n1444gat), .A2(n164gat) );
  NOR2_X1 NOR2_158( .ZN(n1441gat), .A1(n1437gat), .A2(n1378gat) );
  NOR2_X1 NOR2_159( .ZN(n1321gat), .A1(n1442gat), .A2(n837gat) );
  NOR2_X1 NOR2_160( .ZN(n1320gat), .A1(n1444gat), .A2(n278gat) );
  NOR2_X1 NOR2_161( .ZN(n1486gat), .A1(n1482gat), .A2(n1591gat) );
  NOR2_X1 NOR2_162( .ZN(n1440gat), .A1(n1322gat), .A2(n1439gat) );
  NOR2_X1 NOR2_163( .ZN(n1426gat), .A1(n2011gat), .A2(n1591gat) );
  NOR2_X1 NOR2_164( .ZN(n1368gat), .A1(n1442gat), .A2(n613gat) );
  NOR2_X1 NOR2_165( .ZN(n1258gat), .A1(n274gat), .A2(n1444gat) );
  NOR2_X1 NOR2_166( .ZN(n1371gat), .A1(n1370gat), .A2(n1369gat) );
  NOR2_X1 NOR2_167( .ZN(n1365gat), .A1(n1479gat), .A2(n1591gat) );
  NOR2_X1 NOR2_168( .ZN(n1373gat), .A1(n833gat), .A2(n1442gat) );
  NOR2_X1 NOR2_169( .ZN(n1372gat), .A1(n282gat), .A2(n1444gat) );
  NOR2_X1 NOR2_170( .ZN(n1367gat), .A1(n1366gat), .A2(n1374gat) );
  NOR2_X2 NOR2_171( .ZN(n2220gat), .A1(n2290gat), .A2(n2217gat) );
  NOR2_X1 NOR2_172( .ZN(n1423gat), .A1(n2162gat), .A2(n1530gat) );
  NOR2_X1 NOR2_173( .ZN(n1498gat), .A1(n1609gat), .A2(n1427gat) );
  NOR2_X1 NOR2_174( .ZN(n1504gat), .A1(n1450gat), .A2(n1498gat) );
  NOR2_X1 NOR2_175( .ZN(n1607gat), .A1(n2082gat), .A2(n1609gat) );
  NOR2_X1 NOR2_176( .ZN(n1494gat), .A1(n1528gat), .A2(n2162gat) );
  NOR2_X1 NOR2_177( .ZN(n1502gat), .A1(n1607gat), .A2(n1449gat) );
  NOR2_X1 NOR2_178( .ZN(n1250gat), .A1(n1603gat), .A2(n815gat) );
  NOR2_X1 NOR2_179( .ZN(n1103gat), .A1(n956gat), .A2(n1590gat) );
  NOR2_X1 NOR2_180( .ZN(n1417gat), .A1(n2162gat), .A2(n1480gat) );
  NOR2_X1 NOR2_181( .ZN(n1352gat), .A1(n1248gat), .A2(n1418gat) );
  NOR2_X1 NOR2_182( .ZN(n1304gat), .A1(n1590gat), .A2(n1067gat) );
  NOR2_X1 NOR2_183( .ZN(n1249gat), .A1(n679gat), .A2(n1603gat) );
  NOR2_X1 NOR2_184( .ZN(n1419gat), .A1(n2162gat), .A2(n1479gat) );
  NOR2_X1 NOR2_185( .ZN(n1351gat), .A1(n1306gat), .A2(n1353gat) );
  NOR2_X1 NOR2_186( .ZN(n1246gat), .A1(n864gat), .A2(n1590gat) );
  NOR2_X1 NOR2_187( .ZN(n1161gat), .A1(n583gat), .A2(n1603gat) );
  NOR2_X1 NOR2_188( .ZN(n1422gat), .A1(n2011gat), .A2(n2162gat) );
  NOR2_X1 NOR2_189( .ZN(n1303gat), .A1(n1247gat), .A2(n1355gat) );
  NOR2_X1 NOR2_190( .ZN(n1291gat), .A1(n1603gat), .A2(n579gat) );
  NOR2_X1 NOR2_191( .ZN(n1245gat), .A1(n1590gat), .A2(n860gat) );
  NOR2_X1 NOR2_192( .ZN(n1485gat), .A1(n1482gat), .A2(n2162gat) );
  NOR2_X2 NOR2_193( .ZN(n1302gat), .A1(n1300gat), .A2(n1487gat) );
  NOR2_X1 NOR2_194( .ZN(n1163gat), .A1(n882gat), .A2(n1603gat) );
  NOR2_X1 NOR2_195( .ZN(n1102gat), .A1(n1297gat), .A2(n1590gat) );
  NOR2_X1 NOR2_196( .ZN(n1354gat), .A1(n1591gat), .A2(n1530gat) );
  NOR2_X1 NOR2_197( .ZN(n1360gat), .A1(n1164gat), .A2(n1356gat) );
  NOR2_X1 NOR2_198( .ZN(n1435gat), .A1(n1591gat), .A2(n1528gat) );
  NOR2_X1 NOR2_199( .ZN(n1101gat), .A1(n1590gat), .A2(n1293gat) );
  NOR2_X1 NOR2_200( .ZN(n996gat), .A1(n1603gat), .A2(n823gat) );
  NOR2_X1 NOR2_201( .ZN(n1359gat), .A1(n1436gat), .A2(n1106gat) );
  NOR2_X1 NOR2_202( .ZN(n1421gat), .A1(n2162gat), .A2(n2359gat) );
  NOR2_X1 NOR2_203( .ZN(n1104gat), .A1(n1079gat), .A2(n1590gat) );
  NOR2_X1 NOR2_204( .ZN(n887gat), .A1(n1603gat), .A2(n683gat) );
  NOR2_X1 NOR2_205( .ZN(n1358gat), .A1(n1425gat), .A2(n1105gat) );
  NOR2_X1 NOR2_206( .ZN(n1420gat), .A1(n1410gat), .A2(n2162gat) );
  NOR2_X2 NOR2_207( .ZN(n1305gat), .A1(n1147gat), .A2(n1590gat) );
  NOR2_X2 NOR2_208( .ZN(n1162gat), .A1(n698gat), .A2(n1603gat) );
  NOR2_X2 NOR2_209( .ZN(n1357gat), .A1(n1424gat), .A2(n1309gat) );
  NOR3_X1 NOR4_4_A( .ZN(extra4), .A1(n2978gat), .A2(n2982gat), .A3(n2973gat) );
  NOR2_X1 NOR4_4( .ZN(n1428gat), .A1(extra4), .A2(n2977gat) );
  NOR2_X1 NOR2_210( .ZN(n1794gat), .A1(n1673gat), .A2(n1719gat) );
  NOR2_X1 NOR2_211( .ZN(n1796gat), .A1(n1858gat), .A2(n1635gat) );
  NOR2_X1 NOR2_212( .ZN(n1792gat), .A1(n1794gat), .A2(n1796gat) );
  NOR3_X1 NOR3_155( .ZN(n1865gat), .A1(n1989gat), .A2(n1918gat), .A3(n1986gat) );
  NOR3_X1 NOR3_156( .ZN(n1861gat), .A1(n1866gat), .A2(n2216gat), .A3(n1988gat) );
  NOR2_X1 NOR2_213( .ZN(n1793gat), .A1(n1792gat), .A2(n1735gat) );
  NOR2_X1 NOR2_214( .ZN(n1406gat), .A1(n1428gat), .A2(n1387gat) );
  NOR3_X1 NOR3_157( .ZN(n1780gat), .A1(n1777gat), .A2(n1625gat), .A3(n1626gat) );
  NOR2_X1 NOR2_215( .ZN(n2016gat), .A1(n2019gat), .A2(n1878gat) );
  NOR2_X1 NOR2_216( .ZN(n2664gat), .A1(n2850gat), .A2(n3018gat) );
  NOR3_X1 NOR3_158( .ZN(n1666gat), .A1(n1986gat), .A2(n2212gat), .A3(n1991gat) );
  NOR3_X1 NOR3_159( .ZN(n1578gat), .A1(n2152gat), .A2(n2351gat), .A3(n1665gat) );
  NOR2_X1 NOR2_217( .ZN(n1516gat), .A1(n1551gat), .A2(n1517gat) );
  NOR3_X1 NOR3_160( .ZN(n1864gat), .A1(n1858gat), .A2(n1495gat), .A3(n2090gat) );
  NOR2_X1 NOR2_218( .ZN(n1565gat), .A1(n1735gat), .A2(n1552gat) );
  NOR2_X1 NOR2_219( .ZN(n1921gat), .A1(n1738gat), .A2(n1673gat) );
  NOR2_X1 NOR2_220( .ZN(n1798gat), .A1(n1739gat), .A2(n1673gat) );
  NOR3_X1 NOR3_161( .ZN(n1920gat), .A1(n1864gat), .A2(n1921gat), .A3(n1798gat) );
  NOR2_X1 NOR2_221( .ZN(n1926gat), .A1(n1925gat), .A2(n1635gat) );
  NOR2_X1 NOR2_222( .ZN(n1916gat), .A1(n1917gat), .A2(n1859gat) );
  NOR2_X1 NOR2_223( .ZN(n1994gat), .A1(n1719gat), .A2(n1922gat) );
  NOR2_X1 NOR2_224( .ZN(n1924gat), .A1(n1743gat), .A2(n1923gat) );
  NOR3_X1 NOR4_5_A( .ZN(extra5), .A1(n1926gat), .A2(n1916gat), .A3(n1994gat) );
  NOR2_X1 NOR4_5( .ZN(n2078gat), .A1(extra5), .A2(n1924gat) );
  NOR2_X1 NOR2_225( .ZN(n1690gat), .A1(n1700gat), .A2(n1702gat) );
  NOR3_X1 NOR3_162( .ZN(n1660gat), .A1(n1918gat), .A2(n1986gat), .A3(n2212gat) );
  NOR3_X1 NOR3_163( .ZN(n1576gat), .A1(n2351gat), .A2(n1988gat), .A3(n1661gat) );
  NOR2_X1 NOR2_226( .ZN(n1733gat), .A1(n1673gat), .A2(n1572gat) );
  NOR3_X1 NOR3_164( .ZN(n1582gat), .A1(n2283gat), .A2(n1991gat), .A3(n2212gat) );
  NOR3_X1 NOR3_165( .ZN(n1577gat), .A1(n1520gat), .A2(n2351gat), .A3(n1988gat) );
  NOR2_X1 NOR2_227( .ZN(n1581gat), .A1(n1858gat), .A2(n1580gat) );
  NOR3_X1 NOR3_166( .ZN(n2129gat), .A1(n2189gat), .A2(n2134gat), .A3(n2261gat) );
  NOR3_X1 NOR4_6_A( .ZN(extra6), .A1(n2078gat), .A2(n2178gat), .A3(n1990gat) );
  NOR2_X1 NOR4_6( .ZN(n2079gat), .A1(extra6), .A2(n2128gat) );
  NOR3_X1 NOR4_7_A( .ZN(extra7), .A1(n1609gat), .A2(n1778gat), .A3(n1704gat) );
  NOR2_X1 NOR4_7( .ZN(n1695gat), .A1(extra7), .A2(n1703gat) );
  NOR3_X1 NOR3_167( .ZN(n2073gat), .A1(n2078gat), .A2(n1990gat), .A3(n2181gat) );
  NOR2_X1 NOR2_228( .ZN(n1696gat), .A1(n1707gat), .A2(n1698gat) );
  NOR2_X1 NOR2_229( .ZN(n1758gat), .A1(n1311gat), .A2(n1773gat) );
  NOR3_X1 NOR3_168( .ZN(n1574gat), .A1(n1719gat), .A2(n1673gat), .A3(n1444gat) );
  NOR3_X1 NOR3_169( .ZN(n1573gat), .A1(n1444gat), .A2(n1858gat), .A3(n1635gat) );
  NOR2_X1 NOR2_230( .ZN(n1521gat), .A1(n2283gat), .A2(n1991gat) );
  NOR2_X1 NOR2_231( .ZN(n1737gat), .A1(n2212gat), .A2(n2152gat) );
  NOR3_X1 NOR3_170( .ZN(n1732gat), .A1(n1515gat), .A2(n1736gat), .A3(n1658gat) );
  NOR3_X1 NOR3_171( .ZN(n1723gat), .A1(n1659gat), .A2(n1722gat), .A3(n1724gat) );
  NOR2_X1 NOR2_232( .ZN(n1663gat), .A1(n1986gat), .A2(n1918gat) );
  NOR3_X1 NOR3_172( .ZN(n1655gat), .A1(n1736gat), .A2(n1662gat), .A3(n1658gat) );
  NOR3_X1 NOR3_173( .ZN(n1647gat), .A1(n1656gat), .A2(n1659gat), .A3(n1554gat) );
  NOR2_X1 NOR2_233( .ZN(n1667gat), .A1(n1991gat), .A2(n1986gat) );
  NOR3_X1 NOR3_174( .ZN(n1570gat), .A1(n1736gat), .A2(n1658gat), .A3(n1670gat) );
  NOR3_X1 NOR3_175( .ZN(n1646gat), .A1(n1569gat), .A2(n1659gat), .A3(n1566gat) );
  NOR2_X1 NOR2_234( .ZN(n1575gat), .A1(n1918gat), .A2(n2283gat) );
  NOR3_X1 NOR3_176( .ZN(n1728gat), .A1(n1568gat), .A2(n1736gat), .A3(n1658gat) );
  NOR3_X1 NOR3_177( .ZN(n1650gat), .A1(n1727gat), .A2(n1659gat), .A3(n1640gat) );
  NOR2_X1 NOR2_235( .ZN(n1801gat), .A1(n2152gat), .A2(n1989gat) );
  NOR3_X1 NOR3_178( .ZN(n1731gat), .A1(n1658gat), .A2(n1515gat), .A3(n1797gat) );
  NOR3_X1 NOR3_179( .ZN(n1649gat), .A1(n1560gat), .A2(n1659gat), .A3(n1730gat) );
  NOR3_X1 NOR3_180( .ZN(n1571gat), .A1(n1670gat), .A2(n1658gat), .A3(n1797gat) );
  NOR3_X1 NOR3_181( .ZN(n1563gat), .A1(n1561gat), .A2(n1562gat), .A3(n1659gat) );
  NOR2_X1 NOR2_236( .ZN(n1734gat), .A1(n1988gat), .A2(n2212gat) );
  NOR3_X1 NOR3_182( .ZN(n1669gat), .A1(n1668gat), .A2(n1742gat), .A3(n1670gat) );
  NOR2_X1 NOR2_237( .ZN(n1654gat), .A1(n1671gat), .A2(n1659gat) );
  NOR3_X1 NOR3_183( .ZN(n1657gat), .A1(n1662gat), .A2(n1797gat), .A3(n1658gat) );
  NOR3_X2 NOR3_184( .ZN(n1653gat), .A1(n1651gat), .A2(n1652gat), .A3(n1659gat) );
  NOR3_X2 NOR3_185( .ZN(n1729gat), .A1(n1658gat), .A2(n1797gat), .A3(n1568gat) );
  NOR3_X1 NOR3_186( .ZN(n1644gat), .A1(n1643gat), .A2(n1648gat), .A3(n1659gat) );
  NOR3_X1 NOR3_187( .ZN(n1726gat), .A1(n2992gat), .A2(n2986gat), .A3(n2991gat) );
  NOR2_X1 NOR2_238( .ZN(n1929gat), .A1(n1758gat), .A2(n1790gat) );
  NOR3_X1 NOR3_188( .ZN(n2009gat), .A1(n2016gat), .A2(n2664gat), .A3(n2004gat) );
  NOR3_X1 NOR3_189( .ZN(n1413gat), .A1(n1869gat), .A2(n672gat), .A3(n2591gat) );
  NOR2_X1 NOR2_239( .ZN(n1636gat), .A1(n1584gat), .A2(n1718gat) );
  NOR2_X1 NOR2_240( .ZN(n1401gat), .A1(n1584gat), .A2(n1590gat) );
  NOR3_X1 NOR3_190( .ZN(n1408gat), .A1(n1507gat), .A2(n1396gat), .A3(n1393gat) );
  NOR2_X1 NOR2_241( .ZN(n1476gat), .A1(n1858gat), .A2(n1590gat) );
  NOR3_X1 NOR3_191( .ZN(n1407gat), .A1(n1393gat), .A2(n1409gat), .A3(n1677gat) );
  NOR3_X1 NOR3_192( .ZN(n1412gat), .A1(n1411gat), .A2(n1406gat), .A3(n2981gat) );
  NOR3_X1 NOR3_193( .ZN(n2663gat), .A1(n2586gat), .A2(n2660gat), .A3(n2307gat) );
  NOR2_X1 NOR2_242( .ZN(n2662gat), .A1(n2660gat), .A2(n2586gat) );
  NOR2_X1 NOR2_243( .ZN(n2238gat), .A1(n2448gat), .A2(n2444gat) );
  NOR3_X1 NOR3_194( .ZN(n87gat), .A1(n743gat), .A2(n17gat), .A3(n293gat) );
  NOR2_X1 NOR2_244( .ZN(n200gat), .A1(n199gat), .A2(n92gat) );
  NOR3_X1 NOR3_195( .ZN(n184gat), .A1(n189gat), .A2(n188gat), .A3(n179gat) );
  NOR2_X1 NOR2_245( .ZN(n196gat), .A1(n297gat), .A2(n195gat) );
  NOR2_X1 NOR2_246( .ZN(n204gat), .A1(n200gat), .A2(n196gat) );
  NOR3_X1 NOR4_8_A( .ZN(extra8), .A1(n1790gat), .A2(n1310gat), .A3(n2664gat) );
  NOR2_X1 NOR4_8( .ZN(n2163gat), .A1(extra8), .A2(n2168gat) );
  NOR2_X1 NOR2_247( .ZN(n2258gat), .A1(n2260gat), .A2(n2189gat) );
  NOR2_X1 NOR2_248( .ZN(n2255gat), .A1(n2261gat), .A2(n2188gat) );
  NOR3_X1 NOR3_196( .ZN(n2015gat), .A1(n2039gat), .A2(n1774gat), .A3(n1315gat) );
  NOR2_X2 NOR2_249( .ZN(n2017gat), .A1(n1790gat), .A2(n2016gat) );
  NOR2_X1 NOR2_250( .ZN(n2018gat), .A1(n2016gat), .A2(n2097gat) );
  NOR3_X1 NOR4_9_A( .ZN(extra9), .A1(n2035gat), .A2(n2093gat), .A3(n2018gat) );
  NOR2_X1 NOR4_9( .ZN(n2014gat), .A1(extra9), .A2(n2664gat) );
  NOR2_X1 NOR2_251( .ZN(n2194gat), .A1(n2187gat), .A2(n1855gat) );
  NOR2_X1 NOR2_252( .ZN(n2192gat), .A1(n2184gat), .A2(n1855gat) );
  NOR2_X1 NOR2_253( .ZN(n2185gat), .A1(n2261gat), .A2(n2189gat) );
  NOR2_X1 NOR2_254( .ZN(n2132gat), .A1(n2133gat), .A2(n2131gat) );
  NOR2_X1 NOR2_255( .ZN(n2130gat), .A1(n2134gat), .A2(n2185gat) );
  NOR2_X1 NOR2_256( .ZN(n2057gat), .A1(n2049gat), .A2(n1855gat) );
  NOR2_X1 NOR2_257( .ZN(n2250gat), .A1(n2248gat), .A2(n2264gat) );
  NOR2_X1 NOR2_258( .ZN(n2249gat), .A1(n2265gat), .A2(n3006gat) );
  NOR2_X1 NOR2_259( .ZN(n2329gat), .A1(n1855gat), .A2(n3007gat) );
  NOR2_X1 NOR2_260( .ZN(n1958gat), .A1(n1963gat), .A2(n1886gat) );
  NOR3_X1 NOR3_197( .ZN(n1895gat), .A1(n1845gat), .A2(n1891gat), .A3(n1968gat) );
  NOR2_X1 NOR2_261( .ZN(n1710gat), .A1(n1709gat), .A2(n1629gat) );
  NOR2_X1 NOR2_262( .ZN(n1630gat), .A1(n1895gat), .A2(n1631gat) );
  NOR2_X1 NOR2_263( .ZN(n2195gat), .A1(n2200gat), .A2(n1855gat) );
  NOR2_X1 NOR2_264( .ZN(n2556gat), .A1(n1711gat), .A2(n2437gat) );
  NOR2_X1 NOR2_265( .ZN(n2539gat), .A1(n2048gat), .A2(n2437gat) );
  NOR3_X1 NOR3_198( .ZN(n1894gat), .A1(n1968gat), .A2(n1891gat), .A3(n1969gat) );
  NOR2_X2 NOR2_266( .ZN(n1847gat), .A1(n1958gat), .A2(n1845gat) );
  NOR2_X2 NOR2_267( .ZN(n1846gat), .A1(n1845gat), .A2(n1893gat) );
  NOR2_X1 NOR2_268( .ZN(n2436gat), .A1(n2437gat), .A2(n1892gat) );
  NOR2_X1 NOR2_269( .ZN(n2055gat), .A1(n1891gat), .A2(n1958gat) );
  NOR2_X1 NOR2_270( .ZN(n1967gat), .A1(n1893gat), .A2(n1968gat) );
  NOR2_X1 NOR2_271( .ZN(n2387gat), .A1(n2056gat), .A2(n2437gat) );
  NOR2_X1 NOR2_272( .ZN(n1959gat), .A1(n1956gat), .A2(n1963gat) );
  NOR2_X1 NOR2_273( .ZN(n1957gat), .A1(n1886gat), .A2(n1887gat) );
  NOR2_X1 NOR2_274( .ZN(n2330gat), .A1(n2437gat), .A2(n1961gat) );
  NOR2_X1 NOR2_275( .ZN(n2147gat), .A1(n2988gat), .A2(n1855gat) );
  NOR2_X1 NOR2_276( .ZN(n2498gat), .A1(n2199gat), .A2(n2328gat) );
  NOR2_X1 NOR2_277( .ZN(n2193gat), .A1(n2393gat), .A2(n2439gat) );
  NOR2_X1 NOR2_278( .ZN(n2211gat), .A1(n2193gat), .A2(n2402gat) );
  NOR2_X1 NOR2_279( .ZN(n2210gat), .A1(n2401gat), .A2(n2151gat) );
  NOR2_X1 NOR2_280( .ZN(n2396gat), .A1(n2199gat), .A2(n2209gat) );
  NOR2_X1 NOR2_281( .ZN(n2053gat), .A1(n2393gat), .A2(n2438gat) );
  NOR2_X1 NOR2_282( .ZN(n1964gat), .A1(n2392gat), .A2(n2439gat) );
  NOR2_X1 NOR2_283( .ZN(n2198gat), .A1(n2199gat), .A2(n2058gat) );
  NOR3_X1 NOR3_199( .ZN(n2215gat), .A1(n2346gat), .A2(n2151gat), .A3(n2402gat) );
  NOR2_X1 NOR2_284( .ZN(n2350gat), .A1(n2405gat), .A2(n2349gat) );
  NOR2_X1 NOR2_285( .ZN(n2282gat), .A1(n2406gat), .A2(n2215gat) );
  NOR2_X1 NOR2_286( .ZN(n2197gat), .A1(n2199gat), .A2(n2281gat) );
  NOR3_X1 NOR3_200( .ZN(n2213gat), .A1(n2402gat), .A2(n2151gat), .A3(n2345gat) );
  NOR2_X1 NOR2_287( .ZN(n2150gat), .A1(n2401gat), .A2(n2346gat) );
  NOR2_X1 NOR2_288( .ZN(n2149gat), .A1(n2193gat), .A2(n2346gat) );
  NOR2_X1 NOR2_289( .ZN(n2196gat), .A1(n2199gat), .A2(n2146gat) );
  NOR3_X1 NOR3_201( .ZN(n1882gat), .A1(n2124gat), .A2(n2115gat), .A3(n2239gat) );
  NOR2_X1 NOR2_290( .ZN(n1962gat), .A1(n1963gat), .A2(n1893gat) );
  NOR2_X1 NOR2_291( .ZN(n1896gat), .A1(n2995gat), .A2(n1895gat) );
  NOR2_X1 NOR2_292( .ZN(n1972gat), .A1(n1974gat), .A2(n1970gat) );
  NOR2_X1 NOR2_293( .ZN(n1971gat), .A1(n1896gat), .A2(n1973gat) );
  NOR2_X1 NOR2_294( .ZN(n2559gat), .A1(n2999gat), .A2(n2437gat) );
  NOR2_X1 NOR2_295( .ZN(n2331gat), .A1(n2393gat), .A2(n2401gat) );
  NOR2_X2 NOR2_296( .ZN(n2352gat), .A1(n3011gat), .A2(n2215gat) );
  NOR2_X1 NOR2_297( .ZN(n2566gat), .A1(n2643gat), .A2(n2564gat) );
  NOR2_X1 NOR2_298( .ZN(n2565gat), .A1(n2352gat), .A2(n2642gat) );
  NOR2_X1 NOR2_299( .ZN(n2637gat), .A1(n3015gat), .A2(n2199gat) );
  NOR3_X1 NOR3_202( .ZN(n84gat), .A1(n296gat), .A2(n17gat), .A3(n294gat) );
  NOR2_X1 NOR2_300( .ZN(n89gat), .A1(n88gat), .A2(n2784gat) );
  NOR2_X1 NOR2_301( .ZN(n110gat), .A1(n182gat), .A2(n89gat) );
  NOR2_X1 NOR2_302( .ZN(n1074gat), .A1(n2775gat), .A2(n110gat) );
  NOR3_X1 NOR3_203( .ZN(n141gat), .A1(n155gat), .A2(n253gat), .A3(n150gat) );
  NOR2_X1 NOR2_303( .ZN(n38gat), .A1(n151gat), .A2(n233gat) );
  NOR2_X1 NOR2_304( .ZN(n37gat), .A1(n151gat), .A2(n154gat) );
  NOR2_X1 NOR2_305( .ZN(n872gat), .A1(n375gat), .A2(n800gat) );
  NOR2_X1 NOR2_306( .ZN(n234gat), .A1(n155gat), .A2(n233gat) );
  NOR2_X1 NOR2_307( .ZN(n137gat), .A1(n154gat), .A2(n253gat) );
  NOR2_X1 NOR2_308( .ZN(n378gat), .A1(n375gat), .A2(n235gat) );
  NOR2_X1 NOR2_309( .ZN(n377gat), .A1(n110gat), .A2(n2778gat) );
  NOR2_X1 NOR2_310( .ZN(n869gat), .A1(n219gat), .A2(n2792gat) );
  NOR2_X1 NOR2_311( .ZN(n212gat), .A1(n182gat), .A2(n78gat) );
  NOR3_X1 NOR3_204( .ZN(n250gat), .A1(n329gat), .A2(n387gat), .A3(n334gat) );
  NOR2_X1 NOR2_312( .ZN(n249gat), .A1(n386gat), .A2(n330gat) );
  NOR2_X1 NOR2_313( .ZN(n248gat), .A1(n330gat), .A2(n1490gat) );
  NOR2_X1 NOR2_314( .ZN(n453gat), .A1(n372gat), .A2(n452gat) );
  NOR2_X1 NOR2_315( .ZN(n448gat), .A1(n111gat), .A2(n2846gat) );
  NOR2_X1 NOR2_316( .ZN(n974gat), .A1(n2844gat), .A2(n111gat) );
  NOR2_X1 NOR2_317( .ZN(n251gat), .A1(n1490gat), .A2(n387gat) );
  NOR2_X1 NOR2_318( .ZN(n244gat), .A1(n334gat), .A2(n386gat) );
  NOR2_X1 NOR2_319( .ZN(n973gat), .A1(n372gat), .A2(n333gat) );
  NOR2_X1 NOR2_320( .ZN(n870gat), .A1(n2669gat), .A2(n219gat) );
  NOR2_X1 NOR2_321( .ZN(n975gat), .A1(n111gat), .A2(n2852gat) );
  NOR3_X1 NOR3_205( .ZN(n246gat), .A1(n330gat), .A2(n325gat), .A3(n334gat) );
  NOR2_X1 NOR2_322( .ZN(n245gat), .A1(n386gat), .A2(n334gat) );
  NOR2_X1 NOR2_323( .ZN(n460gat), .A1(n462gat), .A2(n2884gat) );
  NOR2_X1 NOR2_324( .ZN(n459gat), .A1(n457gat), .A2(n461gat) );
  NOR2_X1 NOR2_325( .ZN(n972gat), .A1(n372gat), .A2(n458gat) );
  NOR2_X1 NOR2_326( .ZN(n969gat), .A1(n219gat), .A2(n2672gat) );
  NOR2_X1 NOR2_327( .ZN(n971gat), .A1(n111gat), .A2(n2840gat) );
  NOR3_X1 NOR3_206( .ZN(n247gat), .A1(n334gat), .A2(n387gat), .A3(n330gat) );
  NOR2_X1 NOR2_328( .ZN(n145gat), .A1(n144gat), .A2(n325gat) );
  NOR2_X1 NOR2_329( .ZN(n143gat), .A1(n326gat), .A2(n247gat) );
  NOR2_X1 NOR2_330( .ZN(n970gat), .A1(n372gat), .A2(n878gat) );
  NOR2_X1 NOR2_331( .ZN(n968gat), .A1(n2789gat), .A2(n219gat) );
  NOR2_X1 NOR2_332( .ZN(n772gat), .A1(n111gat), .A2(n2842gat) );
  NOR3_X1 NOR3_207( .ZN(n142gat), .A1(n382gat), .A2(n326gat), .A3(n144gat) );
  NOR2_X1 NOR2_333( .ZN(n40gat), .A1(n325gat), .A2(n383gat) );
  NOR2_X1 NOR2_334( .ZN(n39gat), .A1(n383gat), .A2(n247gat) );
  NOR2_X1 NOR2_335( .ZN(n451gat), .A1(n134gat), .A2(n372gat) );
  NOR2_X1 NOR2_336( .ZN(n446gat), .A1(n219gat), .A2(n2781gat) );
  NOR3_X1 NOR3_208( .ZN(n139gat), .A1(n253gat), .A2(n151gat), .A3(n254gat) );
  NOR2_X1 NOR2_337( .ZN(n136gat), .A1(n253gat), .A2(n154gat) );
  NOR2_X1 NOR2_338( .ZN(n391gat), .A1(n252gat), .A2(n468gat) );
  NOR2_X1 NOR2_339( .ZN(n390gat), .A1(n469gat), .A2(n2877gat) );
  NOR2_X2 NOR2_340( .ZN(n1083gat), .A1(n381gat), .A2(n375gat) );
  NOR2_X1 NOR2_341( .ZN(n1077gat), .A1(n110gat), .A2(n2672gat) );
  NOR3_X1 NOR3_209( .ZN(n140gat), .A1(n151gat), .A2(n253gat), .A3(n155gat) );
  NOR2_X1 NOR2_342( .ZN(n242gat), .A1(n254gat), .A2(n241gat) );
  NOR2_X1 NOR2_343( .ZN(n240gat), .A1(n255gat), .A2(n140gat) );
  NOR2_X1 NOR2_344( .ZN(n871gat), .A1(n802gat), .A2(n375gat) );
  NOR2_X1 NOR2_345( .ZN(n797gat), .A1(n110gat), .A2(n2734gat) );
  NOR3_X1 NOR3_210( .ZN(n324gat), .A1(n255gat), .A2(n146gat), .A3(n241gat) );
  NOR2_X1 NOR2_346( .ZN(n238gat), .A1(n147gat), .A2(n254gat) );
  NOR2_X1 NOR2_347( .ZN(n237gat), .A1(n140gat), .A2(n147gat) );
  NOR2_X1 NOR2_348( .ZN(n1082gat), .A1(n375gat), .A2(n380gat) );
  NOR2_X1 NOR2_349( .ZN(n796gat), .A1(n2731gat), .A2(n110gat) );
  NOR3_X1 NOR3_211( .ZN(n85gat), .A1(n17gat), .A2(n294gat), .A3(n637gat) );
  NOR3_X1 NOR3_212( .ZN(n180gat), .A1(n286gat), .A2(n188gat), .A3(n287gat) );
  NOR2_X1 NOR2_350( .ZN(n68gat), .A1(n85gat), .A2(n180gat) );
  NOR3_X1 NOR3_213( .ZN(n186gat), .A1(n189gat), .A2(n287gat), .A3(n288gat) );
  NOR2_X1 NOR2_351( .ZN(n357gat), .A1(n2726gat), .A2(n2860gat) );
  NOR3_X1 NOR3_214( .ZN(n82gat), .A1(n16gat), .A2(n295gat), .A3(n637gat) );
  NOR2_X1 NOR2_352( .ZN(n12gat), .A1(n186gat), .A2(n82gat) );
  NOR2_X1 NOR2_353( .ZN(n1599gat), .A1(n1691gat), .A2(n336gat) );
  NOR2_X1 NOR2_354( .ZN(n1613gat), .A1(n1544gat), .A2(n1698gat) );
  NOR3_X1 NOR3_215( .ZN(n1756gat), .A1(n2512gat), .A2(n1769gat), .A3(n1773gat) );
  NOR2_X1 NOR2_355( .ZN(n1586gat), .A1(n1869gat), .A2(n1683gat) );
  NOR3_X1 NOR3_216( .ZN(n1755gat), .A1(n1769gat), .A2(n1773gat), .A3(n2512gat) );
  NOR3_X1 NOR3_217( .ZN(n2538gat), .A1(n2620gat), .A2(n2625gat), .A3(n2488gat) );
  NOR3_X1 NOR3_218( .ZN(n2483gat), .A1(n2537gat), .A2(n2482gat), .A3(n2486gat) );
  NOR2_X1 NOR2_356( .ZN(n1391gat), .A1(n1513gat), .A2(n2442gat) );
  NOR3_X1 NOR3_219( .ZN(n1471gat), .A1(n1334gat), .A2(n1858gat), .A3(n1604gat) );
  NOR2_X1 NOR2_357( .ZN(n1469gat), .A1(n1858gat), .A2(n1608gat) );
  NOR3_X1 NOR3_220( .ZN(n1472gat), .A1(n1476gat), .A2(n1471gat), .A3(n1469gat) );
  NOR2_X1 NOR2_358( .ZN(n1927gat), .A1(n1790gat), .A2(n1635gat) );
  NOR2_X1 NOR2_359( .ZN(n1470gat), .A1(n1472gat), .A2(n1747gat) );
  NOR3_X1 NOR3_221( .ZN(n1402gat), .A1(n1858gat), .A2(n1393gat), .A3(n1604gat) );
  NOR2_X1 NOR2_360( .ZN(n1400gat), .A1(n1674gat), .A2(n1403gat) );
  NOR2_X1 NOR2_361( .ZN(n1567gat), .A1(n1634gat), .A2(n1735gat) );
  NOR3_X1 NOR3_222( .ZN(n1399gat), .A1(n1806gat), .A2(n1338gat), .A3(n1584gat) );
  NOR3_X1 NOR4_10_A( .ZN(extra10), .A1(n1584gat), .A2(n1719gat), .A3(n1790gat) );
  NOR2_X1 NOR4_10( .ZN(n1564gat), .A1(extra10), .A2(n1576gat) );
  NOR2_X1 NOR2_362( .ZN(n1600gat), .A1(n1685gat), .A2(n1427gat) );
  NOR3_X1 NOR3_223( .ZN(n1519gat), .A1(n1584gat), .A2(n1339gat), .A3(n1600gat) );
  NOR2_X1 NOR2_363( .ZN(n1397gat), .A1(n1519gat), .A2(n1401gat) );
  NOR2_X1 NOR2_364( .ZN(n1398gat), .A1(n1455gat), .A2(n1397gat) );
  NOR2_X1 NOR2_365( .ZN(n2008gat), .A1(n2012gat), .A2(n1774gat) );
  NOR2_X1 NOR2_366( .ZN(n2005gat), .A1(n2002gat), .A2(n2857gat) );
  NOR2_X2 NOR2_367( .ZN(n1818gat), .A1(n1823gat), .A2(n2005gat) );
  NOR3_X2 NOR3_224( .ZN(n1759gat), .A1(n1818gat), .A2(n1935gat), .A3(n2765gat) );
  NOR3_X2 NOR3_225( .ZN(n1686gat), .A1(n1774gat), .A2(n1869gat), .A3(n1684gat) );
  NOR2_X1 NOR2_368( .ZN(n1533gat), .A1(n1524gat), .A2(n1403gat) );
  NOR3_X1 NOR3_226( .ZN(n1863gat), .A1(n1991gat), .A2(n2283gat), .A3(n1989gat) );
  NOR3_X1 NOR3_227( .ZN(n1860gat), .A1(n1988gat), .A2(n2216gat), .A3(n1862gat) );
  NOR2_X1 NOR2_369( .ZN(n1915gat), .A1(n1859gat), .A2(n1919gat) );
  NOR2_X1 NOR2_370( .ZN(n1510gat), .A1(n1584gat), .A2(n1460gat) );
  NOR2_X1 NOR2_371( .ZN(n1800gat), .A1(n1635gat), .A2(n1919gat) );
  NOR2_X1 NOR2_372( .ZN(n1459gat), .A1(n1595gat), .A2(n1454gat) );
  NOR2_X1 NOR2_373( .ZN(n1458gat), .A1(n1510gat), .A2(n1459gat) );
  NOR2_X1 NOR2_374( .ZN(n1532gat), .A1(n1677gat), .A2(n1458gat) );
  NOR2_X1 NOR2_375( .ZN(n1467gat), .A1(n2289gat), .A2(n1468gat) );
  NOR3_X1 NOR3_228( .ZN(n1466gat), .A1(n1392gat), .A2(n1461gat), .A3(n1396gat) );
  NOR2_X1 NOR2_376( .ZN(n1531gat), .A1(n1507gat), .A2(n1477gat) );
  NOR2_X1 NOR2_377( .ZN(n1593gat), .A1(n1551gat), .A2(n1310gat) );
  NOR3_X1 NOR3_229( .ZN(n1602gat), .A1(n1594gat), .A2(n1587gat), .A3(n2989gat) );
  NOR3_X1 NOR3_230( .ZN(n1761gat), .A1(n2985gat), .A2(n1602gat), .A3(n1681gat) );
  NOR3_X1 NOR3_231( .ZN(n1760gat), .A1(n1681gat), .A2(n1602gat), .A3(n2985gat) );
  NOR3_X1 NOR3_232( .ZN(n1721gat), .A1(n2442gat), .A2(n1690gat), .A3(n1978gat) );
  NOR2_X1 NOR2_378( .ZN(n520gat), .A1(n374gat), .A2(n2862gat) );
  NOR2_X1 NOR2_379( .ZN(n519gat), .A1(n2854gat), .A2(n374gat) );
  NOR2_X1 NOR2_380( .ZN(n518gat), .A1(n520gat), .A2(n519gat) );
  NOR2_X1 NOR2_381( .ZN(n418gat), .A1(n374gat), .A2(n2723gat) );
  NOR2_X1 NOR2_382( .ZN(n411gat), .A1(n374gat), .A2(n2726gat) );
  NOR2_X1 NOR2_383( .ZN(n522gat), .A1(n374gat), .A2(n2859gat) );
  NOR2_X1 NOR2_384( .ZN(n516gat), .A1(n374gat), .A2(n2715gat) );
  NOR3_X1 NOR4_11_A( .ZN(extra11), .A1(n417gat), .A2(n413gat), .A3(n412gat) );
  NOR2_X1 NOR4_11( .ZN(n410gat), .A1(extra11), .A2(n406gat) );
  NOR2_X1 NOR2_385( .ZN(n354gat), .A1(n411gat), .A2(n522gat) );
  NOR3_X1 NOR3_233( .ZN(n355gat), .A1(n517gat), .A2(n410gat), .A3(n354gat) );
  NOR2_X1 NOR2_386( .ZN(n408gat), .A1(n516gat), .A2(n407gat) );
  NOR2_X1 NOR2_387( .ZN(n526gat), .A1(n2859gat), .A2(n740gat) );
  NOR2_X1 NOR2_388( .ZN(n531gat), .A1(n740gat), .A2(n2854gat) );
  NOR2_X1 NOR2_389( .ZN(n530gat), .A1(n2862gat), .A2(n740gat) );
  NOR3_X1 NOR3_234( .ZN(n525gat), .A1(n526gat), .A2(n531gat), .A3(n530gat) );
  NOR2_X1 NOR2_390( .ZN(n356gat), .A1(n2726gat), .A2(n740gat) );
  NOR2_X1 NOR2_391( .ZN(n415gat), .A1(n2723gat), .A2(n740gat) );
  NOR2_X1 NOR2_392( .ZN(n521gat), .A1(n740gat), .A2(n2715gat) );
  NOR3_X1 NOR3_235( .ZN(n532gat), .A1(n527gat), .A2(n416gat), .A3(n528gat) );
  NOR2_X1 NOR2_393( .ZN(n359gat), .A1(n290gat), .A2(n358gat) );
  NOR2_X1 NOR2_394( .ZN(n420gat), .A1(n408gat), .A2(n359gat) );
  NOR2_X1 NOR2_395( .ZN(n523gat), .A1(n522gat), .A2(n356gat) );
  NOR2_X1 NOR2_396( .ZN(n634gat), .A1(n418gat), .A2(n521gat) );
  NOR2_X1 NOR2_397( .ZN(n414gat), .A1(n411gat), .A2(n415gat) );
  NOR3_X1 NOR3_236( .ZN(n635gat), .A1(n639gat), .A2(n634gat), .A3(n414gat) );
  NOR2_X1 NOR2_398( .ZN(n1100gat), .A1(n1297gat), .A2(n1111gat) );
  NOR3_X1 NOR3_237( .ZN(n630gat), .A1(n634gat), .A2(n523gat), .A3(n524gat) );
  NOR2_X1 NOR2_399( .ZN(n994gat), .A1(n1112gat), .A2(n882gat) );
  NOR3_X1 NOR3_238( .ZN(n629gat), .A1(n414gat), .A2(n634gat), .A3(n523gat) );
  NOR2_X1 NOR2_400( .ZN(n989gat), .A1(n721gat), .A2(n741gat) );
  NOR3_X1 NOR3_239( .ZN(n632gat), .A1(n414gat), .A2(n523gat), .A3(n633gat) );
  NOR2_X1 NOR2_401( .ZN(n880gat), .A1(n926gat), .A2(n566gat) );
  NOR3_X1 NOR3_240( .ZN(n636gat), .A1(n414gat), .A2(n633gat), .A3(n639gat) );
  NOR2_X1 NOR2_402( .ZN(n801gat), .A1(n672gat), .A2(n670gat) );
  NOR2_X1 NOR2_403( .ZN(n879gat), .A1(n2931gat), .A2(n801gat) );
  NOR2_X1 NOR2_404( .ZN(n1003gat), .A1(n420gat), .A2(n879gat) );
  NOR2_X1 NOR2_405( .ZN(n1255gat), .A1(n1123gat), .A2(n1225gat) );
  NOR2_X1 NOR2_406( .ZN(n1012gat), .A1(n1007gat), .A2(n918gat) );
  NOR2_X1 NOR2_407( .ZN(n905gat), .A1(n625gat), .A2(n1006gat) );
  NOR2_X1 NOR2_408( .ZN(n1009gat), .A1(n1255gat), .A2(n2943gat) );
  NOR2_X1 NOR2_409( .ZN(n409gat), .A1(n406gat), .A2(n407gat) );
  NOR2_X1 NOR2_410( .ZN(n292gat), .A1(n415gat), .A2(n356gat) );
  NOR2_X1 NOR2_411( .ZN(n291gat), .A1(n290gat), .A2(n292gat) );
  NOR2_X1 NOR2_412( .ZN(n419gat), .A1(n409gat), .A2(n291gat) );
  NOR2_X1 NOR2_413( .ZN(n902gat), .A1(n1009gat), .A2(n419gat) );
  NOR2_X1 NOR2_414( .ZN(n1099gat), .A1(n1111gat), .A2(n1293gat) );
  NOR2_X1 NOR2_415( .ZN(n998gat), .A1(n725gat), .A2(n741gat) );
  NOR2_X1 NOR2_416( .ZN(n995gat), .A1(n823gat), .A2(n1112gat) );
  NOR2_X1 NOR2_417( .ZN(n980gat), .A1(n875gat), .A2(n926gat) );
  NOR2_X1 NOR2_418( .ZN(n1001gat), .A1(n420gat), .A2(n1002gat) );
  NOR2_X1 NOR2_419( .ZN(n1175gat), .A1(n621gat), .A2(n1006gat) );
  NOR2_X1 NOR2_420( .ZN(n1174gat), .A1(n845gat), .A2(n1007gat) );
  NOR2_X1 NOR2_421( .ZN(n1243gat), .A1(n1281gat), .A2(n1123gat) );
  NOR2_X1 NOR2_422( .ZN(n1171gat), .A1(n2960gat), .A2(n1243gat) );
  NOR2_X1 NOR2_423( .ZN(n999gat), .A1(n419gat), .A2(n1171gat) );
  NOR2_X1 NOR2_424( .ZN(n1244gat), .A1(n1123gat), .A2(n1134gat) );
  NOR2_X1 NOR2_425( .ZN(n1323gat), .A1(n1007gat), .A2(n401gat) );
  NOR2_X1 NOR2_426( .ZN(n1264gat), .A1(n1006gat), .A2(n617gat) );
  NOR2_X2 NOR2_427( .ZN(n1265gat), .A1(n1244gat), .A2(n2969gat) );
  NOR2_X1 NOR2_428( .ZN(n892gat), .A1(n419gat), .A2(n1265gat) );
  NOR2_X1 NOR2_429( .ZN(n981gat), .A1(n926gat), .A2(n873gat) );
  NOR2_X1 NOR2_430( .ZN(n890gat), .A1(n741gat), .A2(n702gat) );
  NOR2_X1 NOR2_431( .ZN(n889gat), .A1(n1111gat), .A2(n1079gat) );
  NOR2_X1 NOR2_432( .ZN(n886gat), .A1(n683gat), .A2(n1112gat) );
  NOR2_X1 NOR2_433( .ZN(n891gat), .A1(n420gat), .A2(n888gat) );
  NOR2_X1 NOR2_434( .ZN(n904gat), .A1(n1006gat), .A2(n490gat) );
  NOR2_X1 NOR2_435( .ZN(n903gat), .A1(n1007gat), .A2(n397gat) );
  NOR2_X1 NOR2_436( .ZN(n1254gat), .A1(n1123gat), .A2(n1044gat) );
  NOR2_X1 NOR2_437( .ZN(n1008gat), .A1(n2942gat), .A2(n1254gat) );
  NOR2_X1 NOR2_438( .ZN(n900gat), .A1(n419gat), .A2(n1008gat) );
  NOR2_X1 NOR2_439( .ZN(n1152gat), .A1(n926gat), .A2(n1150gat) );
  NOR2_X1 NOR2_440( .ZN(n1092gat), .A1(n1147gat), .A2(n1111gat) );
  NOR2_X1 NOR2_441( .ZN(n997gat), .A1(n741gat), .A2(n393gat) );
  NOR2_X1 NOR2_442( .ZN(n993gat), .A1(n1112gat), .A2(n698gat) );
  NOR2_X1 NOR2_443( .ZN(n895gat), .A1(n420gat), .A2(n898gat) );
  NOR2_X1 NOR2_444( .ZN(n1094gat), .A1(n1112gat), .A2(n583gat) );
  NOR2_X1 NOR2_445( .ZN(n1093gat), .A1(n1111gat), .A2(n864gat) );
  NOR2_X1 NOR2_446( .ZN(n988gat), .A1(n340gat), .A2(n741gat) );
  NOR2_X1 NOR2_447( .ZN(n984gat), .A1(n926gat), .A2(n983gat) );
  NOR2_X1 NOR2_448( .ZN(n1178gat), .A1(n420gat), .A2(n1179gat) );
  NOR2_X1 NOR2_449( .ZN(n1267gat), .A1(n613gat), .A2(n1006gat) );
  NOR2_X1 NOR2_450( .ZN(n1257gat), .A1(n1007gat), .A2(n274gat) );
  NOR2_X1 NOR2_451( .ZN(n1253gat), .A1(n930gat), .A2(n1123gat) );
  NOR2_X1 NOR2_452( .ZN(n1266gat), .A1(n2965gat), .A2(n1253gat) );
  NOR2_X1 NOR2_453( .ZN(n1116gat), .A1(n419gat), .A2(n1266gat) );
  NOR2_X1 NOR2_454( .ZN(n1375gat), .A1(n1006gat), .A2(n706gat) );
  NOR2_X1 NOR2_455( .ZN(n1324gat), .A1(n164gat), .A2(n1007gat) );
  NOR2_X1 NOR2_456( .ZN(n1200gat), .A1(n1120gat), .A2(n1123gat) );
  NOR2_X1 NOR2_457( .ZN(n1172gat), .A1(n2961gat), .A2(n1200gat) );
  NOR2_X1 NOR2_458( .ZN(n899gat), .A1(n419gat), .A2(n1172gat) );
  NOR2_X1 NOR2_459( .ZN(n1091gat), .A1(n1111gat), .A2(n956gat) );
  NOR2_X1 NOR2_460( .ZN(n1088gat), .A1(n1085gat), .A2(n926gat) );
  NOR2_X1 NOR2_461( .ZN(n992gat), .A1(n815gat), .A2(n1112gat) );
  NOR2_X1 NOR2_462( .ZN(n987gat), .A1(n741gat), .A2(n159gat) );
  NOR2_X1 NOR2_463( .ZN(n896gat), .A1(n897gat), .A2(n420gat) );
  NOR2_X1 NOR2_464( .ZN(n1262gat), .A1(n837gat), .A2(n1006gat) );
  NOR2_X1 NOR2_465( .ZN(n1260gat), .A1(n1007gat), .A2(n278gat) );
  NOR2_X1 NOR2_466( .ZN(n1251gat), .A1(n1123gat), .A2(n1071gat) );
  NOR2_X1 NOR2_467( .ZN(n1259gat), .A1(n2967gat), .A2(n1251gat) );
  NOR2_X1 NOR2_468( .ZN(n901gat), .A1(n419gat), .A2(n1259gat) );
  NOR2_X1 NOR2_469( .ZN(n1098gat), .A1(n336gat), .A2(n741gat) );
  NOR2_X1 NOR2_470( .ZN(n1090gat), .A1(n1111gat), .A2(n860gat) );
  NOR2_X1 NOR2_471( .ZN(n986gat), .A1(n985gat), .A2(n926gat) );
  NOR2_X1 NOR2_472( .ZN(n885gat), .A1(n579gat), .A2(n1112gat) );
  NOR2_X1 NOR2_473( .ZN(n893gat), .A1(n894gat), .A2(n420gat) );
  NOR2_X1 NOR2_474( .ZN(n1097gat), .A1(n270gat), .A2(n741gat) );
  NOR2_X1 NOR2_475( .ZN(n1089gat), .A1(n1067gat), .A2(n1111gat) );
  NOR2_X1 NOR2_476( .ZN(n1087gat), .A1(n926gat), .A2(n1084gat) );
  NOR2_X1 NOR2_477( .ZN(n991gat), .A1(n1112gat), .A2(n679gat) );
  NOR2_X1 NOR2_478( .ZN(n1177gat), .A1(n1180gat), .A2(n420gat) );
  NOR2_X2 NOR2_479( .ZN(n1212gat), .A1(n1123gat), .A2(n1034gat) );
  NOR2_X2 NOR2_480( .ZN(n1326gat), .A1(n1007gat), .A2(n282gat) );
  NOR2_X1 NOR2_481( .ZN(n1261gat), .A1(n833gat), .A2(n1006gat) );
  NOR2_X1 NOR2_482( .ZN(n1263gat), .A1(n1212gat), .A2(n2968gat) );
  NOR2_X1 NOR2_483( .ZN(n1115gat), .A1(n1263gat), .A2(n419gat) );
  NOR2_X1 NOR2_484( .ZN(n977gat), .A1(n670gat), .A2(n671gat) );
  NOR3_X1 NOR3_241( .ZN(n631gat), .A1(n523gat), .A2(n633gat), .A3(n524gat) );
  NOR2_X1 NOR2_485( .ZN(n1096gat), .A1(n819gat), .A2(n1112gat) );
  NOR2_X1 NOR2_486( .ZN(n1095gat), .A1(n1240gat), .A2(n1111gat) );
  NOR2_X1 NOR2_487( .ZN(n990gat), .A1(n841gat), .A2(n741gat) );
  NOR2_X1 NOR2_488( .ZN(n979gat), .A1(n1601gat), .A2(n926gat) );
  NOR2_X1 NOR2_489( .ZN(n978gat), .A1(n2944gat), .A2(n2945gat) );
  NOR2_X1 NOR2_490( .ZN(n1004gat), .A1(n978gat), .A2(n420gat) );
  NOR2_X1 NOR2_491( .ZN(n1199gat), .A1(n1123gat), .A2(n1284gat) );
  NOR2_X1 NOR2_492( .ZN(n1176gat), .A1(n829gat), .A2(n1006gat) );
  NOR2_X1 NOR2_493( .ZN(n1173gat), .A1(n1007gat), .A2(n1025gat) );
  NOR2_X1 NOR2_494( .ZN(n1252gat), .A1(n1199gat), .A2(n2962gat) );
  NOR2_X1 NOR2_495( .ZN(n1000gat), .A1(n419gat), .A2(n1252gat) );
  NOR2_X1 NOR2_496( .ZN(n1029gat), .A1(n978gat), .A2(n455gat) );
  NOR2_X1 NOR2_497( .ZN(n1028gat), .A1(n455gat), .A2(n879gat) );
  NOR2_X1 NOR2_498( .ZN(n1031gat), .A1(n1002gat), .A2(n455gat) );
  NOR2_X1 NOR2_499( .ZN(n1030gat), .A1(n455gat), .A2(n888gat) );
  NOR2_X1 NOR2_500( .ZN(n1011gat), .A1(n455gat), .A2(n898gat) );
  NOR2_X1 NOR2_501( .ZN(n1181gat), .A1(n455gat), .A2(n1179gat) );
  NOR2_X1 NOR2_502( .ZN(n1010gat), .A1(n897gat), .A2(n455gat) );
  NOR2_X1 NOR2_503( .ZN(n1005gat), .A1(n894gat), .A2(n455gat) );
  NOR2_X1 NOR2_504( .ZN(n1182gat), .A1(n1180gat), .A2(n455gat) );
  NOR2_X1 NOR2_505( .ZN(n1757gat), .A1(n1773gat), .A2(n1769gat) );
  NOR2_X1 NOR2_506( .ZN(n1745gat), .A1(n1869gat), .A2(n1757gat) );
  NOR2_X1 NOR2_507( .ZN(n73gat), .A1(n67gat), .A2(n2784gat) );
  NOR2_X1 NOR2_508( .ZN(n70gat), .A1(n71gat), .A2(n2720gat) );
  NOR2_X2 NOR2_509( .ZN(n77gat), .A1(n76gat), .A2(n2784gat) );
  NOR2_X1 NOR2_510( .ZN(n13gat), .A1(n2720gat), .A2(n14gat) );

endmodule
