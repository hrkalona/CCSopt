// Verilog
// c1908
// Ninputs 33
// Noutputs 25
// NtotalGates 880
// NOT1 277
// NAND2 347
// BUFF1 162
// AND2 30
// AND3 12
// NAND4 2
// NAND3 1
// NAND8 3
// AND4 2
// NAND5 24
// AND5 16
// AND8 3
// NOR2 1

module c1908(N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,N31,N34,N37,N40,N43,N46,N49,N53,
  N56,N60,N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,N94,N99,N104,N2753,N2754,N2755,
  N2756,N2762,N2767,N2768,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,N2889,
  N2890,N2891,N2892,N2899);
input N1,N4,N7,N10,N13,N16,N19,N22,N25,N28,N31,N34,N37,N40,N43,N46,N49,N53,N56,N60,
  N63,N66,N69,N72,N76,N79,N82,N85,N88,N91,N94,N99,N104;
output N2753,N2754,N2755,N2756,N2762,N2767,N2768,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2811,N2886,N2887,N2888,
  N2889,N2890,N2891,N2892,N2899;

  wire N190,N194,N197,N201,N206,N209,N212,N216,N220,N225,N229,N232,N235,N239,N243,N247,
    N251,N252,N253,N256,N257,N260,N263,N266,N269,N272,N275,N276,N277,N280,N283,N290,
    N297,N300,N303,N306,N313,N316,N319,N326,N331,N338,N343,N346,N349,N352,N355,N358,
    N361,N364,N367,N370,N373,N376,N379,N382,N385,N388,N534,N535,N536,N537,N538,N539,
    N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
    N556,N559,N562,N565,N568,N571,N574,N577,N580,N583,N586,N589,N592,N595,N598,N601,
    N602,N603,N608,N612,N616,N619,N622,N625,N628,N631,N634,N637,N640,N643,N646,N649,
    N652,N655,N658,N661,N664,N667,N670,N673,N676,N679,N682,N685,N688,N691,N694,N697,
    N700,N703,N706,N709,N712,N715,N718,N721,N724,N727,N730,N733,N736,N739,N742,N745,
    N748,N751,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
    N903,N907,N910,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N926,N935,
    N938,N939,N942,N943,N946,N947,N950,N951,N954,N955,N958,N959,N962,N965,N968,N969,
    N972,N973,N976,N977,N980,N981,N984,N985,N988,N989,N990,N991,N992,N993,N994,N997,
    N998,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1013,N1016,N1019,N1022,N1025,
    N1028,N1031,N1034,N1037,N1040,N1043,N1046,N1049,N1054,N1055,N1063,N1064,N1067,N1068,N1119,N1120,
    N1121,N1122,N1128,N1129,N1130,N1131,N1132,N1133,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,
    N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1167,N1168,N1171,N1188,N1205,N1206,N1207,
    N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,
    N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1235,N1238,N1239,N1240,N1241,N1242,N1243,
    N1246,N1249,N1252,N1255,N1258,N1261,N1264,N1267,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
    N1317,N1318,N1319,N1322,N1327,N1328,N1334,N1344,N1345,N1346,N1348,N1349,N1350,N1351,N1352,N1355,
    N1358,N1361,N1364,N1367,N1370,N1373,N1376,N1379,N1383,N1386,N1387,N1388,N1389,N1390,N1393,N1396,
    N1397,N1398,N1399,N1409,N1412,N1413,N1416,N1419,N1433,N1434,N1438,N1439,N1440,N1443,N1444,N1445,
    N1446,N1447,N1448,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,
    N1464,N1468,N1469,N1470,N1471,N1472,N1475,N1476,N1478,N1481,N1484,N1487,N1488,N1489,N1490,N1491,
    N1492,N1493,N1494,N1495,N1496,N1498,N1499,N1500,N1501,N1504,N1510,N1513,N1514,N1517,N1520,N1521,
    N1522,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1534,N1537,N1540,N1546,N1554,N1557,N1561,N1567,
    N1568,N1569,N1571,N1576,N1588,N1591,N1593,N1594,N1595,N1596,N1600,N1603,N1606,N1609,N1612,N1615,
    N1620,N1623,N1635,N1636,N1638,N1639,N1640,N1643,N1647,N1651,N1658,N1661,N1664,N1671,N1672,N1675,
    N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1685,N1688,N1697,N1701,N1706,N1707,N1708,N1709,N1710,
    N1711,N1712,N1713,N1714,N1717,N1720,N1721,N1723,N1727,N1728,N1730,N1731,N1734,N1740,N1741,N1742,
    N1746,N1747,N1748,N1751,N1759,N1761,N1762,N1763,N1764,N1768,N1769,N1772,N1773,N1774,N1777,N1783,
    N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1795,N1796,N1798,N1801,N1802,N1807,N1808,N1809,N1810,
    N1812,N1815,N1818,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1830,N1837,N1838,N1841,N1848,N1849,
    N1850,N1852,N1855,N1856,N1857,N1858,N1864,N1865,N1866,N1869,N1872,N1875,N1878,N1879,N1882,N1883,
    N1884,N1885,N1889,N1895,N1896,N1897,N1898,N1902,N1910,N1911,N1912,N1913,N1915,N1919,N1920,N1921,
    N1922,N1923,N1924,N1927,N1930,N1933,N1936,N1937,N1938,N1941,N1942,N1944,N1947,N1950,N1953,N1958,
    N1961,N1965,N1968,N1975,N1976,N1977,N1978,N1979,N1980,N1985,N1987,N1999,N2000,N2002,N2003,N2004,
    N2005,N2006,N2007,N2008,N2009,N2012,N2013,N2014,N2015,N2016,N2018,N2019,N2020,N2021,N2022,N2023,
    N2024,N2025,N2026,N2027,N2030,N2033,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2047,N2052,N2055,
    N2060,N2061,N2062,N2067,N2068,N2071,N2076,N2077,N2078,N2081,N2086,N2089,N2104,N2119,N2129,N2143,
    N2148,N2151,N2196,N2199,N2202,N2205,N2214,N2215,N2216,N2217,N2222,N2223,N2224,N2225,N2226,N2227,
    N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2240,N2241,N2244,N2245,N2250,N2253,
    N2256,N2257,N2260,N2263,N2266,N2269,N2272,N2279,N2286,N2297,N2315,N2326,N2340,N2353,N2361,N2375,
    N2384,N2385,N2386,N2426,N2427,N2537,N2540,N2543,N2546,N2549,N2552,N2555,N2558,N2561,N2564,N2567,
    N2570,N2573,N2576,N2594,N2597,N2600,N2603,N2606,N2611,N2614,N2617,N2620,N2627,N2628,N2629,N2630,
    N2631,N2632,N2633,N2634,N2639,N2642,N2645,N2648,N2651,N2655,N2658,N2661,N2664,N2669,N2670,N2671,
    N2672,N2673,N2674,N2675,N2676,N2682,N2683,N2688,N2689,N2690,N2691,N2710,N2720,N2721,N2722,N2723,
    N2724,N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,
    N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2750,N2757,N2758,N2759,N2760,N2761,N2763,N2764,
    N2765,N2766,N2773,N2776,N2788,N2789,N2800,N2807,N2808,N2809,N2810,N2812,N2815,N2818,N2821,N2824,
    N2827,N2828,N2829,N2843,N2846,N2850,N2851,N2852,N2853,N2854,N2857,N2858,N2859,N2860,N2861,N2862,
    N2863,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,
    N2881,N2882,N2883,N2895,N2896,N2897,N2898,extra0,extra1,extra2,extra3,extra4,extra5,extra6,extra7,extra8,
    extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,extra17,extra18,extra19,extra20,extra21,extra22,extra23,extra24,
    extra25,extra26,extra27,extra28,extra29,extra30,extra31,extra32,extra33,extra34,extra35,extra36,extra37,extra38,extra39,extra40,
    extra41,extra42,extra43,extra44,extra45,extra46,extra47,extra48,extra49,extra50,extra51;

  INV_X4 NOT1_1( .ZN(N190), .A(N1) );
  INV_X1 NOT1_2( .ZN(N194), .A(N4) );
  INV_X1 NOT1_3( .ZN(N197), .A(N7) );
  INV_X1 NOT1_4( .ZN(N201), .A(N10) );
  INV_X1 NOT1_5( .ZN(N206), .A(N13) );
  INV_X1 NOT1_6( .ZN(N209), .A(N16) );
  INV_X1 NOT1_7( .ZN(N212), .A(N19) );
  INV_X1 NOT1_8( .ZN(N216), .A(N22) );
  INV_X1 NOT1_9( .ZN(N220), .A(N25) );
  INV_X1 NOT1_10( .ZN(N225), .A(N28) );
  INV_X4 NOT1_11( .ZN(N229), .A(N31) );
  INV_X1 NOT1_12( .ZN(N232), .A(N34) );
  INV_X1 NOT1_13( .ZN(N235), .A(N37) );
  INV_X1 NOT1_14( .ZN(N239), .A(N40) );
  INV_X1 NOT1_15( .ZN(N243), .A(N43) );
  INV_X1 NOT1_16( .ZN(N247), .A(N46) );
  NAND2_X1 NAND2_17( .ZN(N251), .A1(N63), .A2(N88) );
  NAND2_X1 NAND2_18( .ZN(N252), .A1(N66), .A2(N91) );
  INV_X1 NOT1_19( .ZN(N253), .A(N72) );
  INV_X1 NOT1_20( .ZN(N256), .A(N72) );
  BUF_X2 BUFF1_21( .Z(N257), .A(N69) );
  BUF_X1 BUFF1_22( .Z(N260), .A(N69) );
  INV_X4 NOT1_23( .ZN(N263), .A(N76) );
  INV_X1 NOT1_24( .ZN(N266), .A(N79) );
  INV_X1 NOT1_25( .ZN(N269), .A(N82) );
  INV_X1 NOT1_26( .ZN(N272), .A(N85) );
  INV_X1 NOT1_27( .ZN(N275), .A(N104) );
  INV_X1 NOT1_28( .ZN(N276), .A(N104) );
  INV_X1 NOT1_29( .ZN(N277), .A(N88) );
  INV_X1 NOT1_30( .ZN(N280), .A(N91) );
  BUF_X1 BUFF1_31( .Z(N283), .A(N94) );
  INV_X1 NOT1_32( .ZN(N290), .A(N94) );
  BUF_X1 BUFF1_33( .Z(N297), .A(N94) );
  INV_X1 NOT1_34( .ZN(N300), .A(N94) );
  BUF_X1 BUFF1_35( .Z(N303), .A(N99) );
  INV_X1 NOT1_36( .ZN(N306), .A(N99) );
  INV_X1 NOT1_37( .ZN(N313), .A(N99) );
  BUF_X1 BUFF1_38( .Z(N316), .A(N104) );
  INV_X1 NOT1_39( .ZN(N319), .A(N104) );
  BUF_X1 BUFF1_40( .Z(N326), .A(N104) );
  BUF_X1 BUFF1_41( .Z(N331), .A(N104) );
  INV_X1 NOT1_42( .ZN(N338), .A(N104) );
  BUF_X1 BUFF1_43( .Z(N343), .A(N1) );
  BUF_X1 BUFF1_44( .Z(N346), .A(N4) );
  BUF_X1 BUFF1_45( .Z(N349), .A(N7) );
  BUF_X1 BUFF1_46( .Z(N352), .A(N10) );
  BUF_X1 BUFF1_47( .Z(N355), .A(N13) );
  BUF_X1 BUFF1_48( .Z(N358), .A(N16) );
  BUF_X1 BUFF1_49( .Z(N361), .A(N19) );
  BUF_X1 BUFF1_50( .Z(N364), .A(N22) );
  BUF_X1 BUFF1_51( .Z(N367), .A(N25) );
  BUF_X1 BUFF1_52( .Z(N370), .A(N28) );
  BUF_X1 BUFF1_53( .Z(N373), .A(N31) );
  BUF_X1 BUFF1_54( .Z(N376), .A(N34) );
  BUF_X1 BUFF1_55( .Z(N379), .A(N37) );
  BUF_X1 BUFF1_56( .Z(N382), .A(N40) );
  BUF_X1 BUFF1_57( .Z(N385), .A(N43) );
  BUF_X1 BUFF1_58( .Z(N388), .A(N46) );
  INV_X1 NOT1_59( .ZN(N534), .A(N343) );
  INV_X1 NOT1_60( .ZN(N535), .A(N346) );
  INV_X4 NOT1_61( .ZN(N536), .A(N349) );
  INV_X1 NOT1_62( .ZN(N537), .A(N352) );
  INV_X1 NOT1_63( .ZN(N538), .A(N355) );
  INV_X1 NOT1_64( .ZN(N539), .A(N358) );
  INV_X1 NOT1_65( .ZN(N540), .A(N361) );
  INV_X1 NOT1_66( .ZN(N541), .A(N364) );
  INV_X1 NOT1_67( .ZN(N542), .A(N367) );
  INV_X1 NOT1_68( .ZN(N543), .A(N370) );
  INV_X1 NOT1_69( .ZN(N544), .A(N373) );
  INV_X1 NOT1_70( .ZN(N545), .A(N376) );
  INV_X1 NOT1_71( .ZN(N546), .A(N379) );
  INV_X1 NOT1_72( .ZN(N547), .A(N382) );
  INV_X1 NOT1_73( .ZN(N548), .A(N385) );
  INV_X1 NOT1_74( .ZN(N549), .A(N388) );
  NAND2_X1 NAND2_75( .ZN(N550), .A1(N306), .A2(N331) );
  NAND2_X1 NAND2_76( .ZN(N551), .A1(N306), .A2(N331) );
  NAND2_X1 NAND2_77( .ZN(N552), .A1(N306), .A2(N331) );
  NAND2_X1 NAND2_78( .ZN(N553), .A1(N306), .A2(N331) );
  NAND2_X1 NAND2_79( .ZN(N554), .A1(N306), .A2(N331) );
  NAND2_X1 NAND2_80( .ZN(N555), .A1(N306), .A2(N331) );
  BUF_X1 BUFF1_81( .Z(N556), .A(N190) );
  BUF_X1 BUFF1_82( .Z(N559), .A(N194) );
  BUF_X1 BUFF1_83( .Z(N562), .A(N206) );
  BUF_X1 BUFF1_84( .Z(N565), .A(N209) );
  BUF_X1 BUFF1_85( .Z(N568), .A(N225) );
  BUF_X1 BUFF1_86( .Z(N571), .A(N243) );
  AND2_X1 AND2_87( .ZN(N574), .A1(N63), .A2(N319) );
  BUF_X2 BUFF1_88( .Z(N577), .A(N220) );
  BUF_X2 BUFF1_89( .Z(N580), .A(N229) );
  BUF_X1 BUFF1_90( .Z(N583), .A(N232) );
  AND2_X1 AND2_91( .ZN(N586), .A1(N66), .A2(N319) );
  BUF_X1 BUFF1_92( .Z(N589), .A(N239) );
  AND3_X1 AND3_93( .ZN(N592), .A1(N49), .A2(N253), .A3(N319) );
  BUF_X1 BUFF1_94( .Z(N595), .A(N247) );
  BUF_X1 BUFF1_95( .Z(N598), .A(N239) );
  NAND2_X1 NAND2_96( .ZN(N601), .A1(N326), .A2(N277) );
  NAND2_X1 NAND2_97( .ZN(N602), .A1(N326), .A2(N280) );
  NAND2_X1 NAND2_98( .ZN(N603), .A1(N260), .A2(N72) );
  NAND2_X1 NAND2_99( .ZN(N608), .A1(N260), .A2(N300) );
  NAND2_X2 NAND2_100( .ZN(N612), .A1(N256), .A2(N300) );
  BUF_X1 BUFF1_101( .Z(N616), .A(N201) );
  BUF_X1 BUFF1_102( .Z(N619), .A(N216) );
  BUF_X1 BUFF1_103( .Z(N622), .A(N220) );
  BUF_X1 BUFF1_104( .Z(N625), .A(N239) );
  BUF_X1 BUFF1_105( .Z(N628), .A(N190) );
  BUF_X1 BUFF1_106( .Z(N631), .A(N190) );
  BUF_X1 BUFF1_107( .Z(N634), .A(N194) );
  BUF_X1 BUFF1_108( .Z(N637), .A(N229) );
  BUF_X1 BUFF1_109( .Z(N640), .A(N197) );
  AND3_X1 AND3_110( .ZN(N643), .A1(N56), .A2(N257), .A3(N319) );
  BUF_X1 BUFF1_111( .Z(N646), .A(N232) );
  BUF_X1 BUFF1_112( .Z(N649), .A(N201) );
  BUF_X1 BUFF1_113( .Z(N652), .A(N235) );
  AND3_X1 AND3_114( .ZN(N655), .A1(N60), .A2(N257), .A3(N319) );
  BUF_X1 BUFF1_115( .Z(N658), .A(N263) );
  BUF_X1 BUFF1_116( .Z(N661), .A(N263) );
  BUF_X1 BUFF1_117( .Z(N664), .A(N266) );
  BUF_X1 BUFF1_118( .Z(N667), .A(N266) );
  BUF_X1 BUFF1_119( .Z(N670), .A(N269) );
  BUF_X1 BUFF1_120( .Z(N673), .A(N269) );
  BUF_X1 BUFF1_121( .Z(N676), .A(N272) );
  BUF_X1 BUFF1_122( .Z(N679), .A(N272) );
  AND2_X1 AND2_123( .ZN(N682), .A1(N251), .A2(N316) );
  AND2_X1 AND2_124( .ZN(N685), .A1(N252), .A2(N316) );
  BUF_X1 BUFF1_125( .Z(N688), .A(N197) );
  BUF_X1 BUFF1_126( .Z(N691), .A(N197) );
  BUF_X1 BUFF1_127( .Z(N694), .A(N212) );
  BUF_X1 BUFF1_128( .Z(N697), .A(N212) );
  BUF_X1 BUFF1_129( .Z(N700), .A(N247) );
  BUF_X1 BUFF1_130( .Z(N703), .A(N247) );
  BUF_X1 BUFF1_131( .Z(N706), .A(N235) );
  BUF_X1 BUFF1_132( .Z(N709), .A(N235) );
  BUF_X1 BUFF1_133( .Z(N712), .A(N201) );
  BUF_X1 BUFF1_134( .Z(N715), .A(N201) );
  BUF_X1 BUFF1_135( .Z(N718), .A(N206) );
  BUF_X1 BUFF1_136( .Z(N721), .A(N216) );
  AND3_X1 AND3_137( .ZN(N724), .A1(N53), .A2(N253), .A3(N319) );
  BUF_X1 BUFF1_138( .Z(N727), .A(N243) );
  BUF_X1 BUFF1_139( .Z(N730), .A(N220) );
  BUF_X1 BUFF1_140( .Z(N733), .A(N220) );
  BUF_X1 BUFF1_141( .Z(N736), .A(N209) );
  BUF_X1 BUFF1_142( .Z(N739), .A(N216) );
  BUF_X1 BUFF1_143( .Z(N742), .A(N225) );
  BUF_X1 BUFF1_144( .Z(N745), .A(N243) );
  BUF_X1 BUFF1_145( .Z(N748), .A(N212) );
  BUF_X1 BUFF1_146( .Z(N751), .A(N225) );
  INV_X4 NOT1_147( .ZN(N886), .A(N682) );
  INV_X4 NOT1_148( .ZN(N887), .A(N685) );
  INV_X1 NOT1_149( .ZN(N888), .A(N616) );
  INV_X1 NOT1_150( .ZN(N889), .A(N619) );
  INV_X1 NOT1_151( .ZN(N890), .A(N622) );
  INV_X1 NOT1_152( .ZN(N891), .A(N625) );
  INV_X1 NOT1_153( .ZN(N892), .A(N631) );
  INV_X1 NOT1_154( .ZN(N893), .A(N643) );
  INV_X1 NOT1_155( .ZN(N894), .A(N649) );
  INV_X1 NOT1_156( .ZN(N895), .A(N652) );
  INV_X1 NOT1_157( .ZN(N896), .A(N655) );
  AND2_X1 AND2_158( .ZN(N897), .A1(N49), .A2(N612) );
  AND2_X1 AND2_159( .ZN(N898), .A1(N56), .A2(N608) );
  NAND2_X1 NAND2_160( .ZN(N899), .A1(N53), .A2(N612) );
  NAND2_X1 NAND2_161( .ZN(N903), .A1(N60), .A2(N608) );
  NAND2_X1 NAND2_162( .ZN(N907), .A1(N49), .A2(N612) );
  NAND2_X1 NAND2_163( .ZN(N910), .A1(N56), .A2(N608) );
  INV_X1 NOT1_164( .ZN(N913), .A(N661) );
  INV_X1 NOT1_165( .ZN(N914), .A(N658) );
  INV_X1 NOT1_166( .ZN(N915), .A(N667) );
  INV_X1 NOT1_167( .ZN(N916), .A(N664) );
  INV_X1 NOT1_168( .ZN(N917), .A(N673) );
  INV_X1 NOT1_169( .ZN(N918), .A(N670) );
  INV_X1 NOT1_170( .ZN(N919), .A(N679) );
  INV_X1 NOT1_171( .ZN(N920), .A(N676) );
  NAND4_X1 NAND4_172( .ZN(N921), .A1(N277), .A2(N297), .A3(N326), .A4(N603) );
  NAND4_X1 NAND4_173( .ZN(N922), .A1(N280), .A2(N297), .A3(N326), .A4(N603) );
  NAND3_X1 NAND3_174( .ZN(N923), .A1(N303), .A2(N338), .A3(N603) );
  AND3_X1 AND3_175( .ZN(N926), .A1(N303), .A2(N338), .A3(N603) );
  BUF_X1 BUFF1_176( .Z(N935), .A(N556) );
  INV_X2 NOT1_177( .ZN(N938), .A(N688) );
  BUF_X1 BUFF1_178( .Z(N939), .A(N556) );
  INV_X2 NOT1_179( .ZN(N942), .A(N691) );
  BUF_X1 BUFF1_180( .Z(N943), .A(N562) );
  INV_X1 NOT1_181( .ZN(N946), .A(N694) );
  BUF_X1 BUFF1_182( .Z(N947), .A(N562) );
  INV_X1 NOT1_183( .ZN(N950), .A(N697) );
  BUF_X1 BUFF1_184( .Z(N951), .A(N568) );
  INV_X1 NOT1_185( .ZN(N954), .A(N700) );
  BUF_X1 BUFF1_186( .Z(N955), .A(N568) );
  INV_X1 NOT1_187( .ZN(N958), .A(N703) );
  BUF_X1 BUFF1_188( .Z(N959), .A(N574) );
  BUF_X1 BUFF1_189( .Z(N962), .A(N574) );
  BUF_X1 BUFF1_190( .Z(N965), .A(N580) );
  INV_X1 NOT1_191( .ZN(N968), .A(N706) );
  BUF_X1 BUFF1_192( .Z(N969), .A(N580) );
  INV_X1 NOT1_193( .ZN(N972), .A(N709) );
  BUF_X1 BUFF1_194( .Z(N973), .A(N586) );
  INV_X1 NOT1_195( .ZN(N976), .A(N712) );
  BUF_X2 BUFF1_196( .Z(N977), .A(N586) );
  INV_X1 NOT1_197( .ZN(N980), .A(N715) );
  BUF_X2 BUFF1_198( .Z(N981), .A(N592) );
  INV_X1 NOT1_199( .ZN(N984), .A(N628) );
  BUF_X1 BUFF1_200( .Z(N985), .A(N592) );
  INV_X1 NOT1_201( .ZN(N988), .A(N718) );
  INV_X1 NOT1_202( .ZN(N989), .A(N721) );
  INV_X1 NOT1_203( .ZN(N990), .A(N634) );
  INV_X1 NOT1_204( .ZN(N991), .A(N724) );
  INV_X2 NOT1_205( .ZN(N992), .A(N727) );
  INV_X2 NOT1_206( .ZN(N993), .A(N637) );
  BUF_X1 BUFF1_207( .Z(N994), .A(N595) );
  INV_X1 NOT1_208( .ZN(N997), .A(N730) );
  BUF_X1 BUFF1_209( .Z(N998), .A(N595) );
  INV_X1 NOT1_210( .ZN(N1001), .A(N733) );
  INV_X1 NOT1_211( .ZN(N1002), .A(N736) );
  INV_X1 NOT1_212( .ZN(N1003), .A(N739) );
  INV_X1 NOT1_213( .ZN(N1004), .A(N640) );
  INV_X1 NOT1_214( .ZN(N1005), .A(N742) );
  INV_X1 NOT1_215( .ZN(N1006), .A(N745) );
  INV_X1 NOT1_216( .ZN(N1007), .A(N646) );
  INV_X1 NOT1_217( .ZN(N1008), .A(N748) );
  INV_X1 NOT1_218( .ZN(N1009), .A(N751) );
  BUF_X1 BUFF1_219( .Z(N1010), .A(N559) );
  BUF_X1 BUFF1_220( .Z(N1013), .A(N559) );
  BUF_X1 BUFF1_221( .Z(N1016), .A(N565) );
  BUF_X1 BUFF1_222( .Z(N1019), .A(N565) );
  BUF_X1 BUFF1_223( .Z(N1022), .A(N571) );
  BUF_X1 BUFF1_224( .Z(N1025), .A(N571) );
  BUF_X1 BUFF1_225( .Z(N1028), .A(N577) );
  BUF_X1 BUFF1_226( .Z(N1031), .A(N577) );
  BUF_X1 BUFF1_227( .Z(N1034), .A(N583) );
  BUF_X1 BUFF1_228( .Z(N1037), .A(N583) );
  BUF_X1 BUFF1_229( .Z(N1040), .A(N589) );
  BUF_X1 BUFF1_230( .Z(N1043), .A(N589) );
  BUF_X1 BUFF1_231( .Z(N1046), .A(N598) );
  BUF_X1 BUFF1_232( .Z(N1049), .A(N598) );
  NAND2_X1 NAND2_233( .ZN(N1054), .A1(N619), .A2(N888) );
  NAND2_X1 NAND2_234( .ZN(N1055), .A1(N616), .A2(N889) );
  NAND2_X1 NAND2_235( .ZN(N1063), .A1(N625), .A2(N890) );
  NAND2_X1 NAND2_236( .ZN(N1064), .A1(N622), .A2(N891) );
  NAND2_X1 NAND2_237( .ZN(N1067), .A1(N655), .A2(N895) );
  NAND2_X1 NAND2_238( .ZN(N1068), .A1(N652), .A2(N896) );
  NAND2_X1 NAND2_239( .ZN(N1119), .A1(N721), .A2(N988) );
  NAND2_X1 NAND2_240( .ZN(N1120), .A1(N718), .A2(N989) );
  NAND2_X1 NAND2_241( .ZN(N1121), .A1(N727), .A2(N991) );
  NAND2_X1 NAND2_242( .ZN(N1122), .A1(N724), .A2(N992) );
  NAND2_X1 NAND2_243( .ZN(N1128), .A1(N739), .A2(N1002) );
  NAND2_X1 NAND2_244( .ZN(N1129), .A1(N736), .A2(N1003) );
  NAND2_X1 NAND2_245( .ZN(N1130), .A1(N745), .A2(N1005) );
  NAND2_X1 NAND2_246( .ZN(N1131), .A1(N742), .A2(N1006) );
  NAND2_X1 NAND2_247( .ZN(N1132), .A1(N751), .A2(N1008) );
  NAND2_X1 NAND2_248( .ZN(N1133), .A1(N748), .A2(N1009) );
  INV_X1 NOT1_249( .ZN(N1148), .A(N939) );
  INV_X1 NOT1_250( .ZN(N1149), .A(N935) );
  NAND2_X2 NAND2_251( .ZN(N1150), .A1(N1054), .A2(N1055) );
  INV_X1 NOT1_252( .ZN(N1151), .A(N943) );
  INV_X1 NOT1_253( .ZN(N1152), .A(N947) );
  INV_X1 NOT1_254( .ZN(N1153), .A(N955) );
  INV_X1 NOT1_255( .ZN(N1154), .A(N951) );
  INV_X1 NOT1_256( .ZN(N1155), .A(N962) );
  INV_X1 NOT1_257( .ZN(N1156), .A(N969) );
  INV_X1 NOT1_258( .ZN(N1157), .A(N977) );
  NAND2_X1 NAND2_259( .ZN(N1158), .A1(N1063), .A2(N1064) );
  INV_X1 NOT1_260( .ZN(N1159), .A(N985) );
  NAND2_X1 NAND2_261( .ZN(N1160), .A1(N985), .A2(N892) );
  INV_X1 NOT1_262( .ZN(N1161), .A(N998) );
  NAND2_X1 NAND2_263( .ZN(N1162), .A1(N1067), .A2(N1068) );
  INV_X2 NOT1_264( .ZN(N1163), .A(N899) );
  BUF_X1 BUFF1_265( .Z(N1164), .A(N899) );
  INV_X1 NOT1_266( .ZN(N1167), .A(N903) );
  BUF_X1 BUFF1_267( .Z(N1168), .A(N903) );
  NAND2_X1 NAND2_268( .ZN(N1171), .A1(N921), .A2(N923) );
  NAND2_X1 NAND2_269( .ZN(N1188), .A1(N922), .A2(N923) );
  INV_X1 NOT1_270( .ZN(N1205), .A(N1010) );
  NAND2_X1 NAND2_271( .ZN(N1206), .A1(N1010), .A2(N938) );
  INV_X1 NOT1_272( .ZN(N1207), .A(N1013) );
  NAND2_X1 NAND2_273( .ZN(N1208), .A1(N1013), .A2(N942) );
  INV_X1 NOT1_274( .ZN(N1209), .A(N1016) );
  NAND2_X1 NAND2_275( .ZN(N1210), .A1(N1016), .A2(N946) );
  INV_X1 NOT1_276( .ZN(N1211), .A(N1019) );
  NAND2_X1 NAND2_277( .ZN(N1212), .A1(N1019), .A2(N950) );
  INV_X1 NOT1_278( .ZN(N1213), .A(N1022) );
  NAND2_X1 NAND2_279( .ZN(N1214), .A1(N1022), .A2(N954) );
  INV_X1 NOT1_280( .ZN(N1215), .A(N1025) );
  NAND2_X1 NAND2_281( .ZN(N1216), .A1(N1025), .A2(N958) );
  INV_X1 NOT1_282( .ZN(N1217), .A(N1028) );
  INV_X1 NOT1_283( .ZN(N1218), .A(N959) );
  INV_X1 NOT1_284( .ZN(N1219), .A(N1031) );
  INV_X1 NOT1_285( .ZN(N1220), .A(N1034) );
  NAND2_X1 NAND2_286( .ZN(N1221), .A1(N1034), .A2(N968) );
  INV_X1 NOT1_287( .ZN(N1222), .A(N965) );
  INV_X1 NOT1_288( .ZN(N1223), .A(N1037) );
  NAND2_X1 NAND2_289( .ZN(N1224), .A1(N1037), .A2(N972) );
  INV_X1 NOT1_290( .ZN(N1225), .A(N1040) );
  NAND2_X1 NAND2_291( .ZN(N1226), .A1(N1040), .A2(N976) );
  INV_X1 NOT1_292( .ZN(N1227), .A(N973) );
  INV_X1 NOT1_293( .ZN(N1228), .A(N1043) );
  NAND2_X1 NAND2_294( .ZN(N1229), .A1(N1043), .A2(N980) );
  INV_X1 NOT1_295( .ZN(N1230), .A(N981) );
  NAND2_X1 NAND2_296( .ZN(N1231), .A1(N981), .A2(N984) );
  NAND2_X1 NAND2_297( .ZN(N1232), .A1(N1119), .A2(N1120) );
  NAND2_X1 NAND2_298( .ZN(N1235), .A1(N1121), .A2(N1122) );
  INV_X1 NOT1_299( .ZN(N1238), .A(N1046) );
  NAND2_X1 NAND2_300( .ZN(N1239), .A1(N1046), .A2(N997) );
  INV_X1 NOT1_301( .ZN(N1240), .A(N994) );
  INV_X1 NOT1_302( .ZN(N1241), .A(N1049) );
  NAND2_X1 NAND2_303( .ZN(N1242), .A1(N1049), .A2(N1001) );
  NAND2_X1 NAND2_304( .ZN(N1243), .A1(N1128), .A2(N1129) );
  NAND2_X1 NAND2_305( .ZN(N1246), .A1(N1130), .A2(N1131) );
  NAND2_X1 NAND2_306( .ZN(N1249), .A1(N1132), .A2(N1133) );
  BUF_X1 BUFF1_307( .Z(N1252), .A(N907) );
  BUF_X1 BUFF1_308( .Z(N1255), .A(N907) );
  BUF_X1 BUFF1_309( .Z(N1258), .A(N910) );
  BUF_X1 BUFF1_310( .Z(N1261), .A(N910) );
  INV_X8 NOT1_311( .ZN(N1264), .A(N1150) );
  NAND2_X1 NAND2_312( .ZN(N1267), .A1(N631), .A2(N1159) );
  NAND2_X1 NAND2_313( .ZN(N1309), .A1(N688), .A2(N1205) );
  NAND2_X1 NAND2_314( .ZN(N1310), .A1(N691), .A2(N1207) );
  NAND2_X1 NAND2_315( .ZN(N1311), .A1(N694), .A2(N1209) );
  NAND2_X1 NAND2_316( .ZN(N1312), .A1(N697), .A2(N1211) );
  NAND2_X1 NAND2_317( .ZN(N1313), .A1(N700), .A2(N1213) );
  NAND2_X1 NAND2_318( .ZN(N1314), .A1(N703), .A2(N1215) );
  NAND2_X1 NAND2_319( .ZN(N1315), .A1(N706), .A2(N1220) );
  NAND2_X1 NAND2_320( .ZN(N1316), .A1(N709), .A2(N1223) );
  NAND2_X1 NAND2_321( .ZN(N1317), .A1(N712), .A2(N1225) );
  NAND2_X1 NAND2_322( .ZN(N1318), .A1(N715), .A2(N1228) );
  INV_X8 NOT1_323( .ZN(N1319), .A(N1158) );
  NAND2_X1 NAND2_324( .ZN(N1322), .A1(N628), .A2(N1230) );
  NAND2_X1 NAND2_325( .ZN(N1327), .A1(N730), .A2(N1238) );
  NAND2_X1 NAND2_326( .ZN(N1328), .A1(N733), .A2(N1241) );
  INV_X8 NOT1_327( .ZN(N1334), .A(N1162) );
  NAND2_X1 NAND2_328( .ZN(N1344), .A1(N1267), .A2(N1160) );
  NAND2_X1 NAND2_329( .ZN(N1345), .A1(N1249), .A2(N894) );
  INV_X8 NOT1_330( .ZN(N1346), .A(N1249) );
  INV_X1 NOT1_331( .ZN(N1348), .A(N1255) );
  INV_X1 NOT1_332( .ZN(N1349), .A(N1252) );
  INV_X1 NOT1_333( .ZN(N1350), .A(N1261) );
  INV_X1 NOT1_334( .ZN(N1351), .A(N1258) );
  NAND2_X1 NAND2_335( .ZN(N1352), .A1(N1309), .A2(N1206) );
  NAND2_X1 NAND2_336( .ZN(N1355), .A1(N1310), .A2(N1208) );
  NAND2_X1 NAND2_337( .ZN(N1358), .A1(N1311), .A2(N1210) );
  NAND2_X1 NAND2_338( .ZN(N1361), .A1(N1312), .A2(N1212) );
  NAND2_X1 NAND2_339( .ZN(N1364), .A1(N1313), .A2(N1214) );
  NAND2_X1 NAND2_340( .ZN(N1367), .A1(N1314), .A2(N1216) );
  NAND2_X1 NAND2_341( .ZN(N1370), .A1(N1315), .A2(N1221) );
  NAND2_X1 NAND2_342( .ZN(N1373), .A1(N1316), .A2(N1224) );
  NAND2_X1 NAND2_343( .ZN(N1376), .A1(N1317), .A2(N1226) );
  NAND2_X1 NAND2_344( .ZN(N1379), .A1(N1318), .A2(N1229) );
  NAND2_X1 NAND2_345( .ZN(N1383), .A1(N1322), .A2(N1231) );
  INV_X1 NOT1_346( .ZN(N1386), .A(N1232) );
  NAND2_X1 NAND2_347( .ZN(N1387), .A1(N1232), .A2(N990) );
  INV_X1 NOT1_348( .ZN(N1388), .A(N1235) );
  NAND2_X2 NAND2_349( .ZN(N1389), .A1(N1235), .A2(N993) );
  NAND2_X2 NAND2_350( .ZN(N1390), .A1(N1327), .A2(N1239) );
  NAND2_X1 NAND2_351( .ZN(N1393), .A1(N1328), .A2(N1242) );
  INV_X1 NOT1_352( .ZN(N1396), .A(N1243) );
  NAND2_X1 NAND2_353( .ZN(N1397), .A1(N1243), .A2(N1004) );
  INV_X1 NOT1_354( .ZN(N1398), .A(N1246) );
  NAND2_X1 NAND2_355( .ZN(N1399), .A1(N1246), .A2(N1007) );
  INV_X1 NOT1_356( .ZN(N1409), .A(N1319) );
  NAND2_X1 NAND2_357( .ZN(N1412), .A1(N649), .A2(N1346) );
  INV_X1 NOT1_358( .ZN(N1413), .A(N1334) );
  BUF_X2 BUFF1_359( .Z(N1416), .A(N1264) );
  BUF_X2 BUFF1_360( .Z(N1419), .A(N1264) );
  NAND2_X1 NAND2_361( .ZN(N1433), .A1(N634), .A2(N1386) );
  NAND2_X1 NAND2_362( .ZN(N1434), .A1(N637), .A2(N1388) );
  NAND2_X1 NAND2_363( .ZN(N1438), .A1(N640), .A2(N1396) );
  NAND2_X1 NAND2_364( .ZN(N1439), .A1(N646), .A2(N1398) );
  INV_X1 NOT1_365( .ZN(N1440), .A(N1344) );
  NAND2_X1 NAND2_366( .ZN(N1443), .A1(N1355), .A2(N1148) );
  INV_X1 NOT1_367( .ZN(N1444), .A(N1355) );
  NAND2_X1 NAND2_368( .ZN(N1445), .A1(N1352), .A2(N1149) );
  INV_X1 NOT1_369( .ZN(N1446), .A(N1352) );
  NAND2_X1 NAND2_370( .ZN(N1447), .A1(N1358), .A2(N1151) );
  INV_X1 NOT1_371( .ZN(N1448), .A(N1358) );
  NAND2_X1 NAND2_372( .ZN(N1451), .A1(N1361), .A2(N1152) );
  INV_X1 NOT1_373( .ZN(N1452), .A(N1361) );
  NAND2_X1 NAND2_374( .ZN(N1453), .A1(N1367), .A2(N1153) );
  INV_X1 NOT1_375( .ZN(N1454), .A(N1367) );
  NAND2_X1 NAND2_376( .ZN(N1455), .A1(N1364), .A2(N1154) );
  INV_X1 NOT1_377( .ZN(N1456), .A(N1364) );
  NAND2_X1 NAND2_378( .ZN(N1457), .A1(N1373), .A2(N1156) );
  INV_X1 NOT1_379( .ZN(N1458), .A(N1373) );
  NAND2_X1 NAND2_380( .ZN(N1459), .A1(N1379), .A2(N1157) );
  INV_X1 NOT1_381( .ZN(N1460), .A(N1379) );
  INV_X1 NOT1_382( .ZN(N1461), .A(N1383) );
  NAND2_X1 NAND2_383( .ZN(N1462), .A1(N1393), .A2(N1161) );
  INV_X1 NOT1_384( .ZN(N1463), .A(N1393) );
  NAND2_X1 NAND2_385( .ZN(N1464), .A1(N1345), .A2(N1412) );
  INV_X1 NOT1_386( .ZN(N1468), .A(N1370) );
  NAND2_X1 NAND2_387( .ZN(N1469), .A1(N1370), .A2(N1222) );
  INV_X1 NOT1_388( .ZN(N1470), .A(N1376) );
  NAND2_X1 NAND2_389( .ZN(N1471), .A1(N1376), .A2(N1227) );
  NAND2_X1 NAND2_390( .ZN(N1472), .A1(N1387), .A2(N1433) );
  INV_X1 NOT1_391( .ZN(N1475), .A(N1390) );
  NAND2_X1 NAND2_392( .ZN(N1476), .A1(N1390), .A2(N1240) );
  NAND2_X1 NAND2_393( .ZN(N1478), .A1(N1389), .A2(N1434) );
  NAND2_X1 NAND2_394( .ZN(N1481), .A1(N1399), .A2(N1439) );
  NAND2_X1 NAND2_395( .ZN(N1484), .A1(N1397), .A2(N1438) );
  NAND2_X1 NAND2_396( .ZN(N1487), .A1(N939), .A2(N1444) );
  NAND2_X1 NAND2_397( .ZN(N1488), .A1(N935), .A2(N1446) );
  NAND2_X1 NAND2_398( .ZN(N1489), .A1(N943), .A2(N1448) );
  INV_X1 NOT1_399( .ZN(N1490), .A(N1419) );
  INV_X1 NOT1_400( .ZN(N1491), .A(N1416) );
  NAND2_X1 NAND2_401( .ZN(N1492), .A1(N947), .A2(N1452) );
  NAND2_X1 NAND2_402( .ZN(N1493), .A1(N955), .A2(N1454) );
  NAND2_X1 NAND2_403( .ZN(N1494), .A1(N951), .A2(N1456) );
  NAND2_X1 NAND2_404( .ZN(N1495), .A1(N969), .A2(N1458) );
  NAND2_X1 NAND2_405( .ZN(N1496), .A1(N977), .A2(N1460) );
  NAND2_X1 NAND2_406( .ZN(N1498), .A1(N998), .A2(N1463) );
  INV_X1 NOT1_407( .ZN(N1499), .A(N1440) );
  NAND2_X1 NAND2_408( .ZN(N1500), .A1(N965), .A2(N1468) );
  NAND2_X1 NAND2_409( .ZN(N1501), .A1(N973), .A2(N1470) );
  NAND2_X1 NAND2_410( .ZN(N1504), .A1(N994), .A2(N1475) );
  INV_X1 NOT1_411( .ZN(N1510), .A(N1464) );
  NAND2_X1 NAND2_412( .ZN(N1513), .A1(N1443), .A2(N1487) );
  NAND2_X1 NAND2_413( .ZN(N1514), .A1(N1445), .A2(N1488) );
  NAND2_X1 NAND2_414( .ZN(N1517), .A1(N1447), .A2(N1489) );
  NAND2_X1 NAND2_415( .ZN(N1520), .A1(N1451), .A2(N1492) );
  NAND2_X1 NAND2_416( .ZN(N1521), .A1(N1453), .A2(N1493) );
  NAND2_X1 NAND2_417( .ZN(N1522), .A1(N1455), .A2(N1494) );
  NAND2_X1 NAND2_418( .ZN(N1526), .A1(N1457), .A2(N1495) );
  NAND2_X1 NAND2_419( .ZN(N1527), .A1(N1459), .A2(N1496) );
  INV_X8 NOT1_420( .ZN(N1528), .A(N1472) );
  NAND2_X1 NAND2_421( .ZN(N1529), .A1(N1462), .A2(N1498) );
  INV_X8 NOT1_422( .ZN(N1530), .A(N1478) );
  INV_X8 NOT1_423( .ZN(N1531), .A(N1481) );
  INV_X1 NOT1_424( .ZN(N1532), .A(N1484) );
  NAND2_X1 NAND2_425( .ZN(N1534), .A1(N1471), .A2(N1501) );
  NAND2_X1 NAND2_426( .ZN(N1537), .A1(N1469), .A2(N1500) );
  NAND2_X1 NAND2_427( .ZN(N1540), .A1(N1476), .A2(N1504) );
  INV_X1 NOT1_428( .ZN(N1546), .A(N1513) );
  INV_X1 NOT1_429( .ZN(N1554), .A(N1521) );
  INV_X1 NOT1_430( .ZN(N1557), .A(N1526) );
  INV_X1 NOT1_431( .ZN(N1561), .A(N1520) );
  NAND2_X1 NAND2_432( .ZN(N1567), .A1(N1484), .A2(N1531) );
  NAND2_X1 NAND2_433( .ZN(N1568), .A1(N1481), .A2(N1532) );
  INV_X1 NOT1_434( .ZN(N1569), .A(N1510) );
  INV_X1 NOT1_435( .ZN(N1571), .A(N1527) );
  INV_X1 NOT1_436( .ZN(N1576), .A(N1529) );
  BUF_X4 BUFF1_437( .Z(N1588), .A(N1522) );
  INV_X1 NOT1_438( .ZN(N1591), .A(N1534) );
  INV_X1 NOT1_439( .ZN(N1593), .A(N1537) );
  NAND2_X1 NAND2_440( .ZN(N1594), .A1(N1540), .A2(N1530) );
  INV_X1 NOT1_441( .ZN(N1595), .A(N1540) );
  NAND2_X1 NAND2_442( .ZN(N1596), .A1(N1567), .A2(N1568) );
  BUF_X1 BUFF1_443( .Z(N1600), .A(N1517) );
  BUF_X1 BUFF1_444( .Z(N1603), .A(N1517) );
  BUF_X1 BUFF1_445( .Z(N1606), .A(N1522) );
  BUF_X1 BUFF1_446( .Z(N1609), .A(N1522) );
  BUF_X1 BUFF1_447( .Z(N1612), .A(N1514) );
  BUF_X1 BUFF1_448( .Z(N1615), .A(N1514) );
  BUF_X1 BUFF1_449( .Z(N1620), .A(N1557) );
  BUF_X1 BUFF1_450( .Z(N1623), .A(N1554) );
  INV_X1 NOT1_451( .ZN(N1635), .A(N1571) );
  NAND2_X1 NAND2_452( .ZN(N1636), .A1(N1478), .A2(N1595) );
  NAND2_X1 NAND2_453( .ZN(N1638), .A1(N1576), .A2(N1569) );
  INV_X1 NOT1_454( .ZN(N1639), .A(N1576) );
  BUF_X1 BUFF1_455( .Z(N1640), .A(N1561) );
  BUF_X1 BUFF1_456( .Z(N1643), .A(N1561) );
  BUF_X1 BUFF1_457( .Z(N1647), .A(N1546) );
  BUF_X1 BUFF1_458( .Z(N1651), .A(N1546) );
  BUF_X1 BUFF1_459( .Z(N1658), .A(N1554) );
  BUF_X1 BUFF1_460( .Z(N1661), .A(N1557) );
  BUF_X1 BUFF1_461( .Z(N1664), .A(N1557) );
  NAND2_X1 NAND2_462( .ZN(N1671), .A1(N1596), .A2(N893) );
  INV_X1 NOT1_463( .ZN(N1672), .A(N1596) );
  INV_X1 NOT1_464( .ZN(N1675), .A(N1600) );
  INV_X1 NOT1_465( .ZN(N1677), .A(N1603) );
  NAND2_X1 NAND2_466( .ZN(N1678), .A1(N1606), .A2(N1217) );
  INV_X1 NOT1_467( .ZN(N1679), .A(N1606) );
  NAND2_X1 NAND2_468( .ZN(N1680), .A1(N1609), .A2(N1219) );
  INV_X1 NOT1_469( .ZN(N1681), .A(N1609) );
  INV_X1 NOT1_470( .ZN(N1682), .A(N1612) );
  INV_X1 NOT1_471( .ZN(N1683), .A(N1615) );
  NAND2_X1 NAND2_472( .ZN(N1685), .A1(N1594), .A2(N1636) );
  NAND2_X1 NAND2_473( .ZN(N1688), .A1(N1510), .A2(N1639) );
  BUF_X1 BUFF1_474( .Z(N1697), .A(N1588) );
  BUF_X1 BUFF1_475( .Z(N1701), .A(N1588) );
  NAND2_X1 NAND2_476( .ZN(N1706), .A1(N643), .A2(N1672) );
  INV_X1 NOT1_477( .ZN(N1707), .A(N1643) );
  NAND2_X1 NAND2_478( .ZN(N1708), .A1(N1647), .A2(N1675) );
  INV_X1 NOT1_479( .ZN(N1709), .A(N1647) );
  NAND2_X1 NAND2_480( .ZN(N1710), .A1(N1651), .A2(N1677) );
  INV_X1 NOT1_481( .ZN(N1711), .A(N1651) );
  NAND2_X1 NAND2_482( .ZN(N1712), .A1(N1028), .A2(N1679) );
  NAND2_X1 NAND2_483( .ZN(N1713), .A1(N1031), .A2(N1681) );
  BUF_X1 BUFF1_484( .Z(N1714), .A(N1620) );
  BUF_X1 BUFF1_485( .Z(N1717), .A(N1620) );
  NAND2_X1 NAND2_486( .ZN(N1720), .A1(N1658), .A2(N1593) );
  INV_X1 NOT1_487( .ZN(N1721), .A(N1658) );
  NAND2_X1 NAND2_488( .ZN(N1723), .A1(N1638), .A2(N1688) );
  INV_X1 NOT1_489( .ZN(N1727), .A(N1661) );
  INV_X1 NOT1_490( .ZN(N1728), .A(N1640) );
  INV_X1 NOT1_491( .ZN(N1730), .A(N1664) );
  BUF_X1 BUFF1_492( .Z(N1731), .A(N1623) );
  BUF_X1 BUFF1_493( .Z(N1734), .A(N1623) );
  NAND2_X1 NAND2_494( .ZN(N1740), .A1(N1685), .A2(N1528) );
  INV_X1 NOT1_495( .ZN(N1741), .A(N1685) );
  NAND2_X1 NAND2_496( .ZN(N1742), .A1(N1671), .A2(N1706) );
  NAND2_X1 NAND2_497( .ZN(N1746), .A1(N1600), .A2(N1709) );
  NAND2_X1 NAND2_498( .ZN(N1747), .A1(N1603), .A2(N1711) );
  NAND2_X1 NAND2_499( .ZN(N1748), .A1(N1678), .A2(N1712) );
  NAND2_X1 NAND2_500( .ZN(N1751), .A1(N1680), .A2(N1713) );
  NAND2_X1 NAND2_501( .ZN(N1759), .A1(N1537), .A2(N1721) );
  INV_X1 NOT1_502( .ZN(N1761), .A(N1697) );
  NAND2_X1 NAND2_503( .ZN(N1762), .A1(N1697), .A2(N1727) );
  INV_X1 NOT1_504( .ZN(N1763), .A(N1701) );
  NAND2_X1 NAND2_505( .ZN(N1764), .A1(N1701), .A2(N1730) );
  INV_X1 NOT1_506( .ZN(N1768), .A(N1717) );
  NAND2_X1 NAND2_507( .ZN(N1769), .A1(N1472), .A2(N1741) );
  NAND2_X1 NAND2_508( .ZN(N1772), .A1(N1723), .A2(N1413) );
  INV_X4 NOT1_509( .ZN(N1773), .A(N1723) );
  NAND2_X1 NAND2_510( .ZN(N1774), .A1(N1708), .A2(N1746) );
  NAND2_X1 NAND2_511( .ZN(N1777), .A1(N1710), .A2(N1747) );
  INV_X4 NOT1_512( .ZN(N1783), .A(N1731) );
  NAND2_X1 NAND2_513( .ZN(N1784), .A1(N1731), .A2(N1682) );
  INV_X1 NOT1_514( .ZN(N1785), .A(N1714) );
  INV_X1 NOT1_515( .ZN(N1786), .A(N1734) );
  NAND2_X1 NAND2_516( .ZN(N1787), .A1(N1734), .A2(N1683) );
  NAND2_X1 NAND2_517( .ZN(N1788), .A1(N1720), .A2(N1759) );
  NAND2_X1 NAND2_518( .ZN(N1791), .A1(N1661), .A2(N1761) );
  NAND2_X1 NAND2_519( .ZN(N1792), .A1(N1664), .A2(N1763) );
  NAND2_X1 NAND2_520( .ZN(N1795), .A1(N1751), .A2(N1155) );
  INV_X1 NOT1_521( .ZN(N1796), .A(N1751) );
  NAND2_X1 NAND2_522( .ZN(N1798), .A1(N1740), .A2(N1769) );
  NAND2_X1 NAND2_523( .ZN(N1801), .A1(N1334), .A2(N1773) );
  NAND2_X1 NAND2_524( .ZN(N1802), .A1(N1742), .A2(N290) );
  INV_X1 NOT1_525( .ZN(N1807), .A(N1748) );
  NAND2_X1 NAND2_526( .ZN(N1808), .A1(N1748), .A2(N1218) );
  NAND2_X1 NAND2_527( .ZN(N1809), .A1(N1612), .A2(N1783) );
  NAND2_X1 NAND2_528( .ZN(N1810), .A1(N1615), .A2(N1786) );
  NAND2_X1 NAND2_529( .ZN(N1812), .A1(N1791), .A2(N1762) );
  NAND2_X1 NAND2_530( .ZN(N1815), .A1(N1792), .A2(N1764) );
  BUF_X1 BUFF1_531( .Z(N1818), .A(N1742) );
  NAND2_X1 NAND2_532( .ZN(N1821), .A1(N1777), .A2(N1490) );
  INV_X1 NOT1_533( .ZN(N1822), .A(N1777) );
  NAND2_X1 NAND2_534( .ZN(N1823), .A1(N1774), .A2(N1491) );
  INV_X1 NOT1_535( .ZN(N1824), .A(N1774) );
  NAND2_X1 NAND2_536( .ZN(N1825), .A1(N962), .A2(N1796) );
  NAND2_X1 NAND2_537( .ZN(N1826), .A1(N1788), .A2(N1409) );
  INV_X1 NOT1_538( .ZN(N1827), .A(N1788) );
  NAND2_X1 NAND2_539( .ZN(N1830), .A1(N1772), .A2(N1801) );
  NAND2_X1 NAND2_540( .ZN(N1837), .A1(N959), .A2(N1807) );
  NAND2_X1 NAND2_541( .ZN(N1838), .A1(N1809), .A2(N1784) );
  NAND2_X1 NAND2_542( .ZN(N1841), .A1(N1810), .A2(N1787) );
  NAND2_X2 NAND2_543( .ZN(N1848), .A1(N1419), .A2(N1822) );
  NAND2_X2 NAND2_544( .ZN(N1849), .A1(N1416), .A2(N1824) );
  NAND2_X2 NAND2_545( .ZN(N1850), .A1(N1795), .A2(N1825) );
  NAND2_X1 NAND2_546( .ZN(N1852), .A1(N1319), .A2(N1827) );
  NAND2_X1 NAND2_547( .ZN(N1855), .A1(N1815), .A2(N1707) );
  INV_X1 NOT1_548( .ZN(N1856), .A(N1815) );
  INV_X1 NOT1_549( .ZN(N1857), .A(N1818) );
  NAND2_X1 NAND2_550( .ZN(N1858), .A1(N1798), .A2(N290) );
  INV_X1 NOT1_551( .ZN(N1864), .A(N1812) );
  NAND2_X1 NAND2_552( .ZN(N1865), .A1(N1812), .A2(N1728) );
  BUF_X1 BUFF1_553( .Z(N1866), .A(N1798) );
  BUF_X1 BUFF1_554( .Z(N1869), .A(N1802) );
  BUF_X1 BUFF1_555( .Z(N1872), .A(N1802) );
  NAND2_X1 NAND2_556( .ZN(N1875), .A1(N1808), .A2(N1837) );
  NAND2_X1 NAND2_557( .ZN(N1878), .A1(N1821), .A2(N1848) );
  NAND2_X1 NAND2_558( .ZN(N1879), .A1(N1823), .A2(N1849) );
  NAND2_X1 NAND2_559( .ZN(N1882), .A1(N1841), .A2(N1768) );
  INV_X1 NOT1_560( .ZN(N1883), .A(N1841) );
  NAND2_X1 NAND2_561( .ZN(N1884), .A1(N1826), .A2(N1852) );
  NAND2_X1 NAND2_562( .ZN(N1885), .A1(N1643), .A2(N1856) );
  NAND2_X1 NAND2_563( .ZN(N1889), .A1(N1830), .A2(N290) );
  INV_X1 NOT1_564( .ZN(N1895), .A(N1838) );
  NAND2_X1 NAND2_565( .ZN(N1896), .A1(N1838), .A2(N1785) );
  NAND2_X1 NAND2_566( .ZN(N1897), .A1(N1640), .A2(N1864) );
  INV_X1 NOT1_567( .ZN(N1898), .A(N1850) );
  BUF_X1 BUFF1_568( .Z(N1902), .A(N1830) );
  INV_X1 NOT1_569( .ZN(N1910), .A(N1878) );
  NAND2_X1 NAND2_570( .ZN(N1911), .A1(N1717), .A2(N1883) );
  INV_X1 NOT1_571( .ZN(N1912), .A(N1884) );
  NAND2_X1 NAND2_572( .ZN(N1913), .A1(N1855), .A2(N1885) );
  INV_X1 NOT1_573( .ZN(N1915), .A(N1866) );
  NAND2_X1 NAND2_574( .ZN(N1919), .A1(N1872), .A2(N919) );
  INV_X1 NOT1_575( .ZN(N1920), .A(N1872) );
  NAND2_X1 NAND2_576( .ZN(N1921), .A1(N1869), .A2(N920) );
  INV_X1 NOT1_577( .ZN(N1922), .A(N1869) );
  INV_X1 NOT1_578( .ZN(N1923), .A(N1875) );
  NAND2_X1 NAND2_579( .ZN(N1924), .A1(N1714), .A2(N1895) );
  BUF_X4 BUFF1_580( .Z(N1927), .A(N1858) );
  BUF_X4 BUFF1_581( .Z(N1930), .A(N1858) );
  NAND2_X1 NAND2_582( .ZN(N1933), .A1(N1865), .A2(N1897) );
  NAND2_X1 NAND2_583( .ZN(N1936), .A1(N1882), .A2(N1911) );
  INV_X1 NOT1_584( .ZN(N1937), .A(N1898) );
  INV_X1 NOT1_585( .ZN(N1938), .A(N1902) );
  NAND2_X1 NAND2_586( .ZN(N1941), .A1(N679), .A2(N1920) );
  NAND2_X1 NAND2_587( .ZN(N1942), .A1(N676), .A2(N1922) );
  BUF_X1 BUFF1_588( .Z(N1944), .A(N1879) );
  INV_X1 NOT1_589( .ZN(N1947), .A(N1913) );
  BUF_X1 BUFF1_590( .Z(N1950), .A(N1889) );
  BUF_X1 BUFF1_591( .Z(N1953), .A(N1889) );
  BUF_X1 BUFF1_592( .Z(N1958), .A(N1879) );
  NAND2_X1 NAND2_593( .ZN(N1961), .A1(N1896), .A2(N1924) );
  AND2_X1 AND2_594( .ZN(N1965), .A1(N1910), .A2(N601) );
  AND2_X1 AND2_595( .ZN(N1968), .A1(N602), .A2(N1912) );
  NAND2_X1 NAND2_596( .ZN(N1975), .A1(N1930), .A2(N917) );
  INV_X1 NOT1_597( .ZN(N1976), .A(N1930) );
  NAND2_X1 NAND2_598( .ZN(N1977), .A1(N1927), .A2(N918) );
  INV_X1 NOT1_599( .ZN(N1978), .A(N1927) );
  NAND2_X1 NAND2_600( .ZN(N1979), .A1(N1919), .A2(N1941) );
  NAND2_X1 NAND2_601( .ZN(N1980), .A1(N1921), .A2(N1942) );
  INV_X1 NOT1_602( .ZN(N1985), .A(N1933) );
  INV_X1 NOT1_603( .ZN(N1987), .A(N1936) );
  INV_X1 NOT1_604( .ZN(N1999), .A(N1944) );
  NAND2_X1 NAND2_605( .ZN(N2000), .A1(N1944), .A2(N1937) );
  INV_X1 NOT1_606( .ZN(N2002), .A(N1947) );
  NAND2_X1 NAND2_607( .ZN(N2003), .A1(N1947), .A2(N1499) );
  NAND2_X1 NAND2_608( .ZN(N2004), .A1(N1953), .A2(N1350) );
  INV_X1 NOT1_609( .ZN(N2005), .A(N1953) );
  NAND2_X1 NAND2_610( .ZN(N2006), .A1(N1950), .A2(N1351) );
  INV_X1 NOT1_611( .ZN(N2007), .A(N1950) );
  NAND2_X1 NAND2_612( .ZN(N2008), .A1(N673), .A2(N1976) );
  NAND2_X1 NAND2_613( .ZN(N2009), .A1(N670), .A2(N1978) );
  INV_X1 NOT1_614( .ZN(N2012), .A(N1979) );
  INV_X1 NOT1_615( .ZN(N2013), .A(N1958) );
  NAND2_X1 NAND2_616( .ZN(N2014), .A1(N1958), .A2(N1923) );
  INV_X1 NOT1_617( .ZN(N2015), .A(N1961) );
  NAND2_X1 NAND2_618( .ZN(N2016), .A1(N1961), .A2(N1635) );
  INV_X1 NOT1_619( .ZN(N2018), .A(N1965) );
  INV_X1 NOT1_620( .ZN(N2019), .A(N1968) );
  NAND2_X1 NAND2_621( .ZN(N2020), .A1(N1898), .A2(N1999) );
  INV_X1 NOT1_622( .ZN(N2021), .A(N1987) );
  NAND2_X1 NAND2_623( .ZN(N2022), .A1(N1987), .A2(N1591) );
  NAND2_X1 NAND2_624( .ZN(N2023), .A1(N1440), .A2(N2002) );
  NAND2_X1 NAND2_625( .ZN(N2024), .A1(N1261), .A2(N2005) );
  NAND2_X1 NAND2_626( .ZN(N2025), .A1(N1258), .A2(N2007) );
  NAND2_X1 NAND2_627( .ZN(N2026), .A1(N1975), .A2(N2008) );
  NAND2_X1 NAND2_628( .ZN(N2027), .A1(N1977), .A2(N2009) );
  INV_X1 NOT1_629( .ZN(N2030), .A(N1980) );
  BUF_X1 BUFF1_630( .Z(N2033), .A(N1980) );
  NAND2_X1 NAND2_631( .ZN(N2036), .A1(N1875), .A2(N2013) );
  NAND2_X1 NAND2_632( .ZN(N2037), .A1(N1571), .A2(N2015) );
  NAND2_X1 NAND2_633( .ZN(N2038), .A1(N2020), .A2(N2000) );
  NAND2_X1 NAND2_634( .ZN(N2039), .A1(N1534), .A2(N2021) );
  NAND2_X1 NAND2_635( .ZN(N2040), .A1(N2023), .A2(N2003) );
  NAND2_X1 NAND2_636( .ZN(N2041), .A1(N2004), .A2(N2024) );
  NAND2_X1 NAND2_637( .ZN(N2042), .A1(N2006), .A2(N2025) );
  INV_X1 NOT1_638( .ZN(N2047), .A(N2026) );
  NAND2_X1 NAND2_639( .ZN(N2052), .A1(N2036), .A2(N2014) );
  NAND2_X1 NAND2_640( .ZN(N2055), .A1(N2037), .A2(N2016) );
  INV_X1 NOT1_641( .ZN(N2060), .A(N2038) );
  NAND2_X1 NAND2_642( .ZN(N2061), .A1(N2039), .A2(N2022) );
  NAND2_X1 NAND2_643( .ZN(N2062), .A1(N2040), .A2(N290) );
  INV_X1 NOT1_644( .ZN(N2067), .A(N2041) );
  INV_X1 NOT1_645( .ZN(N2068), .A(N2027) );
  BUF_X1 BUFF1_646( .Z(N2071), .A(N2027) );
  INV_X1 NOT1_647( .ZN(N2076), .A(N2052) );
  INV_X1 NOT1_648( .ZN(N2077), .A(N2055) );
  NAND2_X1 NAND2_649( .ZN(N2078), .A1(N2060), .A2(N290) );
  NAND2_X1 NAND2_650( .ZN(N2081), .A1(N2061), .A2(N290) );
  INV_X1 NOT1_651( .ZN(N2086), .A(N2042) );
  BUF_X1 BUFF1_652( .Z(N2089), .A(N2042) );
  AND2_X1 AND2_653( .ZN(N2104), .A1(N2030), .A2(N2068) );
  AND2_X1 AND2_654( .ZN(N2119), .A1(N2033), .A2(N2068) );
  AND2_X1 AND2_655( .ZN(N2129), .A1(N2030), .A2(N2071) );
  AND2_X1 AND2_656( .ZN(N2143), .A1(N2033), .A2(N2071) );
  BUF_X1 BUFF1_657( .Z(N2148), .A(N2062) );
  BUF_X1 BUFF1_658( .Z(N2151), .A(N2062) );
  BUF_X1 BUFF1_659( .Z(N2196), .A(N2078) );
  BUF_X1 BUFF1_660( .Z(N2199), .A(N2078) );
  BUF_X1 BUFF1_661( .Z(N2202), .A(N2081) );
  BUF_X1 BUFF1_662( .Z(N2205), .A(N2081) );
  NAND2_X1 NAND2_663( .ZN(N2214), .A1(N2151), .A2(N915) );
  INV_X1 NOT1_664( .ZN(N2215), .A(N2151) );
  NAND2_X1 NAND2_665( .ZN(N2216), .A1(N2148), .A2(N916) );
  INV_X1 NOT1_666( .ZN(N2217), .A(N2148) );
  NAND2_X1 NAND2_667( .ZN(N2222), .A1(N2199), .A2(N1348) );
  INV_X1 NOT1_668( .ZN(N2223), .A(N2199) );
  NAND2_X1 NAND2_669( .ZN(N2224), .A1(N2196), .A2(N1349) );
  INV_X1 NOT1_670( .ZN(N2225), .A(N2196) );
  NAND2_X1 NAND2_671( .ZN(N2226), .A1(N2205), .A2(N913) );
  INV_X1 NOT1_672( .ZN(N2227), .A(N2205) );
  NAND2_X1 NAND2_673( .ZN(N2228), .A1(N2202), .A2(N914) );
  INV_X1 NOT1_674( .ZN(N2229), .A(N2202) );
  NAND2_X1 NAND2_675( .ZN(N2230), .A1(N667), .A2(N2215) );
  NAND2_X1 NAND2_676( .ZN(N2231), .A1(N664), .A2(N2217) );
  NAND2_X1 NAND2_677( .ZN(N2232), .A1(N1255), .A2(N2223) );
  NAND2_X1 NAND2_678( .ZN(N2233), .A1(N1252), .A2(N2225) );
  NAND2_X1 NAND2_679( .ZN(N2234), .A1(N661), .A2(N2227) );
  NAND2_X1 NAND2_680( .ZN(N2235), .A1(N658), .A2(N2229) );
  NAND2_X1 NAND2_681( .ZN(N2236), .A1(N2214), .A2(N2230) );
  NAND2_X1 NAND2_682( .ZN(N2237), .A1(N2216), .A2(N2231) );
  NAND2_X1 NAND2_683( .ZN(N2240), .A1(N2222), .A2(N2232) );
  NAND2_X1 NAND2_684( .ZN(N2241), .A1(N2224), .A2(N2233) );
  NAND2_X1 NAND2_685( .ZN(N2244), .A1(N2226), .A2(N2234) );
  NAND2_X1 NAND2_686( .ZN(N2245), .A1(N2228), .A2(N2235) );
  INV_X1 NOT1_687( .ZN(N2250), .A(N2236) );
  INV_X1 NOT1_688( .ZN(N2253), .A(N2240) );
  INV_X1 NOT1_689( .ZN(N2256), .A(N2244) );
  INV_X1 NOT1_690( .ZN(N2257), .A(N2237) );
  BUF_X4 BUFF1_691( .Z(N2260), .A(N2237) );
  INV_X1 NOT1_692( .ZN(N2263), .A(N2241) );
  AND2_X1 AND2_693( .ZN(N2266), .A1(N1164), .A2(N2241) );
  INV_X1 NOT1_694( .ZN(N2269), .A(N2245) );
  AND2_X1 AND2_695( .ZN(N2272), .A1(N1168), .A2(N2245) );
  NAND4_X1 NAND8_696_A( .ZN(extra0), .A1(N2067), .A2(N2012), .A3(N2047), .A4(N2250) );
  NAND4_X1 NAND8_696_B( .ZN(extra1), .A1(extra0), .A2(N899), .A3(N2256), .A4(N2253) );
  NAND2_X1 NAND8_696( .ZN(N2279), .A1(extra1), .A2(N903) );
  BUF_X1 BUFF1_697( .Z(N2286), .A(N2266) );
  BUF_X1 BUFF1_698( .Z(N2297), .A(N2266) );
  BUF_X1 BUFF1_699( .Z(N2315), .A(N2272) );
  BUF_X1 BUFF1_700( .Z(N2326), .A(N2272) );
  AND2_X1 AND2_701( .ZN(N2340), .A1(N2086), .A2(N2257) );
  AND2_X1 AND2_702( .ZN(N2353), .A1(N2089), .A2(N2257) );
  AND2_X1 AND2_703( .ZN(N2361), .A1(N2086), .A2(N2260) );
  AND2_X1 AND2_704( .ZN(N2375), .A1(N2089), .A2(N2260) );
  AND4_X1 AND4_705( .ZN(N2384), .A1(N338), .A2(N2279), .A3(N313), .A4(N313) );
  AND2_X1 AND2_706( .ZN(N2385), .A1(N1163), .A2(N2263) );
  AND2_X1 AND2_707( .ZN(N2386), .A1(N1164), .A2(N2263) );
  AND2_X1 AND2_708( .ZN(N2426), .A1(N1167), .A2(N2269) );
  AND2_X1 AND2_709( .ZN(N2427), .A1(N1168), .A2(N2269) );
  NAND4_X1 NAND5_710_A( .ZN(extra2), .A1(N2286), .A2(N2315), .A3(N2361), .A4(N2104) );
  NAND2_X1 NAND5_710( .ZN(N2537), .A1(extra2), .A2(N1171) );
  NAND4_X1 NAND5_711_A( .ZN(extra3), .A1(N2286), .A2(N2315), .A3(N2340), .A4(N2129) );
  NAND2_X1 NAND5_711( .ZN(N2540), .A1(extra3), .A2(N1171) );
  NAND4_X1 NAND5_712_A( .ZN(extra4), .A1(N2286), .A2(N2315), .A3(N2340), .A4(N2119) );
  NAND2_X1 NAND5_712( .ZN(N2543), .A1(extra4), .A2(N1171) );
  NAND4_X1 NAND5_713_A( .ZN(extra5), .A1(N2286), .A2(N2315), .A3(N2353), .A4(N2104) );
  NAND2_X1 NAND5_713( .ZN(N2546), .A1(extra5), .A2(N1171) );
  NAND4_X1 NAND5_714_A( .ZN(extra6), .A1(N2297), .A2(N2315), .A3(N2375), .A4(N2119) );
  NAND2_X1 NAND5_714( .ZN(N2549), .A1(extra6), .A2(N1188) );
  NAND4_X1 NAND5_715_A( .ZN(extra7), .A1(N2297), .A2(N2326), .A3(N2361), .A4(N2143) );
  NAND2_X1 NAND5_715( .ZN(N2552), .A1(extra7), .A2(N1188) );
  NAND4_X1 NAND5_716_A( .ZN(extra8), .A1(N2297), .A2(N2326), .A3(N2375), .A4(N2129) );
  NAND2_X1 NAND5_716( .ZN(N2555), .A1(extra8), .A2(N1188) );
  AND4_X1 AND5_717_A( .ZN(extra9), .A1(N2286), .A2(N2315), .A3(N2361), .A4(N2104) );
  AND2_X1 AND5_717( .ZN(N2558), .A1(extra9), .A2(N1171) );
  AND4_X1 AND5_718_A( .ZN(extra10), .A1(N2286), .A2(N2315), .A3(N2340), .A4(N2129) );
  AND2_X1 AND5_718( .ZN(N2561), .A1(extra10), .A2(N1171) );
  AND4_X1 AND5_719_A( .ZN(extra11), .A1(N2286), .A2(N2315), .A3(N2340), .A4(N2119) );
  AND2_X1 AND5_719( .ZN(N2564), .A1(extra11), .A2(N1171) );
  AND4_X1 AND5_720_A( .ZN(extra12), .A1(N2286), .A2(N2315), .A3(N2353), .A4(N2104) );
  AND2_X1 AND5_720( .ZN(N2567), .A1(extra12), .A2(N1171) );
  AND4_X1 AND5_721_A( .ZN(extra13), .A1(N2297), .A2(N2315), .A3(N2375), .A4(N2119) );
  AND2_X1 AND5_721( .ZN(N2570), .A1(extra13), .A2(N1188) );
  AND4_X1 AND5_722_A( .ZN(extra14), .A1(N2297), .A2(N2326), .A3(N2361), .A4(N2143) );
  AND2_X1 AND5_722( .ZN(N2573), .A1(extra14), .A2(N1188) );
  AND4_X1 AND5_723_A( .ZN(extra15), .A1(N2297), .A2(N2326), .A3(N2375), .A4(N2129) );
  AND2_X1 AND5_723( .ZN(N2576), .A1(extra15), .A2(N1188) );
  NAND4_X1 NAND5_724_A( .ZN(extra16), .A1(N2286), .A2(N2427), .A3(N2361), .A4(N2129) );
  NAND2_X2 NAND5_724( .ZN(N2594), .A1(extra16), .A2(N1171) );
  NAND4_X1 NAND5_725_A( .ZN(extra17), .A1(N2297), .A2(N2427), .A3(N2361), .A4(N2119) );
  NAND2_X2 NAND5_725( .ZN(N2597), .A1(extra17), .A2(N1171) );
  NAND4_X1 NAND5_726_A( .ZN(extra18), .A1(N2297), .A2(N2427), .A3(N2375), .A4(N2104) );
  NAND2_X2 NAND5_726( .ZN(N2600), .A1(extra18), .A2(N1171) );
  NAND4_X1 NAND5_727_A( .ZN(extra19), .A1(N2297), .A2(N2427), .A3(N2340), .A4(N2143) );
  NAND2_X2 NAND5_727( .ZN(N2603), .A1(extra19), .A2(N1171) );
  NAND4_X1 NAND5_728_A( .ZN(extra20), .A1(N2297), .A2(N2427), .A3(N2353), .A4(N2129) );
  NAND2_X2 NAND5_728( .ZN(N2606), .A1(extra20), .A2(N1188) );
  NAND4_X1 NAND5_729_A( .ZN(extra21), .A1(N2386), .A2(N2326), .A3(N2361), .A4(N2129) );
  NAND2_X1 NAND5_729( .ZN(N2611), .A1(extra21), .A2(N1188) );
  NAND4_X1 NAND5_730_A( .ZN(extra22), .A1(N2386), .A2(N2326), .A3(N2361), .A4(N2119) );
  NAND2_X1 NAND5_730( .ZN(N2614), .A1(extra22), .A2(N1188) );
  NAND4_X1 NAND5_731_A( .ZN(extra23), .A1(N2386), .A2(N2326), .A3(N2375), .A4(N2104) );
  NAND2_X1 NAND5_731( .ZN(N2617), .A1(extra23), .A2(N1188) );
  NAND4_X1 NAND5_732_A( .ZN(extra24), .A1(N2386), .A2(N2326), .A3(N2353), .A4(N2129) );
  NAND2_X1 NAND5_732( .ZN(N2620), .A1(extra24), .A2(N1188) );
  NAND4_X1 NAND5_733_A( .ZN(extra25), .A1(N2297), .A2(N2427), .A3(N2340), .A4(N2104) );
  NAND2_X1 NAND5_733( .ZN(N2627), .A1(extra25), .A2(N926) );
  NAND4_X1 NAND5_734_A( .ZN(extra26), .A1(N2386), .A2(N2326), .A3(N2340), .A4(N2104) );
  NAND2_X1 NAND5_734( .ZN(N2628), .A1(extra26), .A2(N926) );
  NAND4_X1 NAND5_735_A( .ZN(extra27), .A1(N2386), .A2(N2427), .A3(N2361), .A4(N2104) );
  NAND2_X1 NAND5_735( .ZN(N2629), .A1(extra27), .A2(N926) );
  NAND4_X1 NAND5_736_A( .ZN(extra28), .A1(N2386), .A2(N2427), .A3(N2340), .A4(N2129) );
  NAND2_X1 NAND5_736( .ZN(N2630), .A1(extra28), .A2(N926) );
  NAND4_X1 NAND5_737_A( .ZN(extra29), .A1(N2386), .A2(N2427), .A3(N2340), .A4(N2119) );
  NAND2_X1 NAND5_737( .ZN(N2631), .A1(extra29), .A2(N926) );
  NAND4_X1 NAND5_738_A( .ZN(extra30), .A1(N2386), .A2(N2427), .A3(N2353), .A4(N2104) );
  NAND2_X1 NAND5_738( .ZN(N2632), .A1(extra30), .A2(N926) );
  NAND4_X1 NAND5_739_A( .ZN(extra31), .A1(N2386), .A2(N2426), .A3(N2340), .A4(N2104) );
  NAND2_X1 NAND5_739( .ZN(N2633), .A1(extra31), .A2(N926) );
  NAND4_X1 NAND5_740_A( .ZN(extra32), .A1(N2385), .A2(N2427), .A3(N2340), .A4(N2104) );
  NAND2_X1 NAND5_740( .ZN(N2634), .A1(extra32), .A2(N926) );
  AND4_X1 AND5_741_A( .ZN(extra33), .A1(N2286), .A2(N2427), .A3(N2361), .A4(N2129) );
  AND2_X1 AND5_741( .ZN(N2639), .A1(extra33), .A2(N1171) );
  AND4_X1 AND5_742_A( .ZN(extra34), .A1(N2297), .A2(N2427), .A3(N2361), .A4(N2119) );
  AND2_X1 AND5_742( .ZN(N2642), .A1(extra34), .A2(N1171) );
  AND4_X1 AND5_743_A( .ZN(extra35), .A1(N2297), .A2(N2427), .A3(N2375), .A4(N2104) );
  AND2_X1 AND5_743( .ZN(N2645), .A1(extra35), .A2(N1171) );
  AND4_X1 AND5_744_A( .ZN(extra36), .A1(N2297), .A2(N2427), .A3(N2340), .A4(N2143) );
  AND2_X1 AND5_744( .ZN(N2648), .A1(extra36), .A2(N1171) );
  AND4_X1 AND5_745_A( .ZN(extra37), .A1(N2297), .A2(N2427), .A3(N2353), .A4(N2129) );
  AND2_X1 AND5_745( .ZN(N2651), .A1(extra37), .A2(N1188) );
  AND4_X1 AND5_746_A( .ZN(extra38), .A1(N2386), .A2(N2326), .A3(N2361), .A4(N2129) );
  AND2_X1 AND5_746( .ZN(N2655), .A1(extra38), .A2(N1188) );
  AND4_X1 AND5_747_A( .ZN(extra39), .A1(N2386), .A2(N2326), .A3(N2361), .A4(N2119) );
  AND2_X1 AND5_747( .ZN(N2658), .A1(extra39), .A2(N1188) );
  AND4_X1 AND5_748_A( .ZN(extra40), .A1(N2386), .A2(N2326), .A3(N2375), .A4(N2104) );
  AND2_X1 AND5_748( .ZN(N2661), .A1(extra40), .A2(N1188) );
  AND4_X1 AND5_749_A( .ZN(extra41), .A1(N2386), .A2(N2326), .A3(N2353), .A4(N2129) );
  AND2_X1 AND5_749( .ZN(N2664), .A1(extra41), .A2(N1188) );
  NAND2_X1 NAND2_750( .ZN(N2669), .A1(N2558), .A2(N534) );
  INV_X1 NOT1_751( .ZN(N2670), .A(N2558) );
  NAND2_X1 NAND2_752( .ZN(N2671), .A1(N2561), .A2(N535) );
  INV_X1 NOT1_753( .ZN(N2672), .A(N2561) );
  NAND2_X1 NAND2_754( .ZN(N2673), .A1(N2564), .A2(N536) );
  INV_X1 NOT1_755( .ZN(N2674), .A(N2564) );
  NAND2_X1 NAND2_756( .ZN(N2675), .A1(N2567), .A2(N537) );
  INV_X1 NOT1_757( .ZN(N2676), .A(N2567) );
  NAND2_X1 NAND2_758( .ZN(N2682), .A1(N2570), .A2(N543) );
  INV_X1 NOT1_759( .ZN(N2683), .A(N2570) );
  NAND2_X1 NAND2_760( .ZN(N2688), .A1(N2573), .A2(N548) );
  INV_X1 NOT1_761( .ZN(N2689), .A(N2573) );
  NAND2_X1 NAND2_762( .ZN(N2690), .A1(N2576), .A2(N549) );
  INV_X1 NOT1_763( .ZN(N2691), .A(N2576) );
  AND4_X1 AND8_764_A( .ZN(extra42), .A1(N2627), .A2(N2628), .A3(N2629), .A4(N2630) );
  AND4_X1 AND8_764_B( .ZN(extra43), .A1(extra42), .A2(N2631), .A3(N2632), .A4(N2633) );
  AND2_X1 AND8_764( .ZN(N2710), .A1(extra43), .A2(N2634) );
  NAND2_X1 NAND2_765( .ZN(N2720), .A1(N343), .A2(N2670) );
  NAND2_X1 NAND2_766( .ZN(N2721), .A1(N346), .A2(N2672) );
  NAND2_X1 NAND2_767( .ZN(N2722), .A1(N349), .A2(N2674) );
  NAND2_X1 NAND2_768( .ZN(N2723), .A1(N352), .A2(N2676) );
  NAND2_X1 NAND2_769( .ZN(N2724), .A1(N2639), .A2(N538) );
  INV_X1 NOT1_770( .ZN(N2725), .A(N2639) );
  NAND2_X1 NAND2_771( .ZN(N2726), .A1(N2642), .A2(N539) );
  INV_X1 NOT1_772( .ZN(N2727), .A(N2642) );
  NAND2_X1 NAND2_773( .ZN(N2728), .A1(N2645), .A2(N540) );
  INV_X1 NOT1_774( .ZN(N2729), .A(N2645) );
  NAND2_X1 NAND2_775( .ZN(N2730), .A1(N2648), .A2(N541) );
  INV_X4 NOT1_776( .ZN(N2731), .A(N2648) );
  NAND2_X1 NAND2_777( .ZN(N2732), .A1(N2651), .A2(N542) );
  INV_X1 NOT1_778( .ZN(N2733), .A(N2651) );
  NAND2_X1 NAND2_779( .ZN(N2734), .A1(N370), .A2(N2683) );
  NAND2_X1 NAND2_780( .ZN(N2735), .A1(N2655), .A2(N544) );
  INV_X1 NOT1_781( .ZN(N2736), .A(N2655) );
  NAND2_X1 NAND2_782( .ZN(N2737), .A1(N2658), .A2(N545) );
  INV_X1 NOT1_783( .ZN(N2738), .A(N2658) );
  NAND2_X1 NAND2_784( .ZN(N2739), .A1(N2661), .A2(N546) );
  INV_X1 NOT1_785( .ZN(N2740), .A(N2661) );
  NAND2_X1 NAND2_786( .ZN(N2741), .A1(N2664), .A2(N547) );
  INV_X1 NOT1_787( .ZN(N2742), .A(N2664) );
  NAND2_X1 NAND2_788( .ZN(N2743), .A1(N385), .A2(N2689) );
  NAND2_X1 NAND2_789( .ZN(N2744), .A1(N388), .A2(N2691) );
  NAND4_X1 NAND8_790_A( .ZN(extra44), .A1(N2537), .A2(N2540), .A3(N2543), .A4(N2546) );
  NAND4_X1 NAND8_790_B( .ZN(extra45), .A1(extra44), .A2(N2594), .A3(N2597), .A4(N2600) );
  NAND2_X1 NAND8_790( .ZN(N2745), .A1(extra45), .A2(N2603) );
  NAND4_X1 NAND8_791_A( .ZN(extra46), .A1(N2606), .A2(N2549), .A3(N2611), .A4(N2614) );
  NAND4_X1 NAND8_791_B( .ZN(extra47), .A1(extra46), .A2(N2617), .A3(N2620), .A4(N2552) );
  NAND2_X1 NAND8_791( .ZN(N2746), .A1(extra47), .A2(N2555) );
  AND4_X1 AND8_792_A( .ZN(extra48), .A1(N2537), .A2(N2540), .A3(N2543), .A4(N2546) );
  AND4_X1 AND8_792_B( .ZN(extra49), .A1(extra48), .A2(N2594), .A3(N2597), .A4(N2600) );
  AND2_X1 AND8_792( .ZN(N2747), .A1(extra49), .A2(N2603) );
  AND4_X1 AND8_793_A( .ZN(extra50), .A1(N2606), .A2(N2549), .A3(N2611), .A4(N2614) );
  AND4_X1 AND8_793_B( .ZN(extra51), .A1(extra50), .A2(N2617), .A3(N2620), .A4(N2552) );
  AND2_X1 AND8_793( .ZN(N2750), .A1(extra51), .A2(N2555) );
  NAND2_X1 NAND2_794( .ZN(N2753), .A1(N2669), .A2(N2720) );
  NAND2_X1 NAND2_795( .ZN(N2754), .A1(N2671), .A2(N2721) );
  NAND2_X1 NAND2_796( .ZN(N2755), .A1(N2673), .A2(N2722) );
  NAND2_X1 NAND2_797( .ZN(N2756), .A1(N2675), .A2(N2723) );
  NAND2_X1 NAND2_798( .ZN(N2757), .A1(N355), .A2(N2725) );
  NAND2_X1 NAND2_799( .ZN(N2758), .A1(N358), .A2(N2727) );
  NAND2_X1 NAND2_800( .ZN(N2759), .A1(N361), .A2(N2729) );
  NAND2_X1 NAND2_801( .ZN(N2760), .A1(N364), .A2(N2731) );
  NAND2_X1 NAND2_802( .ZN(N2761), .A1(N367), .A2(N2733) );
  NAND2_X1 NAND2_803( .ZN(N2762), .A1(N2682), .A2(N2734) );
  NAND2_X1 NAND2_804( .ZN(N2763), .A1(N373), .A2(N2736) );
  NAND2_X1 NAND2_805( .ZN(N2764), .A1(N376), .A2(N2738) );
  NAND2_X1 NAND2_806( .ZN(N2765), .A1(N379), .A2(N2740) );
  NAND2_X1 NAND2_807( .ZN(N2766), .A1(N382), .A2(N2742) );
  NAND2_X1 NAND2_808( .ZN(N2767), .A1(N2688), .A2(N2743) );
  NAND2_X1 NAND2_809( .ZN(N2768), .A1(N2690), .A2(N2744) );
  AND2_X1 AND2_810( .ZN(N2773), .A1(N2745), .A2(N275) );
  AND2_X1 AND2_811( .ZN(N2776), .A1(N2746), .A2(N276) );
  NAND2_X1 NAND2_812( .ZN(N2779), .A1(N2724), .A2(N2757) );
  NAND2_X1 NAND2_813( .ZN(N2780), .A1(N2726), .A2(N2758) );
  NAND2_X1 NAND2_814( .ZN(N2781), .A1(N2728), .A2(N2759) );
  NAND2_X1 NAND2_815( .ZN(N2782), .A1(N2730), .A2(N2760) );
  NAND2_X1 NAND2_816( .ZN(N2783), .A1(N2732), .A2(N2761) );
  NAND2_X1 NAND2_817( .ZN(N2784), .A1(N2735), .A2(N2763) );
  NAND2_X1 NAND2_818( .ZN(N2785), .A1(N2737), .A2(N2764) );
  NAND2_X1 NAND2_819( .ZN(N2786), .A1(N2739), .A2(N2765) );
  NAND2_X1 NAND2_820( .ZN(N2787), .A1(N2741), .A2(N2766) );
  AND3_X1 AND3_821( .ZN(N2788), .A1(N2747), .A2(N2750), .A3(N2710) );
  NAND2_X1 NAND2_822( .ZN(N2789), .A1(N2747), .A2(N2750) );
  AND4_X1 AND4_823( .ZN(N2800), .A1(N338), .A2(N2279), .A3(N99), .A4(N2788) );
  NAND2_X1 NAND2_824( .ZN(N2807), .A1(N2773), .A2(N2018) );
  INV_X1 NOT1_825( .ZN(N2808), .A(N2773) );
  NAND2_X1 NAND2_826( .ZN(N2809), .A1(N2776), .A2(N2019) );
  INV_X1 NOT1_827( .ZN(N2810), .A(N2776) );
  NOR2_X1 NOR2_828( .ZN(N2811), .A1(N2384), .A2(N2800) );
  AND3_X1 AND3_829( .ZN(N2812), .A1(N897), .A2(N283), .A3(N2789) );
  AND3_X1 AND3_830( .ZN(N2815), .A1(N76), .A2(N283), .A3(N2789) );
  AND3_X1 AND3_831( .ZN(N2818), .A1(N82), .A2(N283), .A3(N2789) );
  AND3_X1 AND3_832( .ZN(N2821), .A1(N85), .A2(N283), .A3(N2789) );
  AND3_X1 AND3_833( .ZN(N2824), .A1(N898), .A2(N283), .A3(N2789) );
  NAND2_X1 NAND2_834( .ZN(N2827), .A1(N1965), .A2(N2808) );
  NAND2_X1 NAND2_835( .ZN(N2828), .A1(N1968), .A2(N2810) );
  AND3_X1 AND3_836( .ZN(N2829), .A1(N79), .A2(N283), .A3(N2789) );
  NAND2_X1 NAND2_837( .ZN(N2843), .A1(N2807), .A2(N2827) );
  NAND2_X1 NAND2_838( .ZN(N2846), .A1(N2809), .A2(N2828) );
  NAND2_X1 NAND2_839( .ZN(N2850), .A1(N2812), .A2(N2076) );
  NAND2_X1 NAND2_840( .ZN(N2851), .A1(N2815), .A2(N2077) );
  NAND2_X1 NAND2_841( .ZN(N2852), .A1(N2818), .A2(N1915) );
  NAND2_X1 NAND2_842( .ZN(N2853), .A1(N2821), .A2(N1857) );
  NAND2_X1 NAND2_843( .ZN(N2854), .A1(N2824), .A2(N1938) );
  INV_X1 NOT1_844( .ZN(N2857), .A(N2812) );
  INV_X1 NOT1_845( .ZN(N2858), .A(N2815) );
  INV_X1 NOT1_846( .ZN(N2859), .A(N2818) );
  INV_X1 NOT1_847( .ZN(N2860), .A(N2821) );
  INV_X1 NOT1_848( .ZN(N2861), .A(N2824) );
  INV_X1 NOT1_849( .ZN(N2862), .A(N2829) );
  NAND2_X1 NAND2_850( .ZN(N2863), .A1(N2829), .A2(N1985) );
  NAND2_X1 NAND2_851( .ZN(N2866), .A1(N2052), .A2(N2857) );
  NAND2_X1 NAND2_852( .ZN(N2867), .A1(N2055), .A2(N2858) );
  NAND2_X1 NAND2_853( .ZN(N2868), .A1(N1866), .A2(N2859) );
  NAND2_X1 NAND2_854( .ZN(N2869), .A1(N1818), .A2(N2860) );
  NAND2_X1 NAND2_855( .ZN(N2870), .A1(N1902), .A2(N2861) );
  NAND2_X1 NAND2_856( .ZN(N2871), .A1(N2843), .A2(N886) );
  INV_X1 NOT1_857( .ZN(N2872), .A(N2843) );
  NAND2_X1 NAND2_858( .ZN(N2873), .A1(N2846), .A2(N887) );
  INV_X1 NOT1_859( .ZN(N2874), .A(N2846) );
  NAND2_X1 NAND2_860( .ZN(N2875), .A1(N1933), .A2(N2862) );
  NAND2_X1 NAND2_861( .ZN(N2876), .A1(N2866), .A2(N2850) );
  NAND2_X1 NAND2_862( .ZN(N2877), .A1(N2867), .A2(N2851) );
  NAND2_X1 NAND2_863( .ZN(N2878), .A1(N2868), .A2(N2852) );
  NAND2_X1 NAND2_864( .ZN(N2879), .A1(N2869), .A2(N2853) );
  NAND2_X1 NAND2_865( .ZN(N2880), .A1(N2870), .A2(N2854) );
  NAND2_X1 NAND2_866( .ZN(N2881), .A1(N682), .A2(N2872) );
  NAND2_X1 NAND2_867( .ZN(N2882), .A1(N685), .A2(N2874) );
  NAND2_X1 NAND2_868( .ZN(N2883), .A1(N2875), .A2(N2863) );
  AND2_X1 AND2_869( .ZN(N2886), .A1(N2876), .A2(N550) );
  AND2_X1 AND2_870( .ZN(N2887), .A1(N551), .A2(N2877) );
  AND2_X1 AND2_871( .ZN(N2888), .A1(N553), .A2(N2878) );
  AND2_X1 AND2_872( .ZN(N2889), .A1(N2879), .A2(N554) );
  AND2_X1 AND2_873( .ZN(N2890), .A1(N555), .A2(N2880) );
  NAND2_X1 NAND2_874( .ZN(N2891), .A1(N2871), .A2(N2881) );
  NAND2_X1 NAND2_875( .ZN(N2892), .A1(N2873), .A2(N2882) );
  NAND2_X1 NAND2_876( .ZN(N2895), .A1(N2883), .A2(N1461) );
  INV_X1 NOT1_877( .ZN(N2896), .A(N2883) );
  NAND2_X1 NAND2_878( .ZN(N2897), .A1(N1383), .A2(N2896) );
  NAND2_X1 NAND2_879( .ZN(N2898), .A1(N2895), .A2(N2897) );
  AND2_X1 AND2_880( .ZN(N2899), .A1(N2898), .A2(N552) );

endmodule
