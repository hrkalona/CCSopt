// Verilog
// c7552
// Ninputs 207
// Noutputs 108
// NtotalGates 3513
// BUFF1 535
// NOT1 876
// AND2 534
// AND4 64
// NAND2 1028
// NOR2 40
// OR2 180
// OR3 10
// AND5 32
// AND3 146
// OR5 24
// OR4 30
// NOR3 10
// NOR4 4

module c7552(N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,N35,N38,N41,N44,N47,N50,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N69,N70,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,N97,N100,N103,N106,
  N109,N110,N111,N112,N113,N114,N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,N141,N144,
  N147,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,
  N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,
  N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,
  N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N242,N245,N248,N251,N254,N257,N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
  N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,
  N349,N352,N355,N358,N361,N364,N367,N382,N241_I,N387,N388,N478,N482,N484,N486,N489,N492,N501,
  N505,N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,N541,N543,N545,N547,N549,N551,N553,
  N556,N559,N561,N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,N881,N882,N883,N884,N885,
  N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,N10109,N10110,N10111,
  N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,N10715,
  N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,
  N10905,N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O);
input N1,N5,N9,N12,N15,N18,N23,N26,N29,N32,N35,N38,N41,N44,N47,N50,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N69,N70,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N94,N97,N100,N103,N106,N109,N110,N111,N112,N113,N114,
  N115,N118,N121,N124,N127,N130,N133,N134,N135,N138,N141,N144,N147,N150,N151,N152,N153,N154,N155,N156,
  N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
  N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,N240,N242,N245,N248,N251,N254,N257,N260,N263,N267,N271,N274,N277,N280,N283,N286,N289,
  N293,N296,N299,N303,N307,N310,N313,N316,N319,N322,N325,N328,N331,N334,N337,N340,N343,N346,N349,N352,
  N355,N358,N361,N364,N367,N382,N241_I;
output N387,N388,N478,N482,N484,N486,N489,N492,N501,N505,N507,N509,N511,N513,N515,N517,N519,N535,N537,N539,
  N541,N543,N545,N547,N549,N551,N553,N556,N559,N561,N563,N565,N567,N569,N571,N573,N582,N643,N707,N813,
  N881,N882,N883,N884,N885,N889,N945,N1110,N1111,N1112,N1113,N1114,N1489,N1490,N1781,N10025,N10101,N10102,N10103,N10104,
  N10109,N10110,N10111,N10112,N10350,N10351,N10352,N10353,N10574,N10575,N10576,N10628,N10632,N10641,N10704,N10706,N10711,N10712,N10713,N10714,
  N10715,N10716,N10717,N10718,N10729,N10759,N10760,N10761,N10762,N10763,N10827,N10837,N10838,N10839,N10840,N10868,N10869,N10870,N10871,N10905,
  N10906,N10907,N10908,N11333,N11334,N11340,N11342,N241_O;

  wire N467,N469,N494,N528,N575,N578,N585,N590,N593,N596,N599,N604,N609,N614,N625,N628,
    N632,N636,N641,N642,N644,N651,N657,N660,N666,N672,N673,N674,N676,N682,N688,N689,
    N695,N700,N705,N706,N708,N715,N721,N727,N733,N734,N742,N748,N749,N750,N758,N759,
    N762,N768,N774,N780,N786,N794,N800,N806,N812,N814,N821,N827,N833,N839,N845,N853,
    N859,N865,N871,N886,N887,N957,N1028,N1029,N1109,N1115,N1116,N1119,N1125,N1132,N1136,N1141,
    N1147,N1154,N1160,N1167,N1174,N1175,N1182,N1189,N1194,N1199,N1206,N1211,N1218,N1222,N1227,N1233,
    N1240,N1244,N1249,N1256,N1263,N1270,N1277,N1284,N1287,N1290,N1293,N1296,N1299,N1302,N1305,N1308,
    N1311,N1314,N1317,N1320,N1323,N1326,N1329,N1332,N1335,N1338,N1341,N1344,N1347,N1350,N1353,N1356,
    N1359,N1362,N1365,N1368,N1371,N1374,N1377,N1380,N1383,N1386,N1389,N1392,N1395,N1398,N1401,N1404,
    N1407,N1410,N1413,N1416,N1419,N1422,N1425,N1428,N1431,N1434,N1437,N1440,N1443,N1446,N1449,N1452,
    N1455,N1458,N1461,N1464,N1467,N1470,N1473,N1476,N1479,N1482,N1485,N1537,N1551,N1649,N1703,N1708,
    N1713,N1721,N1758,N1782,N1783,N1789,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1805,N1811,N1812,
    N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1828,N1829,N1830,N1832,N1833,N1834,
    N1835,N1839,N1840,N1841,N1842,N1843,N1845,N1851,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
    N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,
    N1881,N1882,N1883,N1884,N1885,N1892,N1899,N1906,N1913,N1919,N1926,N1927,N1928,N1929,N1930,N1931,
    N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,
    N1953,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,
    N1973,N1974,N1975,N1976,N1977,N1983,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N2003,
    N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2031,
    N2038,N2045,N2052,N2058,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2081,
    N2086,N2107,N2108,N2110,N2111,N2112,N2113,N2114,N2115,N2117,N2171,N2172,N2230,N2231,N2235,N2239,
    N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,
    N2256,N2257,N2267,N2268,N2269,N2274,N2275,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,
    N2286,N2287,N2293,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2315,N2321,
    N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2337,N2338,N2339,N2340,N2341,N2342,
    N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,
    N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2374,N2375,N2376,N2377,N2378,N2379,
    N2380,N2381,N2382,N2383,N2384,N2390,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,
    N2406,N2412,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
    N2432,N2433,N2434,N2435,N2436,N2437,N2441,N2442,N2446,N2450,N2454,N2458,N2462,N2466,N2470,N2474,
    N2478,N2482,N2488,N2496,N2502,N2508,N2523,N2533,N2537,N2538,N2542,N2546,N2550,N2554,N2561,N2567,
    N2573,N2604,N2607,N2611,N2615,N2619,N2626,N2632,N2638,N2644,N2650,N2653,N2654,N2658,N2662,N2666,
    N2670,N2674,N2680,N2688,N2692,N2696,N2700,N2704,N2728,N2729,N2733,N2737,N2741,N2745,N2749,N2753,
    N2757,N2761,N2765,N2766,N2769,N2772,N2775,N2778,N2781,N2784,N2787,N2790,N2793,N2796,N2866,N2867,
    N2868,N2869,N2878,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,
    N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2988,N3005,N3006,N3007,
    N3008,N3009,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3032,N3033,N3034,N3035,
    N3036,N3037,N3038,N3039,N3040,N3041,N3061,N3064,N3067,N3070,N3073,N3080,N3096,N3097,N3101,N3107,
    N3114,N3122,N3126,N3130,N3131,N3134,N3135,N3136,N3137,N3140,N3144,N3149,N3155,N3159,N3167,N3168,
    N3169,N3173,N3178,N3184,N3185,N3189,N3195,N3202,N3210,N3211,N3215,N3221,N3228,N3229,N3232,N3236,
    N3241,N3247,N3251,N3255,N3259,N3263,N3267,N3273,N3281,N3287,N3293,N3299,N3303,N3307,N3311,N3315,
    N3322,N3328,N3334,N3340,N3343,N3349,N3355,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,
    N3370,N3371,N3372,N3373,N3374,N3375,N3379,N3380,N3381,N3384,N3390,N3398,N3404,N3410,N3416,N3420,
    N3424,N3428,N3432,N3436,N3440,N3444,N3448,N3452,N3453,N3454,N3458,N3462,N3466,N3470,N3474,N3478,
    N3482,N3486,N3487,N3490,N3493,N3496,N3499,N3502,N3507,N3510,N3515,N3518,N3521,N3524,N3527,N3530,
    N3535,N3539,N3542,N3545,N3548,N3551,N3552,N3553,N3557,N3560,N3563,N3566,N3569,N3570,N3571,N3574,
    N3577,N3580,N3583,N3586,N3589,N3592,N3595,N3598,N3601,N3604,N3607,N3610,N3613,N3616,N3619,N3622,
    N3625,N3628,N3631,N3634,N3637,N3640,N3643,N3646,N3649,N3652,N3655,N3658,N3661,N3664,N3667,N3670,
    N3673,N3676,N3679,N3682,N3685,N3688,N3691,N3694,N3697,N3700,N3703,N3706,N3709,N3712,N3715,N3718,
    N3721,N3724,N3727,N3730,N3733,N3736,N3739,N3742,N3745,N3748,N3751,N3754,N3757,N3760,N3763,N3766,
    N3769,N3772,N3775,N3778,N3781,N3782,N3783,N3786,N3789,N3792,N3795,N3798,N3801,N3804,N3807,N3810,
    N3813,N3816,N3819,N3822,N3825,N3828,N3831,N3834,N3837,N3840,N3843,N3846,N3849,N3852,N3855,N3858,
    N3861,N3864,N3867,N3870,N3873,N3876,N3879,N3882,N3885,N3888,N3891,N3953,N3954,N3955,N3956,N3958,
    N3964,N4193,N4303,N4308,N4313,N4326,N4327,N4333,N4334,N4411,N4412,N4463,N4464,N4465,N4466,N4467,
    N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,
    N4484,N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,
    N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,
    N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531,
    N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4549,N4555,
    N4562,N4563,N4566,N4570,N4575,N4576,N4577,N4581,N4586,N4592,N4593,N4597,N4603,N4610,N4611,N4612,
    N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,
    N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,
    N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4656,N4657,N4661,N4667,N4674,N4675,N4678,
    N4682,N4687,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4706,N4711,N4717,N4718,
    N4722,N4728,N4735,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,
    N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4775,N4776,
    N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,N4789,N4790,N4793,N4794,N4795,N4796,N4799,N4800,
    N4801,N4802,N4803,N4806,N4809,N4810,N4813,N4814,N4817,N4820,N4823,N4826,N4829,N4832,N4835,N4838,
    N4841,N4844,N4847,N4850,N4853,N4856,N4859,N4862,N4865,N4868,N4871,N4874,N4877,N4880,N4883,N4886,
    N4889,N4892,N4895,N4898,N4901,N4904,N4907,N4910,N4913,N4916,N4919,N4922,N4925,N4928,N4931,N4934,
    N4937,N4940,N4943,N4946,N4949,N4952,N4955,N4958,N4961,N4964,N4967,N4970,N4973,N4976,N4979,N4982,
    N4985,N4988,N4991,N4994,N4997,N5000,N5003,N5006,N5009,N5012,N5015,N5018,N5021,N5024,N5027,N5030,
    N5033,N5036,N5039,N5042,N5045,N5046,N5047,N5048,N5049,N5052,N5055,N5058,N5061,N5064,N5065,N5066,
    N5067,N5068,N5071,N5074,N5077,N5080,N5083,N5086,N5089,N5092,N5095,N5098,N5101,N5104,N5107,N5110,
    N5111,N5112,N5113,N5114,N5117,N5120,N5123,N5126,N5129,N5132,N5135,N5138,N5141,N5144,N5147,N5150,
    N5153,N5156,N5159,N5162,N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,
    N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,
    N5193,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,
    N5211,N5212,N5213,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,
    N5296,N5297,N5298,N5299,N5300,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,
    N5363,N5364,N5365,N5366,N5367,N5425,N5426,N5427,N5429,N5430,N5431,N5432,N5433,N5451,N5452,N5453,
    N5454,N5455,N5456,N5457,N5469,N5474,N5475,N5476,N5477,N5571,N5572,N5573,N5574,N5584,N5585,N5586,
    N5587,N5602,N5603,N5604,N5605,N5631,N5632,N5640,N5654,N5670,N5683,N5690,N5697,N5707,N5718,N5728,
    N5735,N5736,N5740,N5744,N5747,N5751,N5755,N5758,N5762,N5766,N5769,N5770,N5771,N5778,N5789,N5799,
    N5807,N5821,N5837,N5850,N5856,N5863,N5870,N5881,N5892,N5898,N5905,N5915,N5926,N5936,N5943,N5944,
    N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,
    N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,
    N5989,N5990,N5991,N5996,N6000,N6003,N6009,N6014,N6018,N6021,N6022,N6023,N6024,N6025,N6026,N6027,
    N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6047,N6052,
    N6056,N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,
    N6074,N6075,N6076,N6077,N6078,N6079,N6083,N6087,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,
    N6098,N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,
    N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6131,N6135,
    N6136,N6137,N6141,N6145,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,
    N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6170,N6174,N6177,N6181,N6182,N6183,N6184,N6185,N6186,
    N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6199,N6202,N6203,N6204,N6207,N6210,
    N6213,N6214,N6217,N6220,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6235,N6236,
    N6239,N6240,N6241,N6242,N6243,N6246,N6249,N6252,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,
    N6263,N6266,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6555,N6556,N6557,N6558,N6559,N6560,
    N6561,N6569,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6621,
    N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,
    N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6668,
    N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,N6702,N6703,
    N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6729,N6730,N6731,N6732,N6733,N6734,N6735,
    N6736,N6741,N6742,N6743,N6744,N6751,N6752,N6753,N6754,N6755,N6756,N6757,N6758,N6761,N6762,N6766,
    N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,
    N6783,N6784,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,N6800,N6803,N6806,
    N6809,N6812,N6815,N6818,N6821,N6824,N6827,N6830,N6833,N6836,N6837,N6838,N6839,N6840,N6841,N6842,
    N6843,N6844,N6845,N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,
    N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,N6878,
    N6879,N6880,N6881,N6884,N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6901,N6912,
    N6923,N6929,N6936,N6946,N6957,N6967,N6968,N6969,N6970,N6977,N6988,N6998,N7006,N7020,N7036,N7049,
    N7055,N7056,N7057,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7073,N7077,N7080,N7086,
    N7091,N7095,N7098,N7099,N7100,N7103,N7104,N7105,N7106,N7107,N7114,N7125,N7136,N7142,N7149,N7159,
    N7170,N7180,N7187,N7188,N7191,N7194,N7198,N7202,N7205,N7209,N7213,N7216,N7219,N7222,N7229,N7240,
    N7250,N7258,N7272,N7288,N7301,N7307,N7314,N7318,N7322,N7325,N7328,N7331,N7334,N7337,N7340,N7343,
    N7346,N7351,N7355,N7358,N7364,N7369,N7373,N7376,N7377,N7378,N7381,N7384,N7387,N7391,N7394,N7398,
    N7402,N7405,N7408,N7411,N7414,N7417,N7420,N7423,N7426,N7429,N7432,N7435,N7438,N7441,N7444,N7447,
    N7450,N7453,N7456,N7459,N7462,N7465,N7468,N7471,N7474,N7477,N7478,N7479,N7482,N7485,N7488,N7491,
    N7494,N7497,N7500,N7503,N7506,N7509,N7512,N7515,N7518,N7521,N7524,N7527,N7530,N7533,N7536,N7539,
    N7542,N7545,N7548,N7551,N7552,N7553,N7556,N7557,N7558,N7559,N7560,N7563,N7566,N7569,N7572,N7573,
    N7574,N7577,N7580,N7581,N7582,N7585,N7588,N7591,N7609,N7613,N7620,N7649,N7650,N7655,N7659,N7668,
    N7671,N7744,N7822,N7825,N7826,N7852,N8114,N8117,N8131,N8134,N8144,N8145,N8146,N8156,N8166,N8169,
    N8183,N8186,N8196,N8200,N8204,N8208,N8216,N8217,N8218,N8219,N8232,N8233,N8242,N8243,N8244,N8245,
    N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8260,N8261,N8262,N8269,N8274,N8275,N8276,
    N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8288,N8294,N8295,N8296,N8297,N8298,N8307,
    N8315,N8317,N8319,N8321,N8322,N8323,N8324,N8325,N8326,N8333,N8337,N8338,N8339,N8340,N8341,N8342,
    N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,N8356,N8357,N8358,
    N8365,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,N8383,
    N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8404,N8405,N8409,N8410,N8411,
    N8412,N8415,N8416,N8417,N8418,N8421,N8430,N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,
    N8442,N8443,N8444,N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8460,N8463,
    N8466,N8469,N8470,N8471,N8474,N8477,N8480,N8483,N8484,N8485,N8488,N8489,N8490,N8491,N8492,N8493,
    N8494,N8495,N8496,N8497,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,
    N8512,N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8522,N8525,N8528,N8531,N8534,N8537,N8538,N8539,
    N8540,N8541,N8545,N8546,N8547,N8548,N8551,N8552,N8553,N8554,N8555,N8558,N8561,N8564,N8565,N8566,
    N8569,N8572,N8575,N8578,N8579,N8580,N8583,N8586,N8589,N8592,N8595,N8598,N8601,N8604,N8607,N8608,
    N8609,N8610,N8615,N8616,N8617,N8618,N8619,N8624,N8625,N8626,N8627,N8632,N8633,N8634,N8637,N8638,
    N8639,N8644,N8645,N8646,N8647,N8648,N8653,N8654,N8655,N8660,N8663,N8666,N8669,N8672,N8675,N8678,
    N8681,N8684,N8687,N8690,N8693,N8696,N8699,N8702,N8705,N8708,N8711,N8714,N8717,N8718,N8721,N8724,
    N8727,N8730,N8733,N8734,N8735,N8738,N8741,N8744,N8747,N8750,N8753,N8754,N8755,N8756,N8757,N8760,
    N8763,N8766,N8769,N8772,N8775,N8778,N8781,N8784,N8787,N8790,N8793,N8796,N8799,N8802,N8805,N8808,
    N8811,N8814,N8815,N8816,N8817,N8818,N8840,N8857,N8861,N8862,N8863,N8864,N8865,N8866,N8871,N8874,
    N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8898,N8902,N8920,N8924,N8927,
    N8931,N8943,N8950,N8956,N8959,N8960,N8963,N8966,N8991,N8992,N8995,N8996,N9001,N9005,N9024,N9025,
    N9029,N9035,N9053,N9054,N9064,N9065,N9066,N9067,N9068,N9071,N9072,N9073,N9074,N9077,N9079,N9082,
    N9083,N9086,N9087,N9088,N9089,N9092,N9093,N9094,N9095,N9098,N9099,N9103,N9107,N9111,N9117,N9127,
    N9146,N9149,N9159,N9160,N9161,N9165,N9169,N9173,N9179,N9180,N9181,N9182,N9183,N9193,N9203,N9206,
    N9220,N9223,N9234,N9235,N9236,N9237,N9238,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,N9250,
    N9251,N9252,N9256,N9257,N9258,N9259,N9260,N9261,N9262,N9265,N9268,N9271,N9272,N9273,N9274,N9275,
    N9276,N9280,N9285,N9286,N9287,N9288,N9290,N9292,N9294,N9296,N9297,N9298,N9299,N9300,N9301,N9307,
    N9314,N9315,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9326,N9332,N9339,N9344,N9352,N9354,N9356,
    N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,N9370,N9371,N9372,N9375,
    N9381,N9382,N9383,N9384,N9385,N9392,N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,
    N9407,N9408,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,N9423,N9426,N9429,
    N9432,N9435,N9442,N9445,N9454,N9455,N9456,N9459,N9460,N9461,N9462,N9465,N9466,N9467,N9468,N9473,
    N9476,N9477,N9478,N9485,N9488,N9493,N9494,N9495,N9498,N9499,N9500,N9505,N9506,N9507,N9508,N9509,
    N9514,N9515,N9516,N9517,N9520,N9526,N9531,N9539,N9540,N9541,N9543,N9551,N9555,N9556,N9557,N9560,
    N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,N9570,N9571,N9575,N9579,N9581,N9582,N9585,
    N9591,N9592,N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9608,
    N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9621,N9622,N9623,N9624,N9626,N9629,N9632,N9635,
    N9642,N9645,N9646,N9649,N9650,N9653,N9656,N9659,N9660,N9661,N9662,N9663,N9666,N9667,N9670,N9671,
    N9674,N9675,N9678,N9679,N9682,N9685,N9690,N9691,N9692,N9695,N9698,N9702,N9707,N9710,N9711,N9714,
    N9715,N9716,N9717,N9720,N9721,N9722,N9723,N9726,N9727,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
    N9739,N9740,N9741,N9742,N9754,N9758,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,N9773,N9774,
    N9775,N9779,N9784,N9785,N9786,N9790,N9791,N9795,N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,
    N9805,N9806,N9809,N9813,N9814,N9815,N9816,N9817,N9820,N9825,N9826,N9827,N9828,N9829,N9830,N9835,
    N9836,N9837,N9838,N9846,N9847,N9862,N9863,N9866,N9873,N9876,N9890,N9891,N9892,N9893,N9894,N9895,
    N9896,N9897,N9898,N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,
    N9917,N9923,N9924,N9925,N9932,N9935,N9938,N9939,N9945,N9946,N9947,N9948,N9949,N9953,N9954,N9955,
    N9956,N9957,N9958,N9959,N9960,N9961,N9964,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974,N9975,
    N9976,N9977,N9978,N9979,N9982,N9983,N9986,N9989,N9992,N9995,N9996,N9997,N9998,N9999,N10002,N10003,
    N10006,N10007,N10010,N10013,N10014,N10015,N10016,N10017,N10018,N10019,N10020,N10021,N10022,N10023,N10024,N10026,
    N10028,N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,N10042,N10043,N10050,N10053,N10054,
    N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10067,N10070,N10073,N10076,N10077,N10082,N10083,N10084,
    N10085,N10086,N10093,N10094,N10105,N10106,N10107,N10108,N10113,N10114,N10115,N10116,N10119,N10124,N10130,N10131,
    N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10148,N10155,N10156,N10157,N10158,N10159,
    N10160,N10161,N10162,N10163,N10164,N10165,N10170,N10173,N10176,N10177,N10178,N10179,N10180,N10183,N10186,N10189,
    N10192,N10195,N10196,N10197,N10200,N10203,N10204,N10205,N10206,N10212,N10213,N10230,N10231,N10232,N10233,N10234,
    N10237,N10238,N10239,N10240,N10241,N10242,N10247,N10248,N10259,N10264,N10265,N10266,N10267,N10268,N10269,N10270,
    N10271,N10272,N10273,N10278,N10279,N10280,N10281,N10282,N10283,N10287,N10288,N10289,N10290,N10291,N10292,N10293,
    N10294,N10295,N10296,N10299,N10300,N10301,N10306,N10307,N10308,N10311,N10314,N10315,N10316,N10317,N10318,N10321,
    N10324,N10325,N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10337,N10338,N10339,N10340,N10341,
    N10344,N10354,N10357,N10360,N10367,N10375,N10381,N10388,N10391,N10399,N10402,N10406,N10409,N10412,N10415,N10419,
    N10422,N10425,N10428,N10431,N10432,N10437,N10438,N10439,N10440,N10441,N10444,N10445,N10450,N10451,N10455,N10456,
    N10465,N10466,N10479,N10497,N10509,N10512,N10515,N10516,N10517,N10518,N10519,N10522,N10525,N10528,N10531,N10534,
    N10535,N10536,N10539,N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,
    N10555,N10556,N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,N10568,N10569,N10570,
    N10571,N10572,N10573,N10577,N10581,N10582,N10583,N10587,N10588,N10589,N10594,N10595,N10596,N10597,N10598,N10602,
    N10609,N10610,N10621,N10626,N10627,N10629,N10631,N10637,N10638,N10639,N10640,N10642,N10643,N10644,N10645,N10647,
    N10648,N10649,N10652,N10659,N10662,N10665,N10668,N10671,N10672,N10673,N10674,N10675,N10678,N10681,N10682,N10683,
    N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10694,N10695,N10696,N10697,N10698,N10701,N10705,N10707,
    N10708,N10709,N10710,N10719,N10720,N10730,N10731,N10737,N10738,N10739,N10746,N10747,N10748,N10749,N10750,N10753,
    N10754,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,N10774,N10775,N10776,N10778,N10781,
    N10784,N10789,N10792,N10796,N10797,N10798,N10799,N10800,N10803,N10806,N10809,N10812,N10815,N10816,N10817,N10820,
    N10823,N10824,N10825,N10826,N10832,N10833,N10834,N10835,N10836,N10845,N10846,N10857,N10862,N10863,N10864,N10865,
    N10866,N10867,N10872,N10873,N10874,N10875,N10876,N10879,N10882,N10883,N10884,N10885,N10886,N10887,N10888,N10889,
    N10890,N10891,N10892,N10895,N10896,N10897,N10898,N10899,N10902,N10909,N10910,N10915,N10916,N10917,N10918,N10919,
    N10922,N10923,N10928,N10931,N10934,N10935,N10936,N10937,N10938,N10941,N10944,N10947,N10950,N10953,N10954,N10955,
    N10958,N10961,N10962,N10963,N10964,N10969,N10970,N10981,N10986,N10987,N10988,N10989,N10990,N10991,N10992,N10995,
    N10998,N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11011,N11012,N11013,N11014,N11015,
    N11018,N11023,N11024,N11027,N11028,N11029,N11030,N11031,N11034,N11035,N11040,N11041,N11042,N11043,N11044,N11047,
    N11050,N11053,N11056,N11059,N11062,N11065,N11066,N11067,N11070,N11073,N11074,N11075,N11076,N11077,N11078,N11095,
    N11098,N11099,N11100,N11103,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,N11117,
    N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11127,N11130,N11137,N11138,N11139,N11140,N11141,N11142,N11143,
    N11144,N11145,N11152,N11153,N11154,N11155,N11156,N11159,N11162,N11165,N11168,N11171,N11174,N11177,N11180,N11183,
    N11184,N11185,N11186,N11187,N11188,N11205,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,
    N11220,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11231,N11232,N11233,N11236,N11239,N11242,N11243,
    N11244,N11245,N11246,N11250,N11252,N11257,N11260,N11261,N11262,N11263,N11264,N11265,N11267,N11268,N11269,N11270,
    N11272,N11277,N11278,N11279,N11280,N11282,N11283,N11284,N11285,N11286,N11288,N11289,N11290,N11291,N11292,N11293,
    N11294,N11295,N11296,N11297,N11298,N11299,N11302,N11307,N11308,N11309,N11312,N11313,N11314,N11315,N11316,N11317,
    N11320,N11321,N11323,N11327,N11328,N11329,N11331,N11335,N11336,N11337,N11338,N11339,N11341,extra0,extra1,extra2,
    extra3,extra4,extra5,extra6,extra7,extra8,extra9,extra10,extra11,extra12,extra13,extra14,extra15,extra16,extra17,extra18,
    extra19,extra20,extra21,extra22,extra23,extra24,extra25,extra26,extra27,extra28,extra29,extra30,extra31,extra32,extra33,extra34,
    extra35,extra36,extra37,extra38,extra39,extra40,extra41,extra42,extra43,extra44,extra45,extra46,extra47,extra48,extra49,extra50,
    extra51,extra52,extra53,extra54,extra55,extra56,extra57,extra58,extra59;

  BUF_X2 BUFF1_1( .Z(N387), .A(N1) );
  BUF_X2 BUFF1_2( .Z(N388), .A(N1) );
  INV_X1 NOT1_3( .ZN(N467), .A(N57) );
  AND2_X1 AND2_4( .ZN(N469), .A1(N134), .A2(N133) );
  BUF_X2 BUFF1_5( .Z(N478), .A(N248) );
  BUF_X1 BUFF1_6( .Z(N482), .A(N254) );
  BUF_X1 BUFF1_7( .Z(N484), .A(N257) );
  BUF_X1 BUFF1_8( .Z(N486), .A(N260) );
  BUF_X1 BUFF1_9( .Z(N489), .A(N263) );
  BUF_X1 BUFF1_10( .Z(N492), .A(N267) );
  AND4_X1 AND4_11( .ZN(N494), .A1(N162), .A2(N172), .A3(N188), .A4(N199) );
  BUF_X1 BUFF1_12( .Z(N501), .A(N274) );
  BUF_X1 BUFF1_13( .Z(N505), .A(N280) );
  BUF_X1 BUFF1_14( .Z(N507), .A(N283) );
  BUF_X1 BUFF1_15( .Z(N509), .A(N286) );
  BUF_X1 BUFF1_16( .Z(N511), .A(N289) );
  BUF_X1 BUFF1_17( .Z(N513), .A(N293) );
  BUF_X1 BUFF1_18( .Z(N515), .A(N296) );
  BUF_X1 BUFF1_19( .Z(N517), .A(N299) );
  BUF_X1 BUFF1_20( .Z(N519), .A(N303) );
  AND4_X1 AND4_21( .ZN(N528), .A1(N150), .A2(N184), .A3(N228), .A4(N240) );
  BUF_X1 BUFF1_22( .Z(N535), .A(N307) );
  BUF_X1 BUFF1_23( .Z(N537), .A(N310) );
  BUF_X1 BUFF1_24( .Z(N539), .A(N313) );
  BUF_X1 BUFF1_25( .Z(N541), .A(N316) );
  BUF_X1 BUFF1_26( .Z(N543), .A(N319) );
  BUF_X1 BUFF1_27( .Z(N545), .A(N322) );
  BUF_X1 BUFF1_28( .Z(N547), .A(N325) );
  BUF_X1 BUFF1_29( .Z(N549), .A(N328) );
  BUF_X1 BUFF1_30( .Z(N551), .A(N331) );
  BUF_X1 BUFF1_31( .Z(N553), .A(N334) );
  BUF_X1 BUFF1_32( .Z(N556), .A(N337) );
  BUF_X1 BUFF1_33( .Z(N559), .A(N343) );
  BUF_X1 BUFF1_34( .Z(N561), .A(N346) );
  BUF_X1 BUFF1_35( .Z(N563), .A(N349) );
  BUF_X1 BUFF1_36( .Z(N565), .A(N352) );
  BUF_X1 BUFF1_37( .Z(N567), .A(N355) );
  BUF_X1 BUFF1_38( .Z(N569), .A(N358) );
  BUF_X1 BUFF1_39( .Z(N571), .A(N361) );
  BUF_X1 BUFF1_40( .Z(N573), .A(N364) );
  AND4_X4 AND4_41( .ZN(N575), .A1(N183), .A2(N182), .A3(N185), .A4(N186) );
  AND4_X1 AND4_42( .ZN(N578), .A1(N210), .A2(N152), .A3(N218), .A4(N230) );
  INV_X1 NOT1_43( .ZN(N582), .A(N15) );
  INV_X1 NOT1_44( .ZN(N585), .A(N5) );
  BUF_X1 BUFF1_45( .Z(N590), .A(N1) );
  INV_X1 NOT1_46( .ZN(N593), .A(N5) );
  INV_X1 NOT1_47( .ZN(N596), .A(N5) );
  INV_X1 NOT1_48( .ZN(N599), .A(N289) );
  INV_X1 NOT1_49( .ZN(N604), .A(N299) );
  INV_X1 NOT1_50( .ZN(N609), .A(N303) );
  BUF_X1 BUFF1_51( .Z(N614), .A(N38) );
  BUF_X1 BUFF1_52( .Z(N625), .A(N15) );
  NAND2_X1 NAND2_53( .ZN(N628), .A1(N12), .A2(N9) );
  NAND2_X1 NAND2_54( .ZN(N632), .A1(N12), .A2(N9) );
  BUF_X1 BUFF1_55( .Z(N636), .A(N38) );
  INV_X2 NOT1_56( .ZN(N641), .A(N245) );
  INV_X2 NOT1_57( .ZN(N642), .A(N248) );
  BUF_X1 BUFF1_58( .Z(N643), .A(N251) );
  INV_X1 NOT1_59( .ZN(N644), .A(N251) );
  INV_X1 NOT1_60( .ZN(N651), .A(N254) );
  BUF_X1 BUFF1_61( .Z(N657), .A(N106) );
  INV_X1 NOT1_62( .ZN(N660), .A(N257) );
  INV_X1 NOT1_63( .ZN(N666), .A(N260) );
  INV_X1 NOT1_64( .ZN(N672), .A(N263) );
  INV_X1 NOT1_65( .ZN(N673), .A(N267) );
  INV_X1 NOT1_66( .ZN(N674), .A(N106) );
  BUF_X1 BUFF1_67( .Z(N676), .A(N18) );
  BUF_X1 BUFF1_68( .Z(N682), .A(N18) );
  AND2_X1 AND2_69( .ZN(N688), .A1(N382), .A2(N263) );
  BUF_X1 BUFF1_70( .Z(N689), .A(N18) );
  INV_X1 NOT1_71( .ZN(N695), .A(N18) );
  NAND2_X1 NAND2_72( .ZN(N700), .A1(N382), .A2(N267) );
  INV_X1 NOT1_73( .ZN(N705), .A(N271) );
  INV_X1 NOT1_74( .ZN(N706), .A(N274) );
  BUF_X1 BUFF1_75( .Z(N707), .A(N277) );
  INV_X1 NOT1_76( .ZN(N708), .A(N277) );
  INV_X1 NOT1_77( .ZN(N715), .A(N280) );
  INV_X1 NOT1_78( .ZN(N721), .A(N283) );
  INV_X1 NOT1_79( .ZN(N727), .A(N286) );
  INV_X1 NOT1_80( .ZN(N733), .A(N289) );
  INV_X1 NOT1_81( .ZN(N734), .A(N293) );
  INV_X1 NOT1_82( .ZN(N742), .A(N296) );
  INV_X1 NOT1_83( .ZN(N748), .A(N299) );
  INV_X1 NOT1_84( .ZN(N749), .A(N303) );
  BUF_X1 BUFF1_85( .Z(N750), .A(N367) );
  INV_X1 NOT1_86( .ZN(N758), .A(N307) );
  INV_X1 NOT1_87( .ZN(N759), .A(N310) );
  INV_X1 NOT1_88( .ZN(N762), .A(N313) );
  INV_X1 NOT1_89( .ZN(N768), .A(N316) );
  INV_X1 NOT1_90( .ZN(N774), .A(N319) );
  INV_X1 NOT1_91( .ZN(N780), .A(N322) );
  INV_X1 NOT1_92( .ZN(N786), .A(N325) );
  INV_X1 NOT1_93( .ZN(N794), .A(N328) );
  INV_X1 NOT1_94( .ZN(N800), .A(N331) );
  INV_X1 NOT1_95( .ZN(N806), .A(N334) );
  INV_X1 NOT1_96( .ZN(N812), .A(N337) );
  BUF_X1 BUFF1_97( .Z(N813), .A(N340) );
  INV_X1 NOT1_98( .ZN(N814), .A(N340) );
  INV_X1 NOT1_99( .ZN(N821), .A(N343) );
  INV_X1 NOT1_100( .ZN(N827), .A(N346) );
  INV_X1 NOT1_101( .ZN(N833), .A(N349) );
  INV_X1 NOT1_102( .ZN(N839), .A(N352) );
  INV_X1 NOT1_103( .ZN(N845), .A(N355) );
  INV_X1 NOT1_104( .ZN(N853), .A(N358) );
  INV_X1 NOT1_105( .ZN(N859), .A(N361) );
  INV_X1 NOT1_106( .ZN(N865), .A(N364) );
  BUF_X1 BUFF1_107( .Z(N871), .A(N367) );
  NAND2_X2 NAND2_108( .ZN(N881), .A1(N467), .A2(N585) );
  INV_X1 NOT1_109( .ZN(N882), .A(N528) );
  INV_X1 NOT1_110( .ZN(N883), .A(N578) );
  INV_X1 NOT1_111( .ZN(N884), .A(N575) );
  INV_X1 NOT1_112( .ZN(N885), .A(N494) );
  AND2_X1 AND2_113( .ZN(N886), .A1(N528), .A2(N578) );
  AND2_X1 AND2_114( .ZN(N887), .A1(N575), .A2(N494) );
  BUF_X2 BUFF1_115( .Z(N889), .A(N590) );
  BUF_X2 BUFF1_116( .Z(N945), .A(N657) );
  INV_X1 NOT1_117( .ZN(N957), .A(N688) );
  AND2_X1 AND2_118( .ZN(N1028), .A1(N382), .A2(N641) );
  NAND2_X1 NAND2_119( .ZN(N1029), .A1(N382), .A2(N705) );
  AND2_X1 AND2_120( .ZN(N1109), .A1(N469), .A2(N596) );
  NAND2_X1 NAND2_121( .ZN(N1110), .A1(N242), .A2(N593) );
  INV_X1 NOT1_122( .ZN(N1111), .A(N625) );
  NAND2_X1 NAND2_123( .ZN(N1112), .A1(N242), .A2(N593) );
  NAND2_X1 NAND2_124( .ZN(N1113), .A1(N469), .A2(N596) );
  INV_X1 NOT1_125( .ZN(N1114), .A(N625) );
  INV_X1 NOT1_126( .ZN(N1115), .A(N871) );
  BUF_X1 BUFF1_127( .Z(N1116), .A(N590) );
  BUF_X1 BUFF1_128( .Z(N1119), .A(N628) );
  BUF_X1 BUFF1_129( .Z(N1125), .A(N682) );
  BUF_X1 BUFF1_130( .Z(N1132), .A(N628) );
  BUF_X1 BUFF1_131( .Z(N1136), .A(N682) );
  BUF_X1 BUFF1_132( .Z(N1141), .A(N628) );
  BUF_X1 BUFF1_133( .Z(N1147), .A(N682) );
  BUF_X1 BUFF1_134( .Z(N1154), .A(N632) );
  BUF_X1 BUFF1_135( .Z(N1160), .A(N676) );
  AND2_X1 AND2_136( .ZN(N1167), .A1(N700), .A2(N614) );
  AND2_X1 AND2_137( .ZN(N1174), .A1(N700), .A2(N614) );
  BUF_X1 BUFF1_138( .Z(N1175), .A(N682) );
  BUF_X1 BUFF1_139( .Z(N1182), .A(N676) );
  INV_X1 NOT1_140( .ZN(N1189), .A(N657) );
  INV_X1 NOT1_141( .ZN(N1194), .A(N676) );
  INV_X1 NOT1_142( .ZN(N1199), .A(N682) );
  INV_X1 NOT1_143( .ZN(N1206), .A(N689) );
  BUF_X1 BUFF1_144( .Z(N1211), .A(N695) );
  INV_X1 NOT1_145( .ZN(N1218), .A(N750) );
  INV_X1 NOT1_146( .ZN(N1222), .A(N1028) );
  BUF_X1 BUFF1_147( .Z(N1227), .A(N632) );
  BUF_X1 BUFF1_148( .Z(N1233), .A(N676) );
  BUF_X1 BUFF1_149( .Z(N1240), .A(N632) );
  BUF_X1 BUFF1_150( .Z(N1244), .A(N676) );
  BUF_X1 BUFF1_151( .Z(N1249), .A(N689) );
  BUF_X1 BUFF1_152( .Z(N1256), .A(N689) );
  BUF_X1 BUFF1_153( .Z(N1263), .A(N695) );
  BUF_X1 BUFF1_154( .Z(N1270), .A(N689) );
  BUF_X1 BUFF1_155( .Z(N1277), .A(N689) );
  BUF_X1 BUFF1_156( .Z(N1284), .A(N700) );
  BUF_X1 BUFF1_157( .Z(N1287), .A(N614) );
  BUF_X1 BUFF1_158( .Z(N1290), .A(N666) );
  BUF_X1 BUFF1_159( .Z(N1293), .A(N660) );
  BUF_X1 BUFF1_160( .Z(N1296), .A(N651) );
  BUF_X1 BUFF1_161( .Z(N1299), .A(N614) );
  BUF_X1 BUFF1_162( .Z(N1302), .A(N644) );
  BUF_X1 BUFF1_163( .Z(N1305), .A(N700) );
  BUF_X1 BUFF1_164( .Z(N1308), .A(N614) );
  BUF_X1 BUFF1_165( .Z(N1311), .A(N614) );
  BUF_X1 BUFF1_166( .Z(N1314), .A(N666) );
  BUF_X1 BUFF1_167( .Z(N1317), .A(N660) );
  BUF_X1 BUFF1_168( .Z(N1320), .A(N651) );
  BUF_X1 BUFF1_169( .Z(N1323), .A(N644) );
  BUF_X1 BUFF1_170( .Z(N1326), .A(N609) );
  BUF_X1 BUFF1_171( .Z(N1329), .A(N604) );
  BUF_X1 BUFF1_172( .Z(N1332), .A(N742) );
  BUF_X1 BUFF1_173( .Z(N1335), .A(N599) );
  BUF_X1 BUFF1_174( .Z(N1338), .A(N727) );
  BUF_X1 BUFF1_175( .Z(N1341), .A(N721) );
  BUF_X1 BUFF1_176( .Z(N1344), .A(N715) );
  BUF_X1 BUFF1_177( .Z(N1347), .A(N734) );
  BUF_X1 BUFF1_178( .Z(N1350), .A(N708) );
  BUF_X1 BUFF1_179( .Z(N1353), .A(N609) );
  BUF_X1 BUFF1_180( .Z(N1356), .A(N604) );
  BUF_X1 BUFF1_181( .Z(N1359), .A(N742) );
  BUF_X1 BUFF1_182( .Z(N1362), .A(N734) );
  BUF_X1 BUFF1_183( .Z(N1365), .A(N599) );
  BUF_X1 BUFF1_184( .Z(N1368), .A(N727) );
  BUF_X1 BUFF1_185( .Z(N1371), .A(N721) );
  BUF_X1 BUFF1_186( .Z(N1374), .A(N715) );
  BUF_X1 BUFF1_187( .Z(N1377), .A(N708) );
  BUF_X1 BUFF1_188( .Z(N1380), .A(N806) );
  BUF_X1 BUFF1_189( .Z(N1383), .A(N800) );
  BUF_X1 BUFF1_190( .Z(N1386), .A(N794) );
  BUF_X1 BUFF1_191( .Z(N1389), .A(N786) );
  BUF_X1 BUFF1_192( .Z(N1392), .A(N780) );
  BUF_X1 BUFF1_193( .Z(N1395), .A(N774) );
  BUF_X1 BUFF1_194( .Z(N1398), .A(N768) );
  BUF_X1 BUFF1_195( .Z(N1401), .A(N762) );
  BUF_X1 BUFF1_196( .Z(N1404), .A(N806) );
  BUF_X1 BUFF1_197( .Z(N1407), .A(N800) );
  BUF_X1 BUFF1_198( .Z(N1410), .A(N794) );
  BUF_X1 BUFF1_199( .Z(N1413), .A(N780) );
  BUF_X1 BUFF1_200( .Z(N1416), .A(N774) );
  BUF_X1 BUFF1_201( .Z(N1419), .A(N768) );
  BUF_X1 BUFF1_202( .Z(N1422), .A(N762) );
  BUF_X1 BUFF1_203( .Z(N1425), .A(N786) );
  BUF_X1 BUFF1_204( .Z(N1428), .A(N636) );
  BUF_X1 BUFF1_205( .Z(N1431), .A(N636) );
  BUF_X1 BUFF1_206( .Z(N1434), .A(N865) );
  BUF_X1 BUFF1_207( .Z(N1437), .A(N859) );
  BUF_X1 BUFF1_208( .Z(N1440), .A(N853) );
  BUF_X1 BUFF1_209( .Z(N1443), .A(N845) );
  BUF_X1 BUFF1_210( .Z(N1446), .A(N839) );
  BUF_X1 BUFF1_211( .Z(N1449), .A(N833) );
  BUF_X1 BUFF1_212( .Z(N1452), .A(N827) );
  BUF_X1 BUFF1_213( .Z(N1455), .A(N821) );
  BUF_X1 BUFF1_214( .Z(N1458), .A(N814) );
  BUF_X2 BUFF1_215( .Z(N1461), .A(N865) );
  BUF_X2 BUFF1_216( .Z(N1464), .A(N859) );
  BUF_X2 BUFF1_217( .Z(N1467), .A(N853) );
  BUF_X4 BUFF1_218( .Z(N1470), .A(N839) );
  BUF_X4 BUFF1_219( .Z(N1473), .A(N833) );
  BUF_X1 BUFF1_220( .Z(N1476), .A(N827) );
  BUF_X1 BUFF1_221( .Z(N1479), .A(N821) );
  BUF_X1 BUFF1_222( .Z(N1482), .A(N845) );
  BUF_X1 BUFF1_223( .Z(N1485), .A(N814) );
  INV_X2 NOT1_224( .ZN(N1489), .A(N1109) );
  BUF_X1 BUFF1_225( .Z(N1490), .A(N1116) );
  AND2_X1 AND2_226( .ZN(N1537), .A1(N957), .A2(N614) );
  AND2_X1 AND2_227( .ZN(N1551), .A1(N614), .A2(N957) );
  AND2_X1 AND2_228( .ZN(N1649), .A1(N1029), .A2(N636) );
  BUF_X1 BUFF1_229( .Z(N1703), .A(N957) );
  NOR2_X1 NOR2_230( .ZN(N1708), .A1(N957), .A2(N614) );
  BUF_X1 BUFF1_231( .Z(N1713), .A(N957) );
  NOR2_X1 NOR2_232( .ZN(N1721), .A1(N614), .A2(N957) );
  BUF_X1 BUFF1_233( .Z(N1758), .A(N1029) );
  AND2_X1 AND2_234( .ZN(N1781), .A1(N163), .A2(N1116) );
  AND2_X1 AND2_235( .ZN(N1782), .A1(N170), .A2(N1125) );
  INV_X2 NOT1_236( .ZN(N1783), .A(N1125) );
  INV_X1 NOT1_237( .ZN(N1789), .A(N1136) );
  AND2_X1 AND2_238( .ZN(N1793), .A1(N169), .A2(N1125) );
  AND2_X1 AND2_239( .ZN(N1794), .A1(N168), .A2(N1125) );
  AND2_X1 AND2_240( .ZN(N1795), .A1(N167), .A2(N1125) );
  AND2_X1 AND2_241( .ZN(N1796), .A1(N166), .A2(N1136) );
  AND2_X1 AND2_242( .ZN(N1797), .A1(N165), .A2(N1136) );
  AND2_X1 AND2_243( .ZN(N1798), .A1(N164), .A2(N1136) );
  INV_X1 NOT1_244( .ZN(N1799), .A(N1147) );
  INV_X1 NOT1_245( .ZN(N1805), .A(N1160) );
  AND2_X1 AND2_246( .ZN(N1811), .A1(N177), .A2(N1147) );
  AND2_X1 AND2_247( .ZN(N1812), .A1(N176), .A2(N1147) );
  AND2_X1 AND2_248( .ZN(N1813), .A1(N175), .A2(N1147) );
  AND2_X1 AND2_249( .ZN(N1814), .A1(N174), .A2(N1147) );
  AND2_X1 AND2_250( .ZN(N1815), .A1(N173), .A2(N1147) );
  AND2_X1 AND2_251( .ZN(N1816), .A1(N157), .A2(N1160) );
  AND2_X1 AND2_252( .ZN(N1817), .A1(N156), .A2(N1160) );
  AND2_X1 AND2_253( .ZN(N1818), .A1(N155), .A2(N1160) );
  AND2_X1 AND2_254( .ZN(N1819), .A1(N154), .A2(N1160) );
  AND2_X1 AND2_255( .ZN(N1820), .A1(N153), .A2(N1160) );
  INV_X1 NOT1_256( .ZN(N1821), .A(N1284) );
  INV_X1 NOT1_257( .ZN(N1822), .A(N1287) );
  INV_X1 NOT1_258( .ZN(N1828), .A(N1290) );
  INV_X1 NOT1_259( .ZN(N1829), .A(N1293) );
  INV_X1 NOT1_260( .ZN(N1830), .A(N1296) );
  INV_X1 NOT1_261( .ZN(N1832), .A(N1299) );
  INV_X1 NOT1_262( .ZN(N1833), .A(N1302) );
  INV_X1 NOT1_263( .ZN(N1834), .A(N1305) );
  INV_X1 NOT1_264( .ZN(N1835), .A(N1308) );
  INV_X1 NOT1_265( .ZN(N1839), .A(N1311) );
  INV_X1 NOT1_266( .ZN(N1840), .A(N1314) );
  INV_X1 NOT1_267( .ZN(N1841), .A(N1317) );
  INV_X1 NOT1_268( .ZN(N1842), .A(N1320) );
  INV_X1 NOT1_269( .ZN(N1843), .A(N1323) );
  INV_X1 NOT1_270( .ZN(N1845), .A(N1175) );
  INV_X1 NOT1_271( .ZN(N1851), .A(N1182) );
  AND2_X1 AND2_272( .ZN(N1857), .A1(N181), .A2(N1175) );
  AND2_X1 AND2_273( .ZN(N1858), .A1(N171), .A2(N1175) );
  AND2_X1 AND2_274( .ZN(N1859), .A1(N180), .A2(N1175) );
  AND2_X1 AND2_275( .ZN(N1860), .A1(N179), .A2(N1175) );
  AND2_X1 AND2_276( .ZN(N1861), .A1(N178), .A2(N1175) );
  AND2_X1 AND2_277( .ZN(N1862), .A1(N161), .A2(N1182) );
  AND2_X1 AND2_278( .ZN(N1863), .A1(N151), .A2(N1182) );
  AND2_X1 AND2_279( .ZN(N1864), .A1(N160), .A2(N1182) );
  AND2_X1 AND2_280( .ZN(N1865), .A1(N159), .A2(N1182) );
  AND2_X1 AND2_281( .ZN(N1866), .A1(N158), .A2(N1182) );
  INV_X1 NOT1_282( .ZN(N1867), .A(N1326) );
  INV_X1 NOT1_283( .ZN(N1868), .A(N1329) );
  INV_X1 NOT1_284( .ZN(N1869), .A(N1332) );
  INV_X1 NOT1_285( .ZN(N1870), .A(N1335) );
  INV_X1 NOT1_286( .ZN(N1871), .A(N1338) );
  INV_X1 NOT1_287( .ZN(N1872), .A(N1341) );
  INV_X1 NOT1_288( .ZN(N1873), .A(N1344) );
  INV_X1 NOT1_289( .ZN(N1874), .A(N1347) );
  INV_X1 NOT1_290( .ZN(N1875), .A(N1350) );
  INV_X1 NOT1_291( .ZN(N1876), .A(N1353) );
  INV_X1 NOT1_292( .ZN(N1877), .A(N1356) );
  INV_X1 NOT1_293( .ZN(N1878), .A(N1359) );
  INV_X1 NOT1_294( .ZN(N1879), .A(N1362) );
  INV_X1 NOT1_295( .ZN(N1880), .A(N1365) );
  INV_X1 NOT1_296( .ZN(N1881), .A(N1368) );
  INV_X1 NOT1_297( .ZN(N1882), .A(N1371) );
  INV_X1 NOT1_298( .ZN(N1883), .A(N1374) );
  INV_X1 NOT1_299( .ZN(N1884), .A(N1377) );
  BUF_X1 BUFF1_300( .Z(N1885), .A(N1199) );
  BUF_X1 BUFF1_301( .Z(N1892), .A(N1194) );
  BUF_X1 BUFF1_302( .Z(N1899), .A(N1199) );
  BUF_X1 BUFF1_303( .Z(N1906), .A(N1194) );
  INV_X1 NOT1_304( .ZN(N1913), .A(N1211) );
  BUF_X1 BUFF1_305( .Z(N1919), .A(N1194) );
  AND2_X1 AND2_306( .ZN(N1926), .A1(N44), .A2(N1211) );
  AND2_X1 AND2_307( .ZN(N1927), .A1(N41), .A2(N1211) );
  AND2_X1 AND2_308( .ZN(N1928), .A1(N29), .A2(N1211) );
  AND2_X1 AND2_309( .ZN(N1929), .A1(N26), .A2(N1211) );
  AND2_X1 AND2_310( .ZN(N1930), .A1(N23), .A2(N1211) );
  INV_X1 NOT1_311( .ZN(N1931), .A(N1380) );
  INV_X1 NOT1_312( .ZN(N1932), .A(N1383) );
  INV_X1 NOT1_313( .ZN(N1933), .A(N1386) );
  INV_X2 NOT1_314( .ZN(N1934), .A(N1389) );
  INV_X2 NOT1_315( .ZN(N1935), .A(N1392) );
  INV_X2 NOT1_316( .ZN(N1936), .A(N1395) );
  INV_X2 NOT1_317( .ZN(N1937), .A(N1398) );
  INV_X2 NOT1_318( .ZN(N1938), .A(N1401) );
  INV_X2 NOT1_319( .ZN(N1939), .A(N1404) );
  INV_X2 NOT1_320( .ZN(N1940), .A(N1407) );
  INV_X1 NOT1_321( .ZN(N1941), .A(N1410) );
  INV_X1 NOT1_322( .ZN(N1942), .A(N1413) );
  INV_X1 NOT1_323( .ZN(N1943), .A(N1416) );
  INV_X1 NOT1_324( .ZN(N1944), .A(N1419) );
  INV_X1 NOT1_325( .ZN(N1945), .A(N1422) );
  INV_X1 NOT1_326( .ZN(N1946), .A(N1425) );
  INV_X1 NOT1_327( .ZN(N1947), .A(N1233) );
  INV_X1 NOT1_328( .ZN(N1953), .A(N1244) );
  AND2_X1 AND2_329( .ZN(N1957), .A1(N209), .A2(N1233) );
  AND2_X1 AND2_330( .ZN(N1958), .A1(N216), .A2(N1233) );
  AND2_X1 AND2_331( .ZN(N1959), .A1(N215), .A2(N1233) );
  AND2_X1 AND2_332( .ZN(N1960), .A1(N214), .A2(N1233) );
  AND2_X1 AND2_333( .ZN(N1961), .A1(N213), .A2(N1244) );
  AND2_X1 AND2_334( .ZN(N1962), .A1(N212), .A2(N1244) );
  AND2_X1 AND2_335( .ZN(N1963), .A1(N211), .A2(N1244) );
  INV_X1 NOT1_336( .ZN(N1965), .A(N1428) );
  AND2_X1 AND2_337( .ZN(N1966), .A1(N1222), .A2(N636) );
  INV_X1 NOT1_338( .ZN(N1967), .A(N1431) );
  INV_X1 NOT1_339( .ZN(N1968), .A(N1434) );
  INV_X1 NOT1_340( .ZN(N1969), .A(N1437) );
  INV_X1 NOT1_341( .ZN(N1970), .A(N1440) );
  INV_X1 NOT1_342( .ZN(N1971), .A(N1443) );
  INV_X1 NOT1_343( .ZN(N1972), .A(N1446) );
  INV_X1 NOT1_344( .ZN(N1973), .A(N1449) );
  INV_X1 NOT1_345( .ZN(N1974), .A(N1452) );
  INV_X1 NOT1_346( .ZN(N1975), .A(N1455) );
  INV_X1 NOT1_347( .ZN(N1976), .A(N1458) );
  INV_X1 NOT1_348( .ZN(N1977), .A(N1249) );
  INV_X1 NOT1_349( .ZN(N1983), .A(N1256) );
  AND2_X1 AND2_350( .ZN(N1989), .A1(N642), .A2(N1249) );
  AND2_X1 AND2_351( .ZN(N1990), .A1(N644), .A2(N1249) );
  AND2_X1 AND2_352( .ZN(N1991), .A1(N651), .A2(N1249) );
  AND2_X1 AND2_353( .ZN(N1992), .A1(N674), .A2(N1249) );
  AND2_X1 AND2_354( .ZN(N1993), .A1(N660), .A2(N1249) );
  AND2_X1 AND2_355( .ZN(N1994), .A1(N666), .A2(N1256) );
  AND2_X1 AND2_356( .ZN(N1995), .A1(N672), .A2(N1256) );
  AND2_X1 AND2_357( .ZN(N1996), .A1(N673), .A2(N1256) );
  INV_X1 NOT1_358( .ZN(N1997), .A(N1263) );
  BUF_X4 BUFF1_359( .Z(N2003), .A(N1194) );
  AND2_X1 AND2_360( .ZN(N2010), .A1(N47), .A2(N1263) );
  AND2_X1 AND2_361( .ZN(N2011), .A1(N35), .A2(N1263) );
  AND2_X1 AND2_362( .ZN(N2012), .A1(N32), .A2(N1263) );
  AND2_X1 AND2_363( .ZN(N2013), .A1(N50), .A2(N1263) );
  AND2_X1 AND2_364( .ZN(N2014), .A1(N66), .A2(N1263) );
  INV_X1 NOT1_365( .ZN(N2015), .A(N1461) );
  INV_X1 NOT1_366( .ZN(N2016), .A(N1464) );
  INV_X1 NOT1_367( .ZN(N2017), .A(N1467) );
  INV_X1 NOT1_368( .ZN(N2018), .A(N1470) );
  INV_X1 NOT1_369( .ZN(N2019), .A(N1473) );
  INV_X1 NOT1_370( .ZN(N2020), .A(N1476) );
  INV_X1 NOT1_371( .ZN(N2021), .A(N1479) );
  INV_X1 NOT1_372( .ZN(N2022), .A(N1482) );
  INV_X1 NOT1_373( .ZN(N2023), .A(N1485) );
  BUF_X1 BUFF1_374( .Z(N2024), .A(N1206) );
  BUF_X1 BUFF1_375( .Z(N2031), .A(N1206) );
  BUF_X1 BUFF1_376( .Z(N2038), .A(N1206) );
  BUF_X1 BUFF1_377( .Z(N2045), .A(N1206) );
  INV_X1 NOT1_378( .ZN(N2052), .A(N1270) );
  INV_X1 NOT1_379( .ZN(N2058), .A(N1277) );
  AND2_X1 AND2_380( .ZN(N2064), .A1(N706), .A2(N1270) );
  AND2_X1 AND2_381( .ZN(N2065), .A1(N708), .A2(N1270) );
  AND2_X1 AND2_382( .ZN(N2066), .A1(N715), .A2(N1270) );
  AND2_X1 AND2_383( .ZN(N2067), .A1(N721), .A2(N1270) );
  AND2_X1 AND2_384( .ZN(N2068), .A1(N727), .A2(N1270) );
  AND2_X1 AND2_385( .ZN(N2069), .A1(N733), .A2(N1277) );
  AND2_X1 AND2_386( .ZN(N2070), .A1(N734), .A2(N1277) );
  AND2_X1 AND2_387( .ZN(N2071), .A1(N742), .A2(N1277) );
  AND2_X1 AND2_388( .ZN(N2072), .A1(N748), .A2(N1277) );
  AND2_X1 AND2_389( .ZN(N2073), .A1(N749), .A2(N1277) );
  BUF_X1 BUFF1_390( .Z(N2074), .A(N1189) );
  BUF_X1 BUFF1_391( .Z(N2081), .A(N1189) );
  BUF_X1 BUFF1_392( .Z(N2086), .A(N1222) );
  NAND2_X2 NAND2_393( .ZN(N2107), .A1(N1287), .A2(N1821) );
  NAND2_X1 NAND2_394( .ZN(N2108), .A1(N1284), .A2(N1822) );
  INV_X1 NOT1_395( .ZN(N2110), .A(N1703) );
  NAND2_X1 NAND2_396( .ZN(N2111), .A1(N1703), .A2(N1832) );
  NAND2_X1 NAND2_397( .ZN(N2112), .A1(N1308), .A2(N1834) );
  NAND2_X1 NAND2_398( .ZN(N2113), .A1(N1305), .A2(N1835) );
  INV_X1 NOT1_399( .ZN(N2114), .A(N1713) );
  NAND2_X1 NAND2_400( .ZN(N2115), .A1(N1713), .A2(N1839) );
  INV_X1 NOT1_401( .ZN(N2117), .A(N1721) );
  INV_X1 NOT1_402( .ZN(N2171), .A(N1758) );
  NAND2_X1 NAND2_403( .ZN(N2172), .A1(N1758), .A2(N1965) );
  INV_X1 NOT1_404( .ZN(N2230), .A(N1708) );
  BUF_X1 BUFF1_405( .Z(N2231), .A(N1537) );
  BUF_X1 BUFF1_406( .Z(N2235), .A(N1551) );
  OR2_X1 OR2_407( .ZN(N2239), .A1(N1783), .A2(N1782) );
  OR2_X1 OR2_408( .ZN(N2240), .A1(N1783), .A2(N1125) );
  OR2_X1 OR2_409( .ZN(N2241), .A1(N1783), .A2(N1793) );
  OR2_X1 OR2_410( .ZN(N2242), .A1(N1783), .A2(N1794) );
  OR2_X1 OR2_411( .ZN(N2243), .A1(N1783), .A2(N1795) );
  OR2_X2 OR2_412( .ZN(N2244), .A1(N1789), .A2(N1796) );
  OR2_X2 OR2_413( .ZN(N2245), .A1(N1789), .A2(N1797) );
  OR2_X2 OR2_414( .ZN(N2246), .A1(N1789), .A2(N1798) );
  OR2_X2 OR2_415( .ZN(N2247), .A1(N1799), .A2(N1811) );
  OR2_X2 OR2_416( .ZN(N2248), .A1(N1799), .A2(N1812) );
  OR2_X1 OR2_417( .ZN(N2249), .A1(N1799), .A2(N1813) );
  OR2_X1 OR2_418( .ZN(N2250), .A1(N1799), .A2(N1814) );
  OR2_X1 OR2_419( .ZN(N2251), .A1(N1799), .A2(N1815) );
  OR2_X1 OR2_420( .ZN(N2252), .A1(N1805), .A2(N1816) );
  OR2_X1 OR2_421( .ZN(N2253), .A1(N1805), .A2(N1817) );
  OR2_X1 OR2_422( .ZN(N2254), .A1(N1805), .A2(N1818) );
  OR2_X1 OR2_423( .ZN(N2255), .A1(N1805), .A2(N1819) );
  OR2_X1 OR2_424( .ZN(N2256), .A1(N1805), .A2(N1820) );
  NAND2_X1 NAND2_425( .ZN(N2257), .A1(N2107), .A2(N2108) );
  INV_X1 NOT1_426( .ZN(N2267), .A(N2074) );
  NAND2_X1 NAND2_427( .ZN(N2268), .A1(N1299), .A2(N2110) );
  NAND2_X1 NAND2_428( .ZN(N2269), .A1(N2112), .A2(N2113) );
  NAND2_X1 NAND2_429( .ZN(N2274), .A1(N1311), .A2(N2114) );
  INV_X1 NOT1_430( .ZN(N2275), .A(N2081) );
  AND2_X1 AND2_431( .ZN(N2277), .A1(N141), .A2(N1845) );
  AND2_X1 AND2_432( .ZN(N2278), .A1(N147), .A2(N1845) );
  AND2_X1 AND2_433( .ZN(N2279), .A1(N138), .A2(N1845) );
  AND2_X1 AND2_434( .ZN(N2280), .A1(N144), .A2(N1845) );
  AND2_X1 AND2_435( .ZN(N2281), .A1(N135), .A2(N1845) );
  AND2_X1 AND2_436( .ZN(N2282), .A1(N141), .A2(N1851) );
  AND2_X1 AND2_437( .ZN(N2283), .A1(N147), .A2(N1851) );
  AND2_X1 AND2_438( .ZN(N2284), .A1(N138), .A2(N1851) );
  AND2_X1 AND2_439( .ZN(N2285), .A1(N144), .A2(N1851) );
  AND2_X1 AND2_440( .ZN(N2286), .A1(N135), .A2(N1851) );
  INV_X1 NOT1_441( .ZN(N2287), .A(N1885) );
  INV_X1 NOT1_442( .ZN(N2293), .A(N1892) );
  AND2_X1 AND2_443( .ZN(N2299), .A1(N103), .A2(N1885) );
  AND2_X1 AND2_444( .ZN(N2300), .A1(N130), .A2(N1885) );
  AND2_X1 AND2_445( .ZN(N2301), .A1(N127), .A2(N1885) );
  AND2_X1 AND2_446( .ZN(N2302), .A1(N124), .A2(N1885) );
  AND2_X1 AND2_447( .ZN(N2303), .A1(N100), .A2(N1885) );
  AND2_X1 AND2_448( .ZN(N2304), .A1(N103), .A2(N1892) );
  AND2_X1 AND2_449( .ZN(N2305), .A1(N130), .A2(N1892) );
  AND2_X1 AND2_450( .ZN(N2306), .A1(N127), .A2(N1892) );
  AND2_X1 AND2_451( .ZN(N2307), .A1(N124), .A2(N1892) );
  AND2_X1 AND2_452( .ZN(N2308), .A1(N100), .A2(N1892) );
  INV_X1 NOT1_453( .ZN(N2309), .A(N1899) );
  INV_X1 NOT1_454( .ZN(N2315), .A(N1906) );
  AND2_X1 AND2_455( .ZN(N2321), .A1(N115), .A2(N1899) );
  AND2_X1 AND2_456( .ZN(N2322), .A1(N118), .A2(N1899) );
  AND2_X1 AND2_457( .ZN(N2323), .A1(N97), .A2(N1899) );
  AND2_X1 AND2_458( .ZN(N2324), .A1(N94), .A2(N1899) );
  AND2_X1 AND2_459( .ZN(N2325), .A1(N121), .A2(N1899) );
  AND2_X1 AND2_460( .ZN(N2326), .A1(N115), .A2(N1906) );
  AND2_X1 AND2_461( .ZN(N2327), .A1(N118), .A2(N1906) );
  AND2_X1 AND2_462( .ZN(N2328), .A1(N97), .A2(N1906) );
  AND2_X1 AND2_463( .ZN(N2329), .A1(N94), .A2(N1906) );
  AND2_X1 AND2_464( .ZN(N2330), .A1(N121), .A2(N1906) );
  INV_X2 NOT1_465( .ZN(N2331), .A(N1919) );
  AND2_X1 AND2_466( .ZN(N2337), .A1(N208), .A2(N1913) );
  AND2_X1 AND2_467( .ZN(N2338), .A1(N198), .A2(N1913) );
  AND2_X1 AND2_468( .ZN(N2339), .A1(N207), .A2(N1913) );
  AND2_X1 AND2_469( .ZN(N2340), .A1(N206), .A2(N1913) );
  AND2_X1 AND2_470( .ZN(N2341), .A1(N205), .A2(N1913) );
  AND2_X1 AND2_471( .ZN(N2342), .A1(N44), .A2(N1919) );
  AND2_X1 AND2_472( .ZN(N2343), .A1(N41), .A2(N1919) );
  AND2_X1 AND2_473( .ZN(N2344), .A1(N29), .A2(N1919) );
  AND2_X1 AND2_474( .ZN(N2345), .A1(N26), .A2(N1919) );
  AND2_X1 AND2_475( .ZN(N2346), .A1(N23), .A2(N1919) );
  OR2_X1 OR2_476( .ZN(N2347), .A1(N1947), .A2(N1233) );
  OR2_X1 OR2_477( .ZN(N2348), .A1(N1947), .A2(N1957) );
  OR2_X1 OR2_478( .ZN(N2349), .A1(N1947), .A2(N1958) );
  OR2_X1 OR2_479( .ZN(N2350), .A1(N1947), .A2(N1959) );
  OR2_X1 OR2_480( .ZN(N2351), .A1(N1947), .A2(N1960) );
  OR2_X1 OR2_481( .ZN(N2352), .A1(N1953), .A2(N1961) );
  OR2_X1 OR2_482( .ZN(N2353), .A1(N1953), .A2(N1962) );
  OR2_X1 OR2_483( .ZN(N2354), .A1(N1953), .A2(N1963) );
  NAND2_X1 NAND2_484( .ZN(N2355), .A1(N1428), .A2(N2171) );
  INV_X2 NOT1_485( .ZN(N2356), .A(N2086) );
  NAND2_X1 NAND2_486( .ZN(N2357), .A1(N2086), .A2(N1967) );
  AND2_X1 AND2_487( .ZN(N2358), .A1(N114), .A2(N1977) );
  AND2_X1 AND2_488( .ZN(N2359), .A1(N113), .A2(N1977) );
  AND2_X1 AND2_489( .ZN(N2360), .A1(N111), .A2(N1977) );
  AND2_X1 AND2_490( .ZN(N2361), .A1(N87), .A2(N1977) );
  AND2_X1 AND2_491( .ZN(N2362), .A1(N112), .A2(N1977) );
  AND2_X1 AND2_492( .ZN(N2363), .A1(N88), .A2(N1983) );
  AND2_X1 AND2_493( .ZN(N2364), .A1(N245), .A2(N1983) );
  AND2_X1 AND2_494( .ZN(N2365), .A1(N271), .A2(N1983) );
  AND2_X1 AND2_495( .ZN(N2366), .A1(N759), .A2(N1983) );
  AND2_X1 AND2_496( .ZN(N2367), .A1(N70), .A2(N1983) );
  INV_X1 NOT1_497( .ZN(N2368), .A(N2003) );
  AND2_X1 AND2_498( .ZN(N2374), .A1(N193), .A2(N1997) );
  AND2_X1 AND2_499( .ZN(N2375), .A1(N192), .A2(N1997) );
  AND2_X1 AND2_500( .ZN(N2376), .A1(N191), .A2(N1997) );
  AND2_X1 AND2_501( .ZN(N2377), .A1(N190), .A2(N1997) );
  AND2_X1 AND2_502( .ZN(N2378), .A1(N189), .A2(N1997) );
  AND2_X1 AND2_503( .ZN(N2379), .A1(N47), .A2(N2003) );
  AND2_X1 AND2_504( .ZN(N2380), .A1(N35), .A2(N2003) );
  AND2_X1 AND2_505( .ZN(N2381), .A1(N32), .A2(N2003) );
  AND2_X1 AND2_506( .ZN(N2382), .A1(N50), .A2(N2003) );
  AND2_X1 AND2_507( .ZN(N2383), .A1(N66), .A2(N2003) );
  INV_X1 NOT1_508( .ZN(N2384), .A(N2024) );
  INV_X1 NOT1_509( .ZN(N2390), .A(N2031) );
  AND2_X1 AND2_510( .ZN(N2396), .A1(N58), .A2(N2024) );
  AND2_X1 AND2_511( .ZN(N2397), .A1(N77), .A2(N2024) );
  AND2_X1 AND2_512( .ZN(N2398), .A1(N78), .A2(N2024) );
  AND2_X1 AND2_513( .ZN(N2399), .A1(N59), .A2(N2024) );
  AND2_X1 AND2_514( .ZN(N2400), .A1(N81), .A2(N2024) );
  AND2_X1 AND2_515( .ZN(N2401), .A1(N80), .A2(N2031) );
  AND2_X1 AND2_516( .ZN(N2402), .A1(N79), .A2(N2031) );
  AND2_X1 AND2_517( .ZN(N2403), .A1(N60), .A2(N2031) );
  AND2_X1 AND2_518( .ZN(N2404), .A1(N61), .A2(N2031) );
  AND2_X1 AND2_519( .ZN(N2405), .A1(N62), .A2(N2031) );
  INV_X1 NOT1_520( .ZN(N2406), .A(N2038) );
  INV_X1 NOT1_521( .ZN(N2412), .A(N2045) );
  AND2_X1 AND2_522( .ZN(N2418), .A1(N69), .A2(N2038) );
  AND2_X1 AND2_523( .ZN(N2419), .A1(N70), .A2(N2038) );
  AND2_X1 AND2_524( .ZN(N2420), .A1(N74), .A2(N2038) );
  AND2_X1 AND2_525( .ZN(N2421), .A1(N76), .A2(N2038) );
  AND2_X1 AND2_526( .ZN(N2422), .A1(N75), .A2(N2038) );
  AND2_X1 AND2_527( .ZN(N2423), .A1(N73), .A2(N2045) );
  AND2_X1 AND2_528( .ZN(N2424), .A1(N53), .A2(N2045) );
  AND2_X1 AND2_529( .ZN(N2425), .A1(N54), .A2(N2045) );
  AND2_X1 AND2_530( .ZN(N2426), .A1(N55), .A2(N2045) );
  AND2_X2 AND2_531( .ZN(N2427), .A1(N56), .A2(N2045) );
  AND2_X2 AND2_532( .ZN(N2428), .A1(N82), .A2(N2052) );
  AND2_X2 AND2_533( .ZN(N2429), .A1(N65), .A2(N2052) );
  AND2_X2 AND2_534( .ZN(N2430), .A1(N83), .A2(N2052) );
  AND2_X1 AND2_535( .ZN(N2431), .A1(N84), .A2(N2052) );
  AND2_X1 AND2_536( .ZN(N2432), .A1(N85), .A2(N2052) );
  AND2_X1 AND2_537( .ZN(N2433), .A1(N64), .A2(N2058) );
  AND2_X1 AND2_538( .ZN(N2434), .A1(N63), .A2(N2058) );
  AND2_X1 AND2_539( .ZN(N2435), .A1(N86), .A2(N2058) );
  AND2_X1 AND2_540( .ZN(N2436), .A1(N109), .A2(N2058) );
  AND2_X1 AND2_541( .ZN(N2437), .A1(N110), .A2(N2058) );
  AND2_X1 AND2_542( .ZN(N2441), .A1(N2239), .A2(N1119) );
  AND2_X1 AND2_543( .ZN(N2442), .A1(N2240), .A2(N1119) );
  AND2_X1 AND2_544( .ZN(N2446), .A1(N2241), .A2(N1119) );
  AND2_X1 AND2_545( .ZN(N2450), .A1(N2242), .A2(N1119) );
  AND2_X1 AND2_546( .ZN(N2454), .A1(N2243), .A2(N1119) );
  AND2_X1 AND2_547( .ZN(N2458), .A1(N2244), .A2(N1132) );
  AND2_X1 AND2_548( .ZN(N2462), .A1(N2247), .A2(N1141) );
  AND2_X1 AND2_549( .ZN(N2466), .A1(N2248), .A2(N1141) );
  AND2_X1 AND2_550( .ZN(N2470), .A1(N2249), .A2(N1141) );
  AND2_X1 AND2_551( .ZN(N2474), .A1(N2250), .A2(N1141) );
  AND2_X1 AND2_552( .ZN(N2478), .A1(N2251), .A2(N1141) );
  AND2_X1 AND2_553( .ZN(N2482), .A1(N2252), .A2(N1154) );
  AND2_X1 AND2_554( .ZN(N2488), .A1(N2253), .A2(N1154) );
  AND2_X1 AND2_555( .ZN(N2496), .A1(N2254), .A2(N1154) );
  AND2_X1 AND2_556( .ZN(N2502), .A1(N2255), .A2(N1154) );
  AND2_X1 AND2_557( .ZN(N2508), .A1(N2256), .A2(N1154) );
  NAND2_X2 NAND2_558( .ZN(N2523), .A1(N2268), .A2(N2111) );
  NAND2_X1 NAND2_559( .ZN(N2533), .A1(N2274), .A2(N2115) );
  INV_X1 NOT1_560( .ZN(N2537), .A(N2235) );
  OR2_X1 OR2_561( .ZN(N2538), .A1(N2278), .A2(N1858) );
  OR2_X1 OR2_562( .ZN(N2542), .A1(N2279), .A2(N1859) );
  OR2_X1 OR2_563( .ZN(N2546), .A1(N2280), .A2(N1860) );
  OR2_X1 OR2_564( .ZN(N2550), .A1(N2281), .A2(N1861) );
  OR2_X1 OR2_565( .ZN(N2554), .A1(N2283), .A2(N1863) );
  OR2_X1 OR2_566( .ZN(N2561), .A1(N2284), .A2(N1864) );
  OR2_X1 OR2_567( .ZN(N2567), .A1(N2285), .A2(N1865) );
  OR2_X1 OR2_568( .ZN(N2573), .A1(N2286), .A2(N1866) );
  OR2_X1 OR2_569( .ZN(N2604), .A1(N2338), .A2(N1927) );
  OR2_X1 OR2_570( .ZN(N2607), .A1(N2339), .A2(N1928) );
  OR2_X1 OR2_571( .ZN(N2611), .A1(N2340), .A2(N1929) );
  OR2_X1 OR2_572( .ZN(N2615), .A1(N2341), .A2(N1930) );
  AND2_X1 AND2_573( .ZN(N2619), .A1(N2348), .A2(N1227) );
  AND2_X1 AND2_574( .ZN(N2626), .A1(N2349), .A2(N1227) );
  AND2_X1 AND2_575( .ZN(N2632), .A1(N2350), .A2(N1227) );
  AND2_X1 AND2_576( .ZN(N2638), .A1(N2351), .A2(N1227) );
  AND2_X1 AND2_577( .ZN(N2644), .A1(N2352), .A2(N1240) );
  NAND2_X1 NAND2_578( .ZN(N2650), .A1(N2355), .A2(N2172) );
  NAND2_X1 NAND2_579( .ZN(N2653), .A1(N1431), .A2(N2356) );
  OR2_X1 OR2_580( .ZN(N2654), .A1(N2359), .A2(N1990) );
  OR2_X1 OR2_581( .ZN(N2658), .A1(N2360), .A2(N1991) );
  OR2_X1 OR2_582( .ZN(N2662), .A1(N2361), .A2(N1992) );
  OR2_X1 OR2_583( .ZN(N2666), .A1(N2362), .A2(N1993) );
  OR2_X1 OR2_584( .ZN(N2670), .A1(N2363), .A2(N1994) );
  OR2_X1 OR2_585( .ZN(N2674), .A1(N2366), .A2(N1256) );
  OR2_X1 OR2_586( .ZN(N2680), .A1(N2367), .A2(N1256) );
  OR2_X1 OR2_587( .ZN(N2688), .A1(N2374), .A2(N2010) );
  OR2_X1 OR2_588( .ZN(N2692), .A1(N2375), .A2(N2011) );
  OR2_X1 OR2_589( .ZN(N2696), .A1(N2376), .A2(N2012) );
  OR2_X1 OR2_590( .ZN(N2700), .A1(N2377), .A2(N2013) );
  OR2_X1 OR2_591( .ZN(N2704), .A1(N2378), .A2(N2014) );
  AND2_X1 AND2_592( .ZN(N2728), .A1(N2347), .A2(N1227) );
  OR2_X1 OR2_593( .ZN(N2729), .A1(N2429), .A2(N2065) );
  OR2_X1 OR2_594( .ZN(N2733), .A1(N2430), .A2(N2066) );
  OR2_X1 OR2_595( .ZN(N2737), .A1(N2431), .A2(N2067) );
  OR2_X1 OR2_596( .ZN(N2741), .A1(N2432), .A2(N2068) );
  OR2_X1 OR2_597( .ZN(N2745), .A1(N2433), .A2(N2069) );
  OR2_X1 OR2_598( .ZN(N2749), .A1(N2434), .A2(N2070) );
  OR2_X1 OR2_599( .ZN(N2753), .A1(N2435), .A2(N2071) );
  OR2_X1 OR2_600( .ZN(N2757), .A1(N2436), .A2(N2072) );
  OR2_X1 OR2_601( .ZN(N2761), .A1(N2437), .A2(N2073) );
  INV_X2 NOT1_602( .ZN(N2765), .A(N2231) );
  AND2_X1 AND2_603( .ZN(N2766), .A1(N2354), .A2(N1240) );
  AND2_X1 AND2_604( .ZN(N2769), .A1(N2353), .A2(N1240) );
  AND2_X1 AND2_605( .ZN(N2772), .A1(N2246), .A2(N1132) );
  AND2_X1 AND2_606( .ZN(N2775), .A1(N2245), .A2(N1132) );
  OR2_X1 OR2_607( .ZN(N2778), .A1(N2282), .A2(N1862) );
  OR2_X1 OR2_608( .ZN(N2781), .A1(N2358), .A2(N1989) );
  OR2_X1 OR2_609( .ZN(N2784), .A1(N2365), .A2(N1996) );
  OR2_X1 OR2_610( .ZN(N2787), .A1(N2364), .A2(N1995) );
  OR2_X1 OR2_611( .ZN(N2790), .A1(N2337), .A2(N1926) );
  OR2_X1 OR2_612( .ZN(N2793), .A1(N2277), .A2(N1857) );
  OR2_X1 OR2_613( .ZN(N2796), .A1(N2428), .A2(N2064) );
  AND2_X1 AND2_614( .ZN(N2866), .A1(N2257), .A2(N1537) );
  AND2_X1 AND2_615( .ZN(N2867), .A1(N2257), .A2(N1537) );
  AND2_X1 AND2_616( .ZN(N2868), .A1(N2257), .A2(N1537) );
  AND2_X1 AND2_617( .ZN(N2869), .A1(N2257), .A2(N1537) );
  AND2_X1 AND2_618( .ZN(N2878), .A1(N2269), .A2(N1551) );
  AND2_X1 AND2_619( .ZN(N2913), .A1(N204), .A2(N2287) );
  AND2_X1 AND2_620( .ZN(N2914), .A1(N203), .A2(N2287) );
  AND2_X1 AND2_621( .ZN(N2915), .A1(N202), .A2(N2287) );
  AND2_X1 AND2_622( .ZN(N2916), .A1(N201), .A2(N2287) );
  AND2_X1 AND2_623( .ZN(N2917), .A1(N200), .A2(N2287) );
  AND2_X1 AND2_624( .ZN(N2918), .A1(N235), .A2(N2293) );
  AND2_X1 AND2_625( .ZN(N2919), .A1(N234), .A2(N2293) );
  AND2_X1 AND2_626( .ZN(N2920), .A1(N233), .A2(N2293) );
  AND2_X1 AND2_627( .ZN(N2921), .A1(N232), .A2(N2293) );
  AND2_X1 AND2_628( .ZN(N2922), .A1(N231), .A2(N2293) );
  AND2_X1 AND2_629( .ZN(N2923), .A1(N197), .A2(N2309) );
  AND2_X1 AND2_630( .ZN(N2924), .A1(N187), .A2(N2309) );
  AND2_X1 AND2_631( .ZN(N2925), .A1(N196), .A2(N2309) );
  AND2_X1 AND2_632( .ZN(N2926), .A1(N195), .A2(N2309) );
  AND2_X1 AND2_633( .ZN(N2927), .A1(N194), .A2(N2309) );
  AND2_X1 AND2_634( .ZN(N2928), .A1(N227), .A2(N2315) );
  AND2_X1 AND2_635( .ZN(N2929), .A1(N217), .A2(N2315) );
  AND2_X1 AND2_636( .ZN(N2930), .A1(N226), .A2(N2315) );
  AND2_X1 AND2_637( .ZN(N2931), .A1(N225), .A2(N2315) );
  AND2_X1 AND2_638( .ZN(N2932), .A1(N224), .A2(N2315) );
  AND2_X1 AND2_639( .ZN(N2933), .A1(N239), .A2(N2331) );
  AND2_X1 AND2_640( .ZN(N2934), .A1(N229), .A2(N2331) );
  AND2_X1 AND2_641( .ZN(N2935), .A1(N238), .A2(N2331) );
  AND2_X1 AND2_642( .ZN(N2936), .A1(N237), .A2(N2331) );
  AND2_X1 AND2_643( .ZN(N2937), .A1(N236), .A2(N2331) );
  NAND2_X1 NAND2_644( .ZN(N2988), .A1(N2653), .A2(N2357) );
  AND2_X1 AND2_645( .ZN(N3005), .A1(N223), .A2(N2368) );
  AND2_X1 AND2_646( .ZN(N3006), .A1(N222), .A2(N2368) );
  AND2_X1 AND2_647( .ZN(N3007), .A1(N221), .A2(N2368) );
  AND2_X1 AND2_648( .ZN(N3008), .A1(N220), .A2(N2368) );
  AND2_X1 AND2_649( .ZN(N3009), .A1(N219), .A2(N2368) );
  AND2_X1 AND2_650( .ZN(N3020), .A1(N812), .A2(N2384) );
  AND2_X1 AND2_651( .ZN(N3021), .A1(N814), .A2(N2384) );
  AND2_X1 AND2_652( .ZN(N3022), .A1(N821), .A2(N2384) );
  AND2_X1 AND2_653( .ZN(N3023), .A1(N827), .A2(N2384) );
  AND2_X1 AND2_654( .ZN(N3024), .A1(N833), .A2(N2384) );
  AND2_X1 AND2_655( .ZN(N3025), .A1(N839), .A2(N2390) );
  AND2_X1 AND2_656( .ZN(N3026), .A1(N845), .A2(N2390) );
  AND2_X1 AND2_657( .ZN(N3027), .A1(N853), .A2(N2390) );
  AND2_X1 AND2_658( .ZN(N3028), .A1(N859), .A2(N2390) );
  AND2_X1 AND2_659( .ZN(N3029), .A1(N865), .A2(N2390) );
  AND2_X1 AND2_660( .ZN(N3032), .A1(N758), .A2(N2406) );
  AND2_X1 AND2_661( .ZN(N3033), .A1(N759), .A2(N2406) );
  AND2_X1 AND2_662( .ZN(N3034), .A1(N762), .A2(N2406) );
  AND2_X1 AND2_663( .ZN(N3035), .A1(N768), .A2(N2406) );
  AND2_X1 AND2_664( .ZN(N3036), .A1(N774), .A2(N2406) );
  AND2_X1 AND2_665( .ZN(N3037), .A1(N780), .A2(N2412) );
  AND2_X1 AND2_666( .ZN(N3038), .A1(N786), .A2(N2412) );
  AND2_X1 AND2_667( .ZN(N3039), .A1(N794), .A2(N2412) );
  AND2_X1 AND2_668( .ZN(N3040), .A1(N800), .A2(N2412) );
  AND2_X1 AND2_669( .ZN(N3041), .A1(N806), .A2(N2412) );
  BUF_X4 BUFF1_670( .Z(N3061), .A(N2257) );
  BUF_X4 BUFF1_671( .Z(N3064), .A(N2257) );
  BUF_X1 BUFF1_672( .Z(N3067), .A(N2269) );
  BUF_X1 BUFF1_673( .Z(N3070), .A(N2269) );
  INV_X1 NOT1_674( .ZN(N3073), .A(N2728) );
  INV_X1 NOT1_675( .ZN(N3080), .A(N2441) );
  AND2_X1 AND2_676( .ZN(N3096), .A1(N666), .A2(N2644) );
  AND2_X1 AND2_677( .ZN(N3097), .A1(N660), .A2(N2638) );
  AND2_X1 AND2_678( .ZN(N3101), .A1(N1189), .A2(N2632) );
  AND2_X1 AND2_679( .ZN(N3107), .A1(N651), .A2(N2626) );
  AND2_X1 AND2_680( .ZN(N3114), .A1(N644), .A2(N2619) );
  AND2_X1 AND2_681( .ZN(N3122), .A1(N2523), .A2(N2257) );
  OR2_X1 OR2_682( .ZN(N3126), .A1(N1167), .A2(N2866) );
  AND2_X1 AND2_683( .ZN(N3130), .A1(N2523), .A2(N2257) );
  OR2_X1 OR2_684( .ZN(N3131), .A1(N1167), .A2(N2869) );
  AND2_X1 AND2_685( .ZN(N3134), .A1(N2523), .A2(N2257) );
  INV_X1 NOT1_686( .ZN(N3135), .A(N2533) );
  AND2_X1 AND2_687( .ZN(N3136), .A1(N666), .A2(N2644) );
  AND2_X1 AND2_688( .ZN(N3137), .A1(N660), .A2(N2638) );
  AND2_X1 AND2_689( .ZN(N3140), .A1(N1189), .A2(N2632) );
  AND2_X1 AND2_690( .ZN(N3144), .A1(N651), .A2(N2626) );
  AND2_X1 AND2_691( .ZN(N3149), .A1(N644), .A2(N2619) );
  AND2_X1 AND2_692( .ZN(N3155), .A1(N2533), .A2(N2269) );
  OR2_X1 OR2_693( .ZN(N3159), .A1(N1174), .A2(N2878) );
  INV_X2 NOT1_694( .ZN(N3167), .A(N2778) );
  AND2_X1 AND2_695( .ZN(N3168), .A1(N609), .A2(N2508) );
  AND2_X1 AND2_696( .ZN(N3169), .A1(N604), .A2(N2502) );
  AND2_X1 AND2_697( .ZN(N3173), .A1(N742), .A2(N2496) );
  AND2_X1 AND2_698( .ZN(N3178), .A1(N734), .A2(N2488) );
  AND2_X1 AND2_699( .ZN(N3184), .A1(N599), .A2(N2482) );
  AND2_X1 AND2_700( .ZN(N3185), .A1(N727), .A2(N2573) );
  AND2_X1 AND2_701( .ZN(N3189), .A1(N721), .A2(N2567) );
  AND2_X1 AND2_702( .ZN(N3195), .A1(N715), .A2(N2561) );
  AND2_X1 AND2_703( .ZN(N3202), .A1(N708), .A2(N2554) );
  AND2_X1 AND2_704( .ZN(N3210), .A1(N609), .A2(N2508) );
  AND2_X1 AND2_705( .ZN(N3211), .A1(N604), .A2(N2502) );
  AND2_X1 AND2_706( .ZN(N3215), .A1(N742), .A2(N2496) );
  AND2_X1 AND2_707( .ZN(N3221), .A1(N2488), .A2(N734) );
  AND2_X1 AND2_708( .ZN(N3228), .A1(N599), .A2(N2482) );
  AND2_X1 AND2_709( .ZN(N3229), .A1(N727), .A2(N2573) );
  AND2_X1 AND2_710( .ZN(N3232), .A1(N721), .A2(N2567) );
  AND2_X1 AND2_711( .ZN(N3236), .A1(N715), .A2(N2561) );
  AND2_X1 AND2_712( .ZN(N3241), .A1(N708), .A2(N2554) );
  OR2_X1 OR2_713( .ZN(N3247), .A1(N2913), .A2(N2299) );
  OR2_X1 OR2_714( .ZN(N3251), .A1(N2914), .A2(N2300) );
  OR2_X1 OR2_715( .ZN(N3255), .A1(N2915), .A2(N2301) );
  OR2_X1 OR2_716( .ZN(N3259), .A1(N2916), .A2(N2302) );
  OR2_X1 OR2_717( .ZN(N3263), .A1(N2917), .A2(N2303) );
  OR2_X1 OR2_718( .ZN(N3267), .A1(N2918), .A2(N2304) );
  OR2_X1 OR2_719( .ZN(N3273), .A1(N2919), .A2(N2305) );
  OR2_X1 OR2_720( .ZN(N3281), .A1(N2920), .A2(N2306) );
  OR2_X1 OR2_721( .ZN(N3287), .A1(N2921), .A2(N2307) );
  OR2_X1 OR2_722( .ZN(N3293), .A1(N2922), .A2(N2308) );
  OR2_X1 OR2_723( .ZN(N3299), .A1(N2924), .A2(N2322) );
  OR2_X1 OR2_724( .ZN(N3303), .A1(N2925), .A2(N2323) );
  OR2_X1 OR2_725( .ZN(N3307), .A1(N2926), .A2(N2324) );
  OR2_X1 OR2_726( .ZN(N3311), .A1(N2927), .A2(N2325) );
  OR2_X1 OR2_727( .ZN(N3315), .A1(N2929), .A2(N2327) );
  OR2_X1 OR2_728( .ZN(N3322), .A1(N2930), .A2(N2328) );
  OR2_X1 OR2_729( .ZN(N3328), .A1(N2931), .A2(N2329) );
  OR2_X1 OR2_730( .ZN(N3334), .A1(N2932), .A2(N2330) );
  OR2_X1 OR2_731( .ZN(N3340), .A1(N2934), .A2(N2343) );
  OR2_X1 OR2_732( .ZN(N3343), .A1(N2935), .A2(N2344) );
  OR2_X1 OR2_733( .ZN(N3349), .A1(N2936), .A2(N2345) );
  OR2_X1 OR2_734( .ZN(N3355), .A1(N2937), .A2(N2346) );
  AND2_X1 AND2_735( .ZN(N3361), .A1(N2761), .A2(N2478) );
  AND2_X1 AND2_736( .ZN(N3362), .A1(N2757), .A2(N2474) );
  AND2_X1 AND2_737( .ZN(N3363), .A1(N2753), .A2(N2470) );
  AND2_X1 AND2_738( .ZN(N3364), .A1(N2749), .A2(N2466) );
  AND2_X1 AND2_739( .ZN(N3365), .A1(N2745), .A2(N2462) );
  AND2_X1 AND2_740( .ZN(N3366), .A1(N2741), .A2(N2550) );
  AND2_X1 AND2_741( .ZN(N3367), .A1(N2737), .A2(N2546) );
  AND2_X1 AND2_742( .ZN(N3368), .A1(N2733), .A2(N2542) );
  AND2_X1 AND2_743( .ZN(N3369), .A1(N2729), .A2(N2538) );
  AND2_X1 AND2_744( .ZN(N3370), .A1(N2670), .A2(N2458) );
  AND2_X1 AND2_745( .ZN(N3371), .A1(N2666), .A2(N2454) );
  AND2_X1 AND2_746( .ZN(N3372), .A1(N2662), .A2(N2450) );
  AND2_X1 AND2_747( .ZN(N3373), .A1(N2658), .A2(N2446) );
  AND2_X1 AND2_748( .ZN(N3374), .A1(N2654), .A2(N2442) );
  AND2_X1 AND2_749( .ZN(N3375), .A1(N2988), .A2(N2650) );
  AND2_X1 AND2_750( .ZN(N3379), .A1(N2650), .A2(N1966) );
  INV_X1 NOT1_751( .ZN(N3380), .A(N2781) );
  AND2_X1 AND2_752( .ZN(N3381), .A1(N695), .A2(N2604) );
  OR2_X1 OR2_753( .ZN(N3384), .A1(N3005), .A2(N2379) );
  OR2_X1 OR2_754( .ZN(N3390), .A1(N3006), .A2(N2380) );
  OR2_X1 OR2_755( .ZN(N3398), .A1(N3007), .A2(N2381) );
  OR2_X1 OR2_756( .ZN(N3404), .A1(N3008), .A2(N2382) );
  OR2_X1 OR2_757( .ZN(N3410), .A1(N3009), .A2(N2383) );
  OR2_X1 OR2_758( .ZN(N3416), .A1(N3021), .A2(N2397) );
  OR2_X1 OR2_759( .ZN(N3420), .A1(N3022), .A2(N2398) );
  OR2_X1 OR2_760( .ZN(N3424), .A1(N3023), .A2(N2399) );
  OR2_X1 OR2_761( .ZN(N3428), .A1(N3024), .A2(N2400) );
  OR2_X1 OR2_762( .ZN(N3432), .A1(N3025), .A2(N2401) );
  OR2_X1 OR2_763( .ZN(N3436), .A1(N3026), .A2(N2402) );
  OR2_X1 OR2_764( .ZN(N3440), .A1(N3027), .A2(N2403) );
  OR2_X1 OR2_765( .ZN(N3444), .A1(N3028), .A2(N2404) );
  OR2_X1 OR2_766( .ZN(N3448), .A1(N3029), .A2(N2405) );
  INV_X1 NOT1_767( .ZN(N3452), .A(N2790) );
  INV_X1 NOT1_768( .ZN(N3453), .A(N2793) );
  OR2_X1 OR2_769( .ZN(N3454), .A1(N3034), .A2(N2420) );
  OR2_X1 OR2_770( .ZN(N3458), .A1(N3035), .A2(N2421) );
  OR2_X1 OR2_771( .ZN(N3462), .A1(N3036), .A2(N2422) );
  OR2_X1 OR2_772( .ZN(N3466), .A1(N3037), .A2(N2423) );
  OR2_X1 OR2_773( .ZN(N3470), .A1(N3038), .A2(N2424) );
  OR2_X1 OR2_774( .ZN(N3474), .A1(N3039), .A2(N2425) );
  OR2_X1 OR2_775( .ZN(N3478), .A1(N3040), .A2(N2426) );
  OR2_X1 OR2_776( .ZN(N3482), .A1(N3041), .A2(N2427) );
  INV_X1 NOT1_777( .ZN(N3486), .A(N2796) );
  BUF_X1 BUFF1_778( .Z(N3487), .A(N2644) );
  BUF_X1 BUFF1_779( .Z(N3490), .A(N2638) );
  BUF_X1 BUFF1_780( .Z(N3493), .A(N2632) );
  BUF_X1 BUFF1_781( .Z(N3496), .A(N2626) );
  BUF_X1 BUFF1_782( .Z(N3499), .A(N2619) );
  BUF_X1 BUFF1_783( .Z(N3502), .A(N2523) );
  NOR2_X2 NOR2_784( .ZN(N3507), .A1(N1167), .A2(N2868) );
  BUF_X1 BUFF1_785( .Z(N3510), .A(N2523) );
  NOR2_X1 NOR2_786( .ZN(N3515), .A1(N644), .A2(N2619) );
  BUF_X1 BUFF1_787( .Z(N3518), .A(N2644) );
  BUF_X1 BUFF1_788( .Z(N3521), .A(N2638) );
  BUF_X1 BUFF1_789( .Z(N3524), .A(N2632) );
  BUF_X1 BUFF1_790( .Z(N3527), .A(N2626) );
  BUF_X1 BUFF1_791( .Z(N3530), .A(N2619) );
  BUF_X1 BUFF1_792( .Z(N3535), .A(N2619) );
  BUF_X1 BUFF1_793( .Z(N3539), .A(N2632) );
  BUF_X1 BUFF1_794( .Z(N3542), .A(N2626) );
  BUF_X1 BUFF1_795( .Z(N3545), .A(N2644) );
  BUF_X1 BUFF1_796( .Z(N3548), .A(N2638) );
  INV_X2 NOT1_797( .ZN(N3551), .A(N2766) );
  INV_X1 NOT1_798( .ZN(N3552), .A(N2769) );
  BUF_X1 BUFF1_799( .Z(N3553), .A(N2442) );
  BUF_X1 BUFF1_800( .Z(N3557), .A(N2450) );
  BUF_X1 BUFF1_801( .Z(N3560), .A(N2446) );
  BUF_X1 BUFF1_802( .Z(N3563), .A(N2458) );
  BUF_X1 BUFF1_803( .Z(N3566), .A(N2454) );
  INV_X1 NOT1_804( .ZN(N3569), .A(N2772) );
  INV_X1 NOT1_805( .ZN(N3570), .A(N2775) );
  BUF_X1 BUFF1_806( .Z(N3571), .A(N2554) );
  BUF_X1 BUFF1_807( .Z(N3574), .A(N2567) );
  BUF_X1 BUFF1_808( .Z(N3577), .A(N2561) );
  BUF_X1 BUFF1_809( .Z(N3580), .A(N2482) );
  BUF_X4 BUFF1_810( .Z(N3583), .A(N2573) );
  BUF_X4 BUFF1_811( .Z(N3586), .A(N2496) );
  BUF_X1 BUFF1_812( .Z(N3589), .A(N2488) );
  BUF_X1 BUFF1_813( .Z(N3592), .A(N2508) );
  BUF_X1 BUFF1_814( .Z(N3595), .A(N2502) );
  BUF_X1 BUFF1_815( .Z(N3598), .A(N2508) );
  BUF_X1 BUFF1_816( .Z(N3601), .A(N2502) );
  BUF_X1 BUFF1_817( .Z(N3604), .A(N2496) );
  BUF_X1 BUFF1_818( .Z(N3607), .A(N2482) );
  BUF_X1 BUFF1_819( .Z(N3610), .A(N2573) );
  BUF_X1 BUFF1_820( .Z(N3613), .A(N2567) );
  BUF_X1 BUFF1_821( .Z(N3616), .A(N2561) );
  BUF_X1 BUFF1_822( .Z(N3619), .A(N2488) );
  BUF_X1 BUFF1_823( .Z(N3622), .A(N2554) );
  NOR2_X1 NOR2_824( .ZN(N3625), .A1(N734), .A2(N2488) );
  NOR2_X1 NOR2_825( .ZN(N3628), .A1(N708), .A2(N2554) );
  BUF_X1 BUFF1_826( .Z(N3631), .A(N2508) );
  BUF_X1 BUFF1_827( .Z(N3634), .A(N2502) );
  BUF_X1 BUFF1_828( .Z(N3637), .A(N2496) );
  BUF_X1 BUFF1_829( .Z(N3640), .A(N2488) );
  BUF_X1 BUFF1_830( .Z(N3643), .A(N2482) );
  BUF_X1 BUFF1_831( .Z(N3646), .A(N2573) );
  BUF_X1 BUFF1_832( .Z(N3649), .A(N2567) );
  BUF_X1 BUFF1_833( .Z(N3652), .A(N2561) );
  BUF_X1 BUFF1_834( .Z(N3655), .A(N2554) );
  NOR2_X1 NOR2_835( .ZN(N3658), .A1(N2488), .A2(N734) );
  BUF_X1 BUFF1_836( .Z(N3661), .A(N2674) );
  BUF_X1 BUFF1_837( .Z(N3664), .A(N2674) );
  BUF_X1 BUFF1_838( .Z(N3667), .A(N2761) );
  BUF_X1 BUFF1_839( .Z(N3670), .A(N2478) );
  BUF_X1 BUFF1_840( .Z(N3673), .A(N2757) );
  BUF_X1 BUFF1_841( .Z(N3676), .A(N2474) );
  BUF_X1 BUFF1_842( .Z(N3679), .A(N2753) );
  BUF_X1 BUFF1_843( .Z(N3682), .A(N2470) );
  BUF_X1 BUFF1_844( .Z(N3685), .A(N2745) );
  BUF_X1 BUFF1_845( .Z(N3688), .A(N2462) );
  BUF_X1 BUFF1_846( .Z(N3691), .A(N2741) );
  BUF_X1 BUFF1_847( .Z(N3694), .A(N2550) );
  BUF_X1 BUFF1_848( .Z(N3697), .A(N2737) );
  BUF_X1 BUFF1_849( .Z(N3700), .A(N2546) );
  BUF_X1 BUFF1_850( .Z(N3703), .A(N2733) );
  BUF_X1 BUFF1_851( .Z(N3706), .A(N2542) );
  BUF_X1 BUFF1_852( .Z(N3709), .A(N2749) );
  BUF_X1 BUFF1_853( .Z(N3712), .A(N2466) );
  BUF_X1 BUFF1_854( .Z(N3715), .A(N2729) );
  BUF_X1 BUFF1_855( .Z(N3718), .A(N2538) );
  BUF_X1 BUFF1_856( .Z(N3721), .A(N2704) );
  BUF_X1 BUFF1_857( .Z(N3724), .A(N2700) );
  BUF_X1 BUFF1_858( .Z(N3727), .A(N2696) );
  BUF_X1 BUFF1_859( .Z(N3730), .A(N2688) );
  BUF_X1 BUFF1_860( .Z(N3733), .A(N2692) );
  BUF_X1 BUFF1_861( .Z(N3736), .A(N2670) );
  BUF_X1 BUFF1_862( .Z(N3739), .A(N2458) );
  BUF_X1 BUFF1_863( .Z(N3742), .A(N2666) );
  BUF_X1 BUFF1_864( .Z(N3745), .A(N2454) );
  BUF_X1 BUFF1_865( .Z(N3748), .A(N2662) );
  BUF_X1 BUFF1_866( .Z(N3751), .A(N2450) );
  BUF_X1 BUFF1_867( .Z(N3754), .A(N2658) );
  BUF_X1 BUFF1_868( .Z(N3757), .A(N2446) );
  BUF_X1 BUFF1_869( .Z(N3760), .A(N2654) );
  BUF_X1 BUFF1_870( .Z(N3763), .A(N2442) );
  BUF_X1 BUFF1_871( .Z(N3766), .A(N2654) );
  BUF_X1 BUFF1_872( .Z(N3769), .A(N2662) );
  BUF_X1 BUFF1_873( .Z(N3772), .A(N2658) );
  BUF_X1 BUFF1_874( .Z(N3775), .A(N2670) );
  BUF_X1 BUFF1_875( .Z(N3778), .A(N2666) );
  INV_X1 NOT1_876( .ZN(N3781), .A(N2784) );
  INV_X1 NOT1_877( .ZN(N3782), .A(N2787) );
  OR2_X1 OR2_878( .ZN(N3783), .A1(N2928), .A2(N2326) );
  OR2_X1 OR2_879( .ZN(N3786), .A1(N2933), .A2(N2342) );
  OR2_X1 OR2_880( .ZN(N3789), .A1(N2923), .A2(N2321) );
  BUF_X1 BUFF1_881( .Z(N3792), .A(N2688) );
  BUF_X1 BUFF1_882( .Z(N3795), .A(N2696) );
  BUF_X1 BUFF1_883( .Z(N3798), .A(N2692) );
  BUF_X1 BUFF1_884( .Z(N3801), .A(N2704) );
  BUF_X1 BUFF1_885( .Z(N3804), .A(N2700) );
  BUF_X1 BUFF1_886( .Z(N3807), .A(N2604) );
  BUF_X1 BUFF1_887( .Z(N3810), .A(N2611) );
  BUF_X1 BUFF1_888( .Z(N3813), .A(N2607) );
  BUF_X1 BUFF1_889( .Z(N3816), .A(N2615) );
  BUF_X1 BUFF1_890( .Z(N3819), .A(N2538) );
  BUF_X1 BUFF1_891( .Z(N3822), .A(N2546) );
  BUF_X1 BUFF1_892( .Z(N3825), .A(N2542) );
  BUF_X1 BUFF1_893( .Z(N3828), .A(N2462) );
  BUF_X1 BUFF1_894( .Z(N3831), .A(N2550) );
  BUF_X1 BUFF1_895( .Z(N3834), .A(N2470) );
  BUF_X1 BUFF1_896( .Z(N3837), .A(N2466) );
  BUF_X1 BUFF1_897( .Z(N3840), .A(N2478) );
  BUF_X1 BUFF1_898( .Z(N3843), .A(N2474) );
  BUF_X1 BUFF1_899( .Z(N3846), .A(N2615) );
  BUF_X1 BUFF1_900( .Z(N3849), .A(N2611) );
  BUF_X1 BUFF1_901( .Z(N3852), .A(N2607) );
  BUF_X1 BUFF1_902( .Z(N3855), .A(N2680) );
  BUF_X1 BUFF1_903( .Z(N3858), .A(N2729) );
  BUF_X1 BUFF1_904( .Z(N3861), .A(N2737) );
  BUF_X1 BUFF1_905( .Z(N3864), .A(N2733) );
  BUF_X1 BUFF1_906( .Z(N3867), .A(N2745) );
  BUF_X1 BUFF1_907( .Z(N3870), .A(N2741) );
  BUF_X1 BUFF1_908( .Z(N3873), .A(N2753) );
  BUF_X1 BUFF1_909( .Z(N3876), .A(N2749) );
  BUF_X1 BUFF1_910( .Z(N3879), .A(N2761) );
  BUF_X1 BUFF1_911( .Z(N3882), .A(N2757) );
  OR2_X1 OR2_912( .ZN(N3885), .A1(N3033), .A2(N2419) );
  OR2_X1 OR2_913( .ZN(N3888), .A1(N3032), .A2(N2418) );
  OR2_X1 OR2_914( .ZN(N3891), .A1(N3020), .A2(N2396) );
  NAND2_X2 NAND2_915( .ZN(N3953), .A1(N3067), .A2(N2117) );
  INV_X2 NOT1_916( .ZN(N3954), .A(N3067) );
  NAND2_X1 NAND2_917( .ZN(N3955), .A1(N3070), .A2(N2537) );
  INV_X1 NOT1_918( .ZN(N3956), .A(N3070) );
  INV_X1 NOT1_919( .ZN(N3958), .A(N3073) );
  INV_X1 NOT1_920( .ZN(N3964), .A(N3080) );
  OR2_X1 OR2_921( .ZN(N4193), .A1(N1649), .A2(N3379) );
  OR3_X1 OR3_922( .ZN(N4303), .A1(N1167), .A2(N2867), .A3(N3130) );
  INV_X1 NOT1_923( .ZN(N4308), .A(N3061) );
  INV_X1 NOT1_924( .ZN(N4313), .A(N3064) );
  NAND2_X1 NAND2_925( .ZN(N4326), .A1(N2769), .A2(N3551) );
  NAND2_X1 NAND2_926( .ZN(N4327), .A1(N2766), .A2(N3552) );
  NAND2_X1 NAND2_927( .ZN(N4333), .A1(N2775), .A2(N3569) );
  NAND2_X1 NAND2_928( .ZN(N4334), .A1(N2772), .A2(N3570) );
  NAND2_X1 NAND2_929( .ZN(N4411), .A1(N2787), .A2(N3781) );
  NAND2_X1 NAND2_930( .ZN(N4412), .A1(N2784), .A2(N3782) );
  NAND2_X1 NAND2_931( .ZN(N4463), .A1(N3487), .A2(N1828) );
  INV_X1 NOT1_932( .ZN(N4464), .A(N3487) );
  NAND2_X1 NAND2_933( .ZN(N4465), .A1(N3490), .A2(N1829) );
  INV_X1 NOT1_934( .ZN(N4466), .A(N3490) );
  NAND2_X1 NAND2_935( .ZN(N4467), .A1(N3493), .A2(N2267) );
  INV_X1 NOT1_936( .ZN(N4468), .A(N3493) );
  NAND2_X1 NAND2_937( .ZN(N4469), .A1(N3496), .A2(N1830) );
  INV_X1 NOT1_938( .ZN(N4470), .A(N3496) );
  NAND2_X1 NAND2_939( .ZN(N4471), .A1(N3499), .A2(N1833) );
  INV_X1 NOT1_940( .ZN(N4472), .A(N3499) );
  INV_X1 NOT1_941( .ZN(N4473), .A(N3122) );
  INV_X1 NOT1_942( .ZN(N4474), .A(N3126) );
  NAND2_X1 NAND2_943( .ZN(N4475), .A1(N3518), .A2(N1840) );
  INV_X1 NOT1_944( .ZN(N4476), .A(N3518) );
  NAND2_X1 NAND2_945( .ZN(N4477), .A1(N3521), .A2(N1841) );
  INV_X1 NOT1_946( .ZN(N4478), .A(N3521) );
  NAND2_X1 NAND2_947( .ZN(N4479), .A1(N3524), .A2(N2275) );
  INV_X1 NOT1_948( .ZN(N4480), .A(N3524) );
  NAND2_X1 NAND2_949( .ZN(N4481), .A1(N3527), .A2(N1842) );
  INV_X1 NOT1_950( .ZN(N4482), .A(N3527) );
  NAND2_X1 NAND2_951( .ZN(N4483), .A1(N3530), .A2(N1843) );
  INV_X1 NOT1_952( .ZN(N4484), .A(N3530) );
  INV_X1 NOT1_953( .ZN(N4485), .A(N3155) );
  INV_X1 NOT1_954( .ZN(N4486), .A(N3159) );
  NAND2_X1 NAND2_955( .ZN(N4487), .A1(N1721), .A2(N3954) );
  NAND2_X1 NAND2_956( .ZN(N4488), .A1(N2235), .A2(N3956) );
  INV_X1 NOT1_957( .ZN(N4489), .A(N3535) );
  NAND2_X1 NAND2_958( .ZN(N4490), .A1(N3535), .A2(N3958) );
  INV_X1 NOT1_959( .ZN(N4491), .A(N3539) );
  INV_X1 NOT1_960( .ZN(N4492), .A(N3542) );
  INV_X1 NOT1_961( .ZN(N4493), .A(N3545) );
  INV_X1 NOT1_962( .ZN(N4494), .A(N3548) );
  INV_X1 NOT1_963( .ZN(N4495), .A(N3553) );
  NAND2_X1 NAND2_964( .ZN(N4496), .A1(N3553), .A2(N3964) );
  INV_X1 NOT1_965( .ZN(N4497), .A(N3557) );
  INV_X1 NOT1_966( .ZN(N4498), .A(N3560) );
  INV_X1 NOT1_967( .ZN(N4499), .A(N3563) );
  INV_X1 NOT1_968( .ZN(N4500), .A(N3566) );
  INV_X1 NOT1_969( .ZN(N4501), .A(N3571) );
  NAND2_X1 NAND2_970( .ZN(N4502), .A1(N3571), .A2(N3167) );
  INV_X1 NOT1_971( .ZN(N4503), .A(N3574) );
  INV_X1 NOT1_972( .ZN(N4504), .A(N3577) );
  INV_X1 NOT1_973( .ZN(N4505), .A(N3580) );
  INV_X1 NOT1_974( .ZN(N4506), .A(N3583) );
  NAND2_X1 NAND2_975( .ZN(N4507), .A1(N3598), .A2(N1867) );
  INV_X1 NOT1_976( .ZN(N4508), .A(N3598) );
  NAND2_X1 NAND2_977( .ZN(N4509), .A1(N3601), .A2(N1868) );
  INV_X1 NOT1_978( .ZN(N4510), .A(N3601) );
  NAND2_X1 NAND2_979( .ZN(N4511), .A1(N3604), .A2(N1869) );
  INV_X1 NOT1_980( .ZN(N4512), .A(N3604) );
  NAND2_X1 NAND2_981( .ZN(N4513), .A1(N3607), .A2(N1870) );
  INV_X1 NOT1_982( .ZN(N4514), .A(N3607) );
  NAND2_X1 NAND2_983( .ZN(N4515), .A1(N3610), .A2(N1871) );
  INV_X1 NOT1_984( .ZN(N4516), .A(N3610) );
  NAND2_X1 NAND2_985( .ZN(N4517), .A1(N3613), .A2(N1872) );
  INV_X1 NOT1_986( .ZN(N4518), .A(N3613) );
  NAND2_X1 NAND2_987( .ZN(N4519), .A1(N3616), .A2(N1873) );
  INV_X1 NOT1_988( .ZN(N4520), .A(N3616) );
  NAND2_X1 NAND2_989( .ZN(N4521), .A1(N3619), .A2(N1874) );
  INV_X1 NOT1_990( .ZN(N4522), .A(N3619) );
  NAND2_X1 NAND2_991( .ZN(N4523), .A1(N3622), .A2(N1875) );
  INV_X1 NOT1_992( .ZN(N4524), .A(N3622) );
  NAND2_X1 NAND2_993( .ZN(N4525), .A1(N3631), .A2(N1876) );
  INV_X1 NOT1_994( .ZN(N4526), .A(N3631) );
  NAND2_X1 NAND2_995( .ZN(N4527), .A1(N3634), .A2(N1877) );
  INV_X1 NOT1_996( .ZN(N4528), .A(N3634) );
  NAND2_X1 NAND2_997( .ZN(N4529), .A1(N3637), .A2(N1878) );
  INV_X1 NOT1_998( .ZN(N4530), .A(N3637) );
  NAND2_X1 NAND2_999( .ZN(N4531), .A1(N3640), .A2(N1879) );
  INV_X1 NOT1_1000( .ZN(N4532), .A(N3640) );
  NAND2_X1 NAND2_1001( .ZN(N4533), .A1(N3643), .A2(N1880) );
  INV_X1 NOT1_1002( .ZN(N4534), .A(N3643) );
  NAND2_X1 NAND2_1003( .ZN(N4535), .A1(N3646), .A2(N1881) );
  INV_X2 NOT1_1004( .ZN(N4536), .A(N3646) );
  NAND2_X1 NAND2_1005( .ZN(N4537), .A1(N3649), .A2(N1882) );
  INV_X1 NOT1_1006( .ZN(N4538), .A(N3649) );
  NAND2_X1 NAND2_1007( .ZN(N4539), .A1(N3652), .A2(N1883) );
  INV_X1 NOT1_1008( .ZN(N4540), .A(N3652) );
  NAND2_X1 NAND2_1009( .ZN(N4541), .A1(N3655), .A2(N1884) );
  INV_X1 NOT1_1010( .ZN(N4542), .A(N3655) );
  INV_X1 NOT1_1011( .ZN(N4543), .A(N3658) );
  AND2_X1 AND2_1012( .ZN(N4544), .A1(N806), .A2(N3293) );
  AND2_X1 AND2_1013( .ZN(N4545), .A1(N800), .A2(N3287) );
  AND2_X1 AND2_1014( .ZN(N4549), .A1(N794), .A2(N3281) );
  AND2_X1 AND2_1015( .ZN(N4555), .A1(N3273), .A2(N786) );
  AND2_X1 AND2_1016( .ZN(N4562), .A1(N780), .A2(N3267) );
  AND2_X1 AND2_1017( .ZN(N4563), .A1(N774), .A2(N3355) );
  AND2_X1 AND2_1018( .ZN(N4566), .A1(N768), .A2(N3349) );
  AND2_X1 AND2_1019( .ZN(N4570), .A1(N762), .A2(N3343) );
  INV_X1 NOT1_1020( .ZN(N4575), .A(N3661) );
  AND2_X1 AND2_1021( .ZN(N4576), .A1(N806), .A2(N3293) );
  AND2_X1 AND2_1022( .ZN(N4577), .A1(N800), .A2(N3287) );
  AND2_X1 AND2_1023( .ZN(N4581), .A1(N794), .A2(N3281) );
  AND2_X1 AND2_1024( .ZN(N4586), .A1(N786), .A2(N3273) );
  AND2_X1 AND2_1025( .ZN(N4592), .A1(N780), .A2(N3267) );
  AND2_X1 AND2_1026( .ZN(N4593), .A1(N774), .A2(N3355) );
  AND2_X1 AND2_1027( .ZN(N4597), .A1(N768), .A2(N3349) );
  AND2_X1 AND2_1028( .ZN(N4603), .A1(N762), .A2(N3343) );
  INV_X1 NOT1_1029( .ZN(N4610), .A(N3664) );
  INV_X1 NOT1_1030( .ZN(N4611), .A(N3667) );
  INV_X1 NOT1_1031( .ZN(N4612), .A(N3670) );
  INV_X1 NOT1_1032( .ZN(N4613), .A(N3673) );
  INV_X1 NOT1_1033( .ZN(N4614), .A(N3676) );
  INV_X1 NOT1_1034( .ZN(N4615), .A(N3679) );
  INV_X1 NOT1_1035( .ZN(N4616), .A(N3682) );
  INV_X1 NOT1_1036( .ZN(N4617), .A(N3685) );
  INV_X1 NOT1_1037( .ZN(N4618), .A(N3688) );
  INV_X1 NOT1_1038( .ZN(N4619), .A(N3691) );
  INV_X1 NOT1_1039( .ZN(N4620), .A(N3694) );
  INV_X1 NOT1_1040( .ZN(N4621), .A(N3697) );
  INV_X1 NOT1_1041( .ZN(N4622), .A(N3700) );
  INV_X1 NOT1_1042( .ZN(N4623), .A(N3703) );
  INV_X1 NOT1_1043( .ZN(N4624), .A(N3706) );
  INV_X1 NOT1_1044( .ZN(N4625), .A(N3709) );
  INV_X1 NOT1_1045( .ZN(N4626), .A(N3712) );
  INV_X1 NOT1_1046( .ZN(N4627), .A(N3715) );
  INV_X1 NOT1_1047( .ZN(N4628), .A(N3718) );
  INV_X1 NOT1_1048( .ZN(N4629), .A(N3721) );
  AND2_X1 AND2_1049( .ZN(N4630), .A1(N3448), .A2(N2704) );
  INV_X1 NOT1_1050( .ZN(N4631), .A(N3724) );
  AND2_X1 AND2_1051( .ZN(N4632), .A1(N3444), .A2(N2700) );
  INV_X1 NOT1_1052( .ZN(N4633), .A(N3727) );
  AND2_X1 AND2_1053( .ZN(N4634), .A1(N3440), .A2(N2696) );
  AND2_X1 AND2_1054( .ZN(N4635), .A1(N3436), .A2(N2692) );
  INV_X1 NOT1_1055( .ZN(N4636), .A(N3730) );
  AND2_X1 AND2_1056( .ZN(N4637), .A1(N3432), .A2(N2688) );
  AND2_X1 AND2_1057( .ZN(N4638), .A1(N3428), .A2(N3311) );
  AND2_X1 AND2_1058( .ZN(N4639), .A1(N3424), .A2(N3307) );
  AND2_X1 AND2_1059( .ZN(N4640), .A1(N3420), .A2(N3303) );
  AND2_X1 AND2_1060( .ZN(N4641), .A1(N3416), .A2(N3299) );
  INV_X1 NOT1_1061( .ZN(N4642), .A(N3733) );
  INV_X1 NOT1_1062( .ZN(N4643), .A(N3736) );
  INV_X1 NOT1_1063( .ZN(N4644), .A(N3739) );
  INV_X1 NOT1_1064( .ZN(N4645), .A(N3742) );
  INV_X1 NOT1_1065( .ZN(N4646), .A(N3745) );
  INV_X1 NOT1_1066( .ZN(N4647), .A(N3748) );
  INV_X1 NOT1_1067( .ZN(N4648), .A(N3751) );
  INV_X1 NOT1_1068( .ZN(N4649), .A(N3754) );
  INV_X1 NOT1_1069( .ZN(N4650), .A(N3757) );
  INV_X1 NOT1_1070( .ZN(N4651), .A(N3760) );
  INV_X1 NOT1_1071( .ZN(N4652), .A(N3763) );
  INV_X1 NOT1_1072( .ZN(N4653), .A(N3375) );
  AND2_X1 AND2_1073( .ZN(N4656), .A1(N865), .A2(N3410) );
  AND2_X1 AND2_1074( .ZN(N4657), .A1(N859), .A2(N3404) );
  AND2_X1 AND2_1075( .ZN(N4661), .A1(N853), .A2(N3398) );
  AND2_X1 AND2_1076( .ZN(N4667), .A1(N3390), .A2(N845) );
  AND2_X1 AND2_1077( .ZN(N4674), .A1(N839), .A2(N3384) );
  AND2_X1 AND2_1078( .ZN(N4675), .A1(N833), .A2(N3334) );
  AND2_X1 AND2_1079( .ZN(N4678), .A1(N827), .A2(N3328) );
  AND2_X1 AND2_1080( .ZN(N4682), .A1(N821), .A2(N3322) );
  AND2_X1 AND2_1081( .ZN(N4687), .A1(N814), .A2(N3315) );
  INV_X1 NOT1_1082( .ZN(N4693), .A(N3766) );
  NAND2_X2 NAND2_1083( .ZN(N4694), .A1(N3766), .A2(N3380) );
  INV_X1 NOT1_1084( .ZN(N4695), .A(N3769) );
  INV_X1 NOT1_1085( .ZN(N4696), .A(N3772) );
  INV_X1 NOT1_1086( .ZN(N4697), .A(N3775) );
  INV_X1 NOT1_1087( .ZN(N4698), .A(N3778) );
  INV_X1 NOT1_1088( .ZN(N4699), .A(N3783) );
  INV_X1 NOT1_1089( .ZN(N4700), .A(N3786) );
  AND2_X1 AND2_1090( .ZN(N4701), .A1(N865), .A2(N3410) );
  AND2_X1 AND2_1091( .ZN(N4702), .A1(N859), .A2(N3404) );
  AND2_X1 AND2_1092( .ZN(N4706), .A1(N853), .A2(N3398) );
  AND2_X1 AND2_1093( .ZN(N4711), .A1(N845), .A2(N3390) );
  AND2_X1 AND2_1094( .ZN(N4717), .A1(N839), .A2(N3384) );
  AND2_X1 AND2_1095( .ZN(N4718), .A1(N833), .A2(N3334) );
  AND2_X1 AND2_1096( .ZN(N4722), .A1(N827), .A2(N3328) );
  AND2_X1 AND2_1097( .ZN(N4728), .A1(N821), .A2(N3322) );
  AND2_X1 AND2_1098( .ZN(N4735), .A1(N814), .A2(N3315) );
  INV_X1 NOT1_1099( .ZN(N4743), .A(N3789) );
  INV_X1 NOT1_1100( .ZN(N4744), .A(N3792) );
  INV_X1 NOT1_1101( .ZN(N4745), .A(N3807) );
  NAND2_X1 NAND2_1102( .ZN(N4746), .A1(N3807), .A2(N3452) );
  INV_X1 NOT1_1103( .ZN(N4747), .A(N3810) );
  INV_X1 NOT1_1104( .ZN(N4748), .A(N3813) );
  INV_X1 NOT1_1105( .ZN(N4749), .A(N3816) );
  INV_X1 NOT1_1106( .ZN(N4750), .A(N3819) );
  NAND2_X1 NAND2_1107( .ZN(N4751), .A1(N3819), .A2(N3453) );
  INV_X1 NOT1_1108( .ZN(N4752), .A(N3822) );
  INV_X1 NOT1_1109( .ZN(N4753), .A(N3825) );
  INV_X1 NOT1_1110( .ZN(N4754), .A(N3828) );
  INV_X1 NOT1_1111( .ZN(N4755), .A(N3831) );
  AND2_X1 AND2_1112( .ZN(N4756), .A1(N3482), .A2(N3263) );
  AND2_X1 AND2_1113( .ZN(N4757), .A1(N3478), .A2(N3259) );
  AND2_X1 AND2_1114( .ZN(N4758), .A1(N3474), .A2(N3255) );
  AND2_X1 AND2_1115( .ZN(N4759), .A1(N3470), .A2(N3251) );
  AND2_X1 AND2_1116( .ZN(N4760), .A1(N3466), .A2(N3247) );
  INV_X1 NOT1_1117( .ZN(N4761), .A(N3846) );
  AND2_X1 AND2_1118( .ZN(N4762), .A1(N3462), .A2(N2615) );
  INV_X1 NOT1_1119( .ZN(N4763), .A(N3849) );
  AND2_X1 AND2_1120( .ZN(N4764), .A1(N3458), .A2(N2611) );
  INV_X1 NOT1_1121( .ZN(N4765), .A(N3852) );
  AND2_X1 AND2_1122( .ZN(N4766), .A1(N3454), .A2(N2607) );
  AND2_X1 AND2_1123( .ZN(N4767), .A1(N2680), .A2(N3381) );
  INV_X1 NOT1_1124( .ZN(N4768), .A(N3855) );
  AND2_X1 AND2_1125( .ZN(N4769), .A1(N3340), .A2(N695) );
  INV_X1 NOT1_1126( .ZN(N4775), .A(N3858) );
  NAND2_X1 NAND2_1127( .ZN(N4776), .A1(N3858), .A2(N3486) );
  INV_X1 NOT1_1128( .ZN(N4777), .A(N3861) );
  INV_X1 NOT1_1129( .ZN(N4778), .A(N3864) );
  INV_X1 NOT1_1130( .ZN(N4779), .A(N3867) );
  INV_X1 NOT1_1131( .ZN(N4780), .A(N3870) );
  INV_X1 NOT1_1132( .ZN(N4781), .A(N3885) );
  INV_X1 NOT1_1133( .ZN(N4782), .A(N3888) );
  INV_X1 NOT1_1134( .ZN(N4783), .A(N3891) );
  OR2_X1 OR2_1135( .ZN(N4784), .A1(N3131), .A2(N3134) );
  INV_X1 NOT1_1136( .ZN(N4789), .A(N3502) );
  INV_X1 NOT1_1137( .ZN(N4790), .A(N3131) );
  INV_X1 NOT1_1138( .ZN(N4793), .A(N3507) );
  INV_X1 NOT1_1139( .ZN(N4794), .A(N3510) );
  INV_X1 NOT1_1140( .ZN(N4795), .A(N3515) );
  BUF_X4 BUFF1_1141( .Z(N4796), .A(N3114) );
  INV_X1 NOT1_1142( .ZN(N4799), .A(N3586) );
  INV_X1 NOT1_1143( .ZN(N4800), .A(N3589) );
  INV_X1 NOT1_1144( .ZN(N4801), .A(N3592) );
  INV_X1 NOT1_1145( .ZN(N4802), .A(N3595) );
  NAND2_X1 NAND2_1146( .ZN(N4803), .A1(N4326), .A2(N4327) );
  NAND2_X1 NAND2_1147( .ZN(N4806), .A1(N4333), .A2(N4334) );
  INV_X1 NOT1_1148( .ZN(N4809), .A(N3625) );
  BUF_X1 BUFF1_1149( .Z(N4810), .A(N3178) );
  INV_X2 NOT1_1150( .ZN(N4813), .A(N3628) );
  BUF_X1 BUFF1_1151( .Z(N4814), .A(N3202) );
  BUF_X1 BUFF1_1152( .Z(N4817), .A(N3221) );
  BUF_X1 BUFF1_1153( .Z(N4820), .A(N3293) );
  BUF_X1 BUFF1_1154( .Z(N4823), .A(N3287) );
  BUF_X1 BUFF1_1155( .Z(N4826), .A(N3281) );
  BUF_X1 BUFF1_1156( .Z(N4829), .A(N3273) );
  BUF_X1 BUFF1_1157( .Z(N4832), .A(N3267) );
  BUF_X1 BUFF1_1158( .Z(N4835), .A(N3355) );
  BUF_X1 BUFF1_1159( .Z(N4838), .A(N3349) );
  BUF_X1 BUFF1_1160( .Z(N4841), .A(N3343) );
  NOR2_X2 NOR2_1161( .ZN(N4844), .A1(N3273), .A2(N786) );
  BUF_X1 BUFF1_1162( .Z(N4847), .A(N3293) );
  BUF_X1 BUFF1_1163( .Z(N4850), .A(N3287) );
  BUF_X1 BUFF1_1164( .Z(N4853), .A(N3281) );
  BUF_X1 BUFF1_1165( .Z(N4856), .A(N3267) );
  BUF_X1 BUFF1_1166( .Z(N4859), .A(N3355) );
  BUF_X1 BUFF1_1167( .Z(N4862), .A(N3349) );
  BUF_X1 BUFF1_1168( .Z(N4865), .A(N3343) );
  BUF_X1 BUFF1_1169( .Z(N4868), .A(N3273) );
  NOR2_X1 NOR2_1170( .ZN(N4871), .A1(N786), .A2(N3273) );
  BUF_X1 BUFF1_1171( .Z(N4874), .A(N3448) );
  BUF_X1 BUFF1_1172( .Z(N4877), .A(N3444) );
  BUF_X1 BUFF1_1173( .Z(N4880), .A(N3440) );
  BUF_X1 BUFF1_1174( .Z(N4883), .A(N3432) );
  BUF_X1 BUFF1_1175( .Z(N4886), .A(N3428) );
  BUF_X1 BUFF1_1176( .Z(N4889), .A(N3311) );
  BUF_X1 BUFF1_1177( .Z(N4892), .A(N3424) );
  BUF_X1 BUFF1_1178( .Z(N4895), .A(N3307) );
  BUF_X1 BUFF1_1179( .Z(N4898), .A(N3420) );
  BUF_X1 BUFF1_1180( .Z(N4901), .A(N3303) );
  BUF_X1 BUFF1_1181( .Z(N4904), .A(N3436) );
  BUF_X1 BUFF1_1182( .Z(N4907), .A(N3416) );
  BUF_X1 BUFF1_1183( .Z(N4910), .A(N3299) );
  BUF_X1 BUFF1_1184( .Z(N4913), .A(N3410) );
  BUF_X1 BUFF1_1185( .Z(N4916), .A(N3404) );
  BUF_X1 BUFF1_1186( .Z(N4919), .A(N3398) );
  BUF_X1 BUFF1_1187( .Z(N4922), .A(N3390) );
  BUF_X1 BUFF1_1188( .Z(N4925), .A(N3384) );
  BUF_X1 BUFF1_1189( .Z(N4928), .A(N3334) );
  BUF_X1 BUFF1_1190( .Z(N4931), .A(N3328) );
  BUF_X1 BUFF1_1191( .Z(N4934), .A(N3322) );
  BUF_X1 BUFF1_1192( .Z(N4937), .A(N3315) );
  NOR2_X1 NOR2_1193( .ZN(N4940), .A1(N3390), .A2(N845) );
  BUF_X1 BUFF1_1194( .Z(N4943), .A(N3315) );
  BUF_X1 BUFF1_1195( .Z(N4946), .A(N3328) );
  BUF_X1 BUFF1_1196( .Z(N4949), .A(N3322) );
  BUF_X1 BUFF1_1197( .Z(N4952), .A(N3384) );
  BUF_X1 BUFF1_1198( .Z(N4955), .A(N3334) );
  BUF_X1 BUFF1_1199( .Z(N4958), .A(N3398) );
  BUF_X1 BUFF1_1200( .Z(N4961), .A(N3390) );
  BUF_X1 BUFF1_1201( .Z(N4964), .A(N3410) );
  BUF_X1 BUFF1_1202( .Z(N4967), .A(N3404) );
  BUF_X1 BUFF1_1203( .Z(N4970), .A(N3340) );
  BUF_X1 BUFF1_1204( .Z(N4973), .A(N3349) );
  BUF_X1 BUFF1_1205( .Z(N4976), .A(N3343) );
  BUF_X1 BUFF1_1206( .Z(N4979), .A(N3267) );
  BUF_X1 BUFF1_1207( .Z(N4982), .A(N3355) );
  BUF_X1 BUFF1_1208( .Z(N4985), .A(N3281) );
  BUF_X1 BUFF1_1209( .Z(N4988), .A(N3273) );
  BUF_X1 BUFF1_1210( .Z(N4991), .A(N3293) );
  BUF_X1 BUFF1_1211( .Z(N4994), .A(N3287) );
  NAND2_X1 NAND2_1212( .ZN(N4997), .A1(N4411), .A2(N4412) );
  BUF_X1 BUFF1_1213( .Z(N5000), .A(N3410) );
  BUF_X1 BUFF1_1214( .Z(N5003), .A(N3404) );
  BUF_X1 BUFF1_1215( .Z(N5006), .A(N3398) );
  BUF_X1 BUFF1_1216( .Z(N5009), .A(N3384) );
  BUF_X1 BUFF1_1217( .Z(N5012), .A(N3334) );
  BUF_X1 BUFF1_1218( .Z(N5015), .A(N3328) );
  BUF_X1 BUFF1_1219( .Z(N5018), .A(N3322) );
  BUF_X1 BUFF1_1220( .Z(N5021), .A(N3390) );
  BUF_X1 BUFF1_1221( .Z(N5024), .A(N3315) );
  NOR2_X1 NOR2_1222( .ZN(N5027), .A1(N845), .A2(N3390) );
  NOR2_X1 NOR2_1223( .ZN(N5030), .A1(N814), .A2(N3315) );
  BUF_X1 BUFF1_1224( .Z(N5033), .A(N3299) );
  BUF_X1 BUFF1_1225( .Z(N5036), .A(N3307) );
  BUF_X1 BUFF1_1226( .Z(N5039), .A(N3303) );
  BUF_X1 BUFF1_1227( .Z(N5042), .A(N3311) );
  INV_X2 NOT1_1228( .ZN(N5045), .A(N3795) );
  INV_X1 NOT1_1229( .ZN(N5046), .A(N3798) );
  INV_X1 NOT1_1230( .ZN(N5047), .A(N3801) );
  INV_X1 NOT1_1231( .ZN(N5048), .A(N3804) );
  BUF_X1 BUFF1_1232( .Z(N5049), .A(N3247) );
  BUF_X4 BUFF1_1233( .Z(N5052), .A(N3255) );
  BUF_X1 BUFF1_1234( .Z(N5055), .A(N3251) );
  BUF_X1 BUFF1_1235( .Z(N5058), .A(N3263) );
  BUF_X1 BUFF1_1236( .Z(N5061), .A(N3259) );
  INV_X1 NOT1_1237( .ZN(N5064), .A(N3834) );
  INV_X1 NOT1_1238( .ZN(N5065), .A(N3837) );
  INV_X1 NOT1_1239( .ZN(N5066), .A(N3840) );
  INV_X1 NOT1_1240( .ZN(N5067), .A(N3843) );
  BUF_X1 BUFF1_1241( .Z(N5068), .A(N3482) );
  BUF_X1 BUFF1_1242( .Z(N5071), .A(N3263) );
  BUF_X1 BUFF1_1243( .Z(N5074), .A(N3478) );
  BUF_X1 BUFF1_1244( .Z(N5077), .A(N3259) );
  BUF_X1 BUFF1_1245( .Z(N5080), .A(N3474) );
  BUF_X1 BUFF1_1246( .Z(N5083), .A(N3255) );
  BUF_X1 BUFF1_1247( .Z(N5086), .A(N3466) );
  BUF_X1 BUFF1_1248( .Z(N5089), .A(N3247) );
  BUF_X1 BUFF1_1249( .Z(N5092), .A(N3462) );
  BUF_X1 BUFF1_1250( .Z(N5095), .A(N3458) );
  BUF_X1 BUFF1_1251( .Z(N5098), .A(N3454) );
  BUF_X1 BUFF1_1252( .Z(N5101), .A(N3470) );
  BUF_X1 BUFF1_1253( .Z(N5104), .A(N3251) );
  BUF_X1 BUFF1_1254( .Z(N5107), .A(N3381) );
  INV_X1 NOT1_1255( .ZN(N5110), .A(N3873) );
  INV_X1 NOT1_1256( .ZN(N5111), .A(N3876) );
  INV_X1 NOT1_1257( .ZN(N5112), .A(N3879) );
  INV_X1 NOT1_1258( .ZN(N5113), .A(N3882) );
  BUF_X1 BUFF1_1259( .Z(N5114), .A(N3458) );
  BUF_X1 BUFF1_1260( .Z(N5117), .A(N3454) );
  BUF_X1 BUFF1_1261( .Z(N5120), .A(N3466) );
  BUF_X1 BUFF1_1262( .Z(N5123), .A(N3462) );
  BUF_X1 BUFF1_1263( .Z(N5126), .A(N3474) );
  BUF_X1 BUFF1_1264( .Z(N5129), .A(N3470) );
  BUF_X1 BUFF1_1265( .Z(N5132), .A(N3482) );
  BUF_X1 BUFF1_1266( .Z(N5135), .A(N3478) );
  BUF_X1 BUFF1_1267( .Z(N5138), .A(N3416) );
  BUF_X1 BUFF1_1268( .Z(N5141), .A(N3424) );
  BUF_X1 BUFF1_1269( .Z(N5144), .A(N3420) );
  BUF_X1 BUFF1_1270( .Z(N5147), .A(N3432) );
  BUF_X1 BUFF1_1271( .Z(N5150), .A(N3428) );
  BUF_X1 BUFF1_1272( .Z(N5153), .A(N3440) );
  BUF_X1 BUFF1_1273( .Z(N5156), .A(N3436) );
  BUF_X1 BUFF1_1274( .Z(N5159), .A(N3448) );
  BUF_X1 BUFF1_1275( .Z(N5162), .A(N3444) );
  NAND2_X2 NAND2_1276( .ZN(N5165), .A1(N4486), .A2(N4485) );
  NAND2_X2 NAND2_1277( .ZN(N5166), .A1(N4474), .A2(N4473) );
  NAND2_X2 NAND2_1278( .ZN(N5167), .A1(N1290), .A2(N4464) );
  NAND2_X2 NAND2_1279( .ZN(N5168), .A1(N1293), .A2(N4466) );
  NAND2_X2 NAND2_1280( .ZN(N5169), .A1(N2074), .A2(N4468) );
  NAND2_X2 NAND2_1281( .ZN(N5170), .A1(N1296), .A2(N4470) );
  NAND2_X2 NAND2_1282( .ZN(N5171), .A1(N1302), .A2(N4472) );
  NAND2_X1 NAND2_1283( .ZN(N5172), .A1(N1314), .A2(N4476) );
  NAND2_X1 NAND2_1284( .ZN(N5173), .A1(N1317), .A2(N4478) );
  NAND2_X1 NAND2_1285( .ZN(N5174), .A1(N2081), .A2(N4480) );
  NAND2_X1 NAND2_1286( .ZN(N5175), .A1(N1320), .A2(N4482) );
  NAND2_X1 NAND2_1287( .ZN(N5176), .A1(N1323), .A2(N4484) );
  NAND2_X1 NAND2_1288( .ZN(N5177), .A1(N3953), .A2(N4487) );
  NAND2_X1 NAND2_1289( .ZN(N5178), .A1(N3955), .A2(N4488) );
  NAND2_X1 NAND2_1290( .ZN(N5179), .A1(N3073), .A2(N4489) );
  NAND2_X1 NAND2_1291( .ZN(N5180), .A1(N3542), .A2(N4491) );
  NAND2_X1 NAND2_1292( .ZN(N5181), .A1(N3539), .A2(N4492) );
  NAND2_X1 NAND2_1293( .ZN(N5182), .A1(N3548), .A2(N4493) );
  NAND2_X1 NAND2_1294( .ZN(N5183), .A1(N3545), .A2(N4494) );
  NAND2_X1 NAND2_1295( .ZN(N5184), .A1(N3080), .A2(N4495) );
  NAND2_X1 NAND2_1296( .ZN(N5185), .A1(N3560), .A2(N4497) );
  NAND2_X1 NAND2_1297( .ZN(N5186), .A1(N3557), .A2(N4498) );
  NAND2_X1 NAND2_1298( .ZN(N5187), .A1(N3566), .A2(N4499) );
  NAND2_X1 NAND2_1299( .ZN(N5188), .A1(N3563), .A2(N4500) );
  NAND2_X1 NAND2_1300( .ZN(N5189), .A1(N2778), .A2(N4501) );
  NAND2_X1 NAND2_1301( .ZN(N5190), .A1(N3577), .A2(N4503) );
  NAND2_X1 NAND2_1302( .ZN(N5191), .A1(N3574), .A2(N4504) );
  NAND2_X1 NAND2_1303( .ZN(N5192), .A1(N3583), .A2(N4505) );
  NAND2_X1 NAND2_1304( .ZN(N5193), .A1(N3580), .A2(N4506) );
  NAND2_X1 NAND2_1305( .ZN(N5196), .A1(N1326), .A2(N4508) );
  NAND2_X1 NAND2_1306( .ZN(N5197), .A1(N1329), .A2(N4510) );
  NAND2_X1 NAND2_1307( .ZN(N5198), .A1(N1332), .A2(N4512) );
  NAND2_X1 NAND2_1308( .ZN(N5199), .A1(N1335), .A2(N4514) );
  NAND2_X1 NAND2_1309( .ZN(N5200), .A1(N1338), .A2(N4516) );
  NAND2_X1 NAND2_1310( .ZN(N5201), .A1(N1341), .A2(N4518) );
  NAND2_X1 NAND2_1311( .ZN(N5202), .A1(N1344), .A2(N4520) );
  NAND2_X1 NAND2_1312( .ZN(N5203), .A1(N1347), .A2(N4522) );
  NAND2_X1 NAND2_1313( .ZN(N5204), .A1(N1350), .A2(N4524) );
  NAND2_X1 NAND2_1314( .ZN(N5205), .A1(N1353), .A2(N4526) );
  NAND2_X1 NAND2_1315( .ZN(N5206), .A1(N1356), .A2(N4528) );
  NAND2_X1 NAND2_1316( .ZN(N5207), .A1(N1359), .A2(N4530) );
  NAND2_X1 NAND2_1317( .ZN(N5208), .A1(N1362), .A2(N4532) );
  NAND2_X1 NAND2_1318( .ZN(N5209), .A1(N1365), .A2(N4534) );
  NAND2_X1 NAND2_1319( .ZN(N5210), .A1(N1368), .A2(N4536) );
  NAND2_X1 NAND2_1320( .ZN(N5211), .A1(N1371), .A2(N4538) );
  NAND2_X1 NAND2_1321( .ZN(N5212), .A1(N1374), .A2(N4540) );
  NAND2_X1 NAND2_1322( .ZN(N5213), .A1(N1377), .A2(N4542) );
  NAND2_X1 NAND2_1323( .ZN(N5283), .A1(N3670), .A2(N4611) );
  NAND2_X1 NAND2_1324( .ZN(N5284), .A1(N3667), .A2(N4612) );
  NAND2_X1 NAND2_1325( .ZN(N5285), .A1(N3676), .A2(N4613) );
  NAND2_X1 NAND2_1326( .ZN(N5286), .A1(N3673), .A2(N4614) );
  NAND2_X1 NAND2_1327( .ZN(N5287), .A1(N3682), .A2(N4615) );
  NAND2_X1 NAND2_1328( .ZN(N5288), .A1(N3679), .A2(N4616) );
  NAND2_X1 NAND2_1329( .ZN(N5289), .A1(N3688), .A2(N4617) );
  NAND2_X1 NAND2_1330( .ZN(N5290), .A1(N3685), .A2(N4618) );
  NAND2_X1 NAND2_1331( .ZN(N5291), .A1(N3694), .A2(N4619) );
  NAND2_X1 NAND2_1332( .ZN(N5292), .A1(N3691), .A2(N4620) );
  NAND2_X1 NAND2_1333( .ZN(N5293), .A1(N3700), .A2(N4621) );
  NAND2_X1 NAND2_1334( .ZN(N5294), .A1(N3697), .A2(N4622) );
  NAND2_X1 NAND2_1335( .ZN(N5295), .A1(N3706), .A2(N4623) );
  NAND2_X1 NAND2_1336( .ZN(N5296), .A1(N3703), .A2(N4624) );
  NAND2_X1 NAND2_1337( .ZN(N5297), .A1(N3712), .A2(N4625) );
  NAND2_X1 NAND2_1338( .ZN(N5298), .A1(N3709), .A2(N4626) );
  NAND2_X1 NAND2_1339( .ZN(N5299), .A1(N3718), .A2(N4627) );
  NAND2_X1 NAND2_1340( .ZN(N5300), .A1(N3715), .A2(N4628) );
  NAND2_X1 NAND2_1341( .ZN(N5314), .A1(N3739), .A2(N4643) );
  NAND2_X1 NAND2_1342( .ZN(N5315), .A1(N3736), .A2(N4644) );
  NAND2_X1 NAND2_1343( .ZN(N5316), .A1(N3745), .A2(N4645) );
  NAND2_X1 NAND2_1344( .ZN(N5317), .A1(N3742), .A2(N4646) );
  NAND2_X1 NAND2_1345( .ZN(N5318), .A1(N3751), .A2(N4647) );
  NAND2_X1 NAND2_1346( .ZN(N5319), .A1(N3748), .A2(N4648) );
  NAND2_X1 NAND2_1347( .ZN(N5320), .A1(N3757), .A2(N4649) );
  NAND2_X1 NAND2_1348( .ZN(N5321), .A1(N3754), .A2(N4650) );
  NAND2_X1 NAND2_1349( .ZN(N5322), .A1(N3763), .A2(N4651) );
  NAND2_X1 NAND2_1350( .ZN(N5323), .A1(N3760), .A2(N4652) );
  INV_X1 NOT1_1351( .ZN(N5324), .A(N4193) );
  NAND2_X1 NAND2_1352( .ZN(N5363), .A1(N2781), .A2(N4693) );
  NAND2_X1 NAND2_1353( .ZN(N5364), .A1(N3772), .A2(N4695) );
  NAND2_X1 NAND2_1354( .ZN(N5365), .A1(N3769), .A2(N4696) );
  NAND2_X1 NAND2_1355( .ZN(N5366), .A1(N3778), .A2(N4697) );
  NAND2_X1 NAND2_1356( .ZN(N5367), .A1(N3775), .A2(N4698) );
  NAND2_X1 NAND2_1357( .ZN(N5425), .A1(N2790), .A2(N4745) );
  NAND2_X1 NAND2_1358( .ZN(N5426), .A1(N3813), .A2(N4747) );
  NAND2_X1 NAND2_1359( .ZN(N5427), .A1(N3810), .A2(N4748) );
  NAND2_X1 NAND2_1360( .ZN(N5429), .A1(N2793), .A2(N4750) );
  NAND2_X1 NAND2_1361( .ZN(N5430), .A1(N3825), .A2(N4752) );
  NAND2_X1 NAND2_1362( .ZN(N5431), .A1(N3822), .A2(N4753) );
  NAND2_X1 NAND2_1363( .ZN(N5432), .A1(N3831), .A2(N4754) );
  NAND2_X1 NAND2_1364( .ZN(N5433), .A1(N3828), .A2(N4755) );
  NAND2_X1 NAND2_1365( .ZN(N5451), .A1(N2796), .A2(N4775) );
  NAND2_X1 NAND2_1366( .ZN(N5452), .A1(N3864), .A2(N4777) );
  NAND2_X1 NAND2_1367( .ZN(N5453), .A1(N3861), .A2(N4778) );
  NAND2_X2 NAND2_1368( .ZN(N5454), .A1(N3870), .A2(N4779) );
  NAND2_X2 NAND2_1369( .ZN(N5455), .A1(N3867), .A2(N4780) );
  NAND2_X1 NAND2_1370( .ZN(N5456), .A1(N3888), .A2(N4781) );
  NAND2_X1 NAND2_1371( .ZN(N5457), .A1(N3885), .A2(N4782) );
  INV_X2 NOT1_1372( .ZN(N5469), .A(N4303) );
  NAND2_X1 NAND2_1373( .ZN(N5474), .A1(N3589), .A2(N4799) );
  NAND2_X1 NAND2_1374( .ZN(N5475), .A1(N3586), .A2(N4800) );
  NAND2_X1 NAND2_1375( .ZN(N5476), .A1(N3595), .A2(N4801) );
  NAND2_X1 NAND2_1376( .ZN(N5477), .A1(N3592), .A2(N4802) );
  NAND2_X1 NAND2_1377( .ZN(N5571), .A1(N3798), .A2(N5045) );
  NAND2_X1 NAND2_1378( .ZN(N5572), .A1(N3795), .A2(N5046) );
  NAND2_X1 NAND2_1379( .ZN(N5573), .A1(N3804), .A2(N5047) );
  NAND2_X1 NAND2_1380( .ZN(N5574), .A1(N3801), .A2(N5048) );
  NAND2_X1 NAND2_1381( .ZN(N5584), .A1(N3837), .A2(N5064) );
  NAND2_X1 NAND2_1382( .ZN(N5585), .A1(N3834), .A2(N5065) );
  NAND2_X1 NAND2_1383( .ZN(N5586), .A1(N3843), .A2(N5066) );
  NAND2_X1 NAND2_1384( .ZN(N5587), .A1(N3840), .A2(N5067) );
  NAND2_X1 NAND2_1385( .ZN(N5602), .A1(N3876), .A2(N5110) );
  NAND2_X1 NAND2_1386( .ZN(N5603), .A1(N3873), .A2(N5111) );
  NAND2_X1 NAND2_1387( .ZN(N5604), .A1(N3882), .A2(N5112) );
  NAND2_X1 NAND2_1388( .ZN(N5605), .A1(N3879), .A2(N5113) );
  NAND2_X1 NAND2_1389( .ZN(N5631), .A1(N5324), .A2(N4653) );
  NAND2_X1 NAND2_1390( .ZN(N5632), .A1(N4463), .A2(N5167) );
  NAND2_X1 NAND2_1391( .ZN(N5640), .A1(N4465), .A2(N5168) );
  NAND2_X1 NAND2_1392( .ZN(N5654), .A1(N4467), .A2(N5169) );
  NAND2_X1 NAND2_1393( .ZN(N5670), .A1(N4469), .A2(N5170) );
  NAND2_X1 NAND2_1394( .ZN(N5683), .A1(N4471), .A2(N5171) );
  NAND2_X1 NAND2_1395( .ZN(N5690), .A1(N4475), .A2(N5172) );
  NAND2_X1 NAND2_1396( .ZN(N5697), .A1(N4477), .A2(N5173) );
  NAND2_X1 NAND2_1397( .ZN(N5707), .A1(N4479), .A2(N5174) );
  NAND2_X1 NAND2_1398( .ZN(N5718), .A1(N4481), .A2(N5175) );
  NAND2_X1 NAND2_1399( .ZN(N5728), .A1(N4483), .A2(N5176) );
  INV_X1 NOT1_1400( .ZN(N5735), .A(N5177) );
  NAND2_X1 NAND2_1401( .ZN(N5736), .A1(N5179), .A2(N4490) );
  NAND2_X1 NAND2_1402( .ZN(N5740), .A1(N5180), .A2(N5181) );
  NAND2_X1 NAND2_1403( .ZN(N5744), .A1(N5182), .A2(N5183) );
  NAND2_X1 NAND2_1404( .ZN(N5747), .A1(N5184), .A2(N4496) );
  NAND2_X1 NAND2_1405( .ZN(N5751), .A1(N5185), .A2(N5186) );
  NAND2_X1 NAND2_1406( .ZN(N5755), .A1(N5187), .A2(N5188) );
  NAND2_X1 NAND2_1407( .ZN(N5758), .A1(N5189), .A2(N4502) );
  NAND2_X1 NAND2_1408( .ZN(N5762), .A1(N5190), .A2(N5191) );
  NAND2_X1 NAND2_1409( .ZN(N5766), .A1(N5192), .A2(N5193) );
  INV_X1 NOT1_1410( .ZN(N5769), .A(N4803) );
  INV_X1 NOT1_1411( .ZN(N5770), .A(N4806) );
  NAND2_X1 NAND2_1412( .ZN(N5771), .A1(N4507), .A2(N5196) );
  NAND2_X1 NAND2_1413( .ZN(N5778), .A1(N4509), .A2(N5197) );
  NAND2_X1 NAND2_1414( .ZN(N5789), .A1(N4511), .A2(N5198) );
  NAND2_X1 NAND2_1415( .ZN(N5799), .A1(N4513), .A2(N5199) );
  NAND2_X1 NAND2_1416( .ZN(N5807), .A1(N4515), .A2(N5200) );
  NAND2_X1 NAND2_1417( .ZN(N5821), .A1(N4517), .A2(N5201) );
  NAND2_X1 NAND2_1418( .ZN(N5837), .A1(N4519), .A2(N5202) );
  NAND2_X1 NAND2_1419( .ZN(N5850), .A1(N4521), .A2(N5203) );
  NAND2_X1 NAND2_1420( .ZN(N5856), .A1(N4523), .A2(N5204) );
  NAND2_X1 NAND2_1421( .ZN(N5863), .A1(N4525), .A2(N5205) );
  NAND2_X1 NAND2_1422( .ZN(N5870), .A1(N4527), .A2(N5206) );
  NAND2_X1 NAND2_1423( .ZN(N5881), .A1(N4529), .A2(N5207) );
  NAND2_X1 NAND2_1424( .ZN(N5892), .A1(N4531), .A2(N5208) );
  NAND2_X1 NAND2_1425( .ZN(N5898), .A1(N4533), .A2(N5209) );
  NAND2_X1 NAND2_1426( .ZN(N5905), .A1(N4535), .A2(N5210) );
  NAND2_X2 NAND2_1427( .ZN(N5915), .A1(N4537), .A2(N5211) );
  NAND2_X2 NAND2_1428( .ZN(N5926), .A1(N4539), .A2(N5212) );
  NAND2_X1 NAND2_1429( .ZN(N5936), .A1(N4541), .A2(N5213) );
  INV_X1 NOT1_1430( .ZN(N5943), .A(N4817) );
  NAND2_X1 NAND2_1431( .ZN(N5944), .A1(N4820), .A2(N1931) );
  INV_X1 NOT1_1432( .ZN(N5945), .A(N4820) );
  NAND2_X1 NAND2_1433( .ZN(N5946), .A1(N4823), .A2(N1932) );
  INV_X1 NOT1_1434( .ZN(N5947), .A(N4823) );
  NAND2_X1 NAND2_1435( .ZN(N5948), .A1(N4826), .A2(N1933) );
  INV_X1 NOT1_1436( .ZN(N5949), .A(N4826) );
  NAND2_X1 NAND2_1437( .ZN(N5950), .A1(N4829), .A2(N1934) );
  INV_X1 NOT1_1438( .ZN(N5951), .A(N4829) );
  NAND2_X1 NAND2_1439( .ZN(N5952), .A1(N4832), .A2(N1935) );
  INV_X1 NOT1_1440( .ZN(N5953), .A(N4832) );
  NAND2_X1 NAND2_1441( .ZN(N5954), .A1(N4835), .A2(N1936) );
  INV_X1 NOT1_1442( .ZN(N5955), .A(N4835) );
  NAND2_X1 NAND2_1443( .ZN(N5956), .A1(N4838), .A2(N1937) );
  INV_X1 NOT1_1444( .ZN(N5957), .A(N4838) );
  NAND2_X1 NAND2_1445( .ZN(N5958), .A1(N4841), .A2(N1938) );
  INV_X1 NOT1_1446( .ZN(N5959), .A(N4841) );
  AND2_X1 AND2_1447( .ZN(N5960), .A1(N2674), .A2(N4769) );
  INV_X1 NOT1_1448( .ZN(N5966), .A(N4844) );
  NAND2_X1 NAND2_1449( .ZN(N5967), .A1(N4847), .A2(N1939) );
  INV_X1 NOT1_1450( .ZN(N5968), .A(N4847) );
  NAND2_X1 NAND2_1451( .ZN(N5969), .A1(N4850), .A2(N1940) );
  INV_X1 NOT1_1452( .ZN(N5970), .A(N4850) );
  NAND2_X1 NAND2_1453( .ZN(N5971), .A1(N4853), .A2(N1941) );
  INV_X1 NOT1_1454( .ZN(N5972), .A(N4853) );
  NAND2_X1 NAND2_1455( .ZN(N5973), .A1(N4856), .A2(N1942) );
  INV_X1 NOT1_1456( .ZN(N5974), .A(N4856) );
  NAND2_X1 NAND2_1457( .ZN(N5975), .A1(N4859), .A2(N1943) );
  INV_X1 NOT1_1458( .ZN(N5976), .A(N4859) );
  NAND2_X1 NAND2_1459( .ZN(N5977), .A1(N4862), .A2(N1944) );
  INV_X1 NOT1_1460( .ZN(N5978), .A(N4862) );
  NAND2_X1 NAND2_1461( .ZN(N5979), .A1(N4865), .A2(N1945) );
  INV_X1 NOT1_1462( .ZN(N5980), .A(N4865) );
  AND2_X1 AND2_1463( .ZN(N5981), .A1(N2674), .A2(N4769) );
  NAND2_X1 NAND2_1464( .ZN(N5989), .A1(N4868), .A2(N1946) );
  INV_X1 NOT1_1465( .ZN(N5990), .A(N4868) );
  NAND2_X1 NAND2_1466( .ZN(N5991), .A1(N5283), .A2(N5284) );
  NAND2_X1 NAND2_1467( .ZN(N5996), .A1(N5285), .A2(N5286) );
  NAND2_X1 NAND2_1468( .ZN(N6000), .A1(N5287), .A2(N5288) );
  NAND2_X1 NAND2_1469( .ZN(N6003), .A1(N5289), .A2(N5290) );
  NAND2_X1 NAND2_1470( .ZN(N6009), .A1(N5291), .A2(N5292) );
  NAND2_X1 NAND2_1471( .ZN(N6014), .A1(N5293), .A2(N5294) );
  NAND2_X1 NAND2_1472( .ZN(N6018), .A1(N5295), .A2(N5296) );
  NAND2_X1 NAND2_1473( .ZN(N6021), .A1(N5297), .A2(N5298) );
  NAND2_X1 NAND2_1474( .ZN(N6022), .A1(N5299), .A2(N5300) );
  INV_X1 NOT1_1475( .ZN(N6023), .A(N4874) );
  NAND2_X1 NAND2_1476( .ZN(N6024), .A1(N4874), .A2(N4629) );
  INV_X1 NOT1_1477( .ZN(N6025), .A(N4877) );
  NAND2_X1 NAND2_1478( .ZN(N6026), .A1(N4877), .A2(N4631) );
  INV_X1 NOT1_1479( .ZN(N6027), .A(N4880) );
  NAND2_X1 NAND2_1480( .ZN(N6028), .A1(N4880), .A2(N4633) );
  INV_X1 NOT1_1481( .ZN(N6029), .A(N4883) );
  NAND2_X1 NAND2_1482( .ZN(N6030), .A1(N4883), .A2(N4636) );
  INV_X1 NOT1_1483( .ZN(N6031), .A(N4886) );
  INV_X1 NOT1_1484( .ZN(N6032), .A(N4889) );
  INV_X1 NOT1_1485( .ZN(N6033), .A(N4892) );
  INV_X1 NOT1_1486( .ZN(N6034), .A(N4895) );
  INV_X1 NOT1_1487( .ZN(N6035), .A(N4898) );
  INV_X1 NOT1_1488( .ZN(N6036), .A(N4901) );
  INV_X1 NOT1_1489( .ZN(N6037), .A(N4904) );
  NAND2_X1 NAND2_1490( .ZN(N6038), .A1(N4904), .A2(N4642) );
  INV_X1 NOT1_1491( .ZN(N6039), .A(N4907) );
  INV_X1 NOT1_1492( .ZN(N6040), .A(N4910) );
  NAND2_X1 NAND2_1493( .ZN(N6041), .A1(N5314), .A2(N5315) );
  NAND2_X1 NAND2_1494( .ZN(N6047), .A1(N5316), .A2(N5317) );
  NAND2_X1 NAND2_1495( .ZN(N6052), .A1(N5318), .A2(N5319) );
  NAND2_X1 NAND2_1496( .ZN(N6056), .A1(N5320), .A2(N5321) );
  NAND2_X1 NAND2_1497( .ZN(N6059), .A1(N5322), .A2(N5323) );
  NAND2_X1 NAND2_1498( .ZN(N6060), .A1(N4913), .A2(N1968) );
  INV_X1 NOT1_1499( .ZN(N6061), .A(N4913) );
  NAND2_X1 NAND2_1500( .ZN(N6062), .A1(N4916), .A2(N1969) );
  INV_X1 NOT1_1501( .ZN(N6063), .A(N4916) );
  NAND2_X1 NAND2_1502( .ZN(N6064), .A1(N4919), .A2(N1970) );
  INV_X1 NOT1_1503( .ZN(N6065), .A(N4919) );
  NAND2_X1 NAND2_1504( .ZN(N6066), .A1(N4922), .A2(N1971) );
  INV_X1 NOT1_1505( .ZN(N6067), .A(N4922) );
  NAND2_X1 NAND2_1506( .ZN(N6068), .A1(N4925), .A2(N1972) );
  INV_X1 NOT1_1507( .ZN(N6069), .A(N4925) );
  NAND2_X1 NAND2_1508( .ZN(N6070), .A1(N4928), .A2(N1973) );
  INV_X1 NOT1_1509( .ZN(N6071), .A(N4928) );
  NAND2_X1 NAND2_1510( .ZN(N6072), .A1(N4931), .A2(N1974) );
  INV_X2 NOT1_1511( .ZN(N6073), .A(N4931) );
  NAND2_X1 NAND2_1512( .ZN(N6074), .A1(N4934), .A2(N1975) );
  INV_X1 NOT1_1513( .ZN(N6075), .A(N4934) );
  NAND2_X1 NAND2_1514( .ZN(N6076), .A1(N4937), .A2(N1976) );
  INV_X1 NOT1_1515( .ZN(N6077), .A(N4937) );
  INV_X1 NOT1_1516( .ZN(N6078), .A(N4940) );
  NAND2_X1 NAND2_1517( .ZN(N6079), .A1(N5363), .A2(N4694) );
  NAND2_X1 NAND2_1518( .ZN(N6083), .A1(N5364), .A2(N5365) );
  NAND2_X1 NAND2_1519( .ZN(N6087), .A1(N5366), .A2(N5367) );
  INV_X1 NOT1_1520( .ZN(N6090), .A(N4943) );
  NAND2_X1 NAND2_1521( .ZN(N6091), .A1(N4943), .A2(N4699) );
  INV_X1 NOT1_1522( .ZN(N6092), .A(N4946) );
  INV_X1 NOT1_1523( .ZN(N6093), .A(N4949) );
  INV_X1 NOT1_1524( .ZN(N6094), .A(N4952) );
  INV_X1 NOT1_1525( .ZN(N6095), .A(N4955) );
  INV_X1 NOT1_1526( .ZN(N6096), .A(N4970) );
  NAND2_X1 NAND2_1527( .ZN(N6097), .A1(N4970), .A2(N4700) );
  INV_X1 NOT1_1528( .ZN(N6098), .A(N4973) );
  INV_X1 NOT1_1529( .ZN(N6099), .A(N4976) );
  INV_X1 NOT1_1530( .ZN(N6100), .A(N4979) );
  INV_X1 NOT1_1531( .ZN(N6101), .A(N4982) );
  INV_X1 NOT1_1532( .ZN(N6102), .A(N4997) );
  NAND2_X1 NAND2_1533( .ZN(N6103), .A1(N5000), .A2(N2015) );
  INV_X1 NOT1_1534( .ZN(N6104), .A(N5000) );
  NAND2_X1 NAND2_1535( .ZN(N6105), .A1(N5003), .A2(N2016) );
  INV_X1 NOT1_1536( .ZN(N6106), .A(N5003) );
  NAND2_X1 NAND2_1537( .ZN(N6107), .A1(N5006), .A2(N2017) );
  INV_X1 NOT1_1538( .ZN(N6108), .A(N5006) );
  NAND2_X1 NAND2_1539( .ZN(N6109), .A1(N5009), .A2(N2018) );
  INV_X1 NOT1_1540( .ZN(N6110), .A(N5009) );
  NAND2_X1 NAND2_1541( .ZN(N6111), .A1(N5012), .A2(N2019) );
  INV_X1 NOT1_1542( .ZN(N6112), .A(N5012) );
  NAND2_X1 NAND2_1543( .ZN(N6113), .A1(N5015), .A2(N2020) );
  INV_X1 NOT1_1544( .ZN(N6114), .A(N5015) );
  NAND2_X1 NAND2_1545( .ZN(N6115), .A1(N5018), .A2(N2021) );
  INV_X1 NOT1_1546( .ZN(N6116), .A(N5018) );
  NAND2_X1 NAND2_1547( .ZN(N6117), .A1(N5021), .A2(N2022) );
  INV_X1 NOT1_1548( .ZN(N6118), .A(N5021) );
  NAND2_X1 NAND2_1549( .ZN(N6119), .A1(N5024), .A2(N2023) );
  INV_X1 NOT1_1550( .ZN(N6120), .A(N5024) );
  INV_X1 NOT1_1551( .ZN(N6121), .A(N5033) );
  NAND2_X1 NAND2_1552( .ZN(N6122), .A1(N5033), .A2(N4743) );
  INV_X1 NOT1_1553( .ZN(N6123), .A(N5036) );
  INV_X1 NOT1_1554( .ZN(N6124), .A(N5039) );
  NAND2_X1 NAND2_1555( .ZN(N6125), .A1(N5042), .A2(N4744) );
  INV_X1 NOT1_1556( .ZN(N6126), .A(N5042) );
  NAND2_X1 NAND2_1557( .ZN(N6127), .A1(N5425), .A2(N4746) );
  NAND2_X1 NAND2_1558( .ZN(N6131), .A1(N5426), .A2(N5427) );
  INV_X1 NOT1_1559( .ZN(N6135), .A(N5049) );
  NAND2_X1 NAND2_1560( .ZN(N6136), .A1(N5049), .A2(N4749) );
  NAND2_X1 NAND2_1561( .ZN(N6137), .A1(N5429), .A2(N4751) );
  NAND2_X1 NAND2_1562( .ZN(N6141), .A1(N5430), .A2(N5431) );
  NAND2_X2 NAND2_1563( .ZN(N6145), .A1(N5432), .A2(N5433) );
  INV_X1 NOT1_1564( .ZN(N6148), .A(N5068) );
  INV_X1 NOT1_1565( .ZN(N6149), .A(N5071) );
  INV_X1 NOT1_1566( .ZN(N6150), .A(N5074) );
  INV_X1 NOT1_1567( .ZN(N6151), .A(N5077) );
  INV_X1 NOT1_1568( .ZN(N6152), .A(N5080) );
  INV_X1 NOT1_1569( .ZN(N6153), .A(N5083) );
  INV_X1 NOT1_1570( .ZN(N6154), .A(N5086) );
  INV_X1 NOT1_1571( .ZN(N6155), .A(N5089) );
  INV_X1 NOT1_1572( .ZN(N6156), .A(N5092) );
  NAND2_X1 NAND2_1573( .ZN(N6157), .A1(N5092), .A2(N4761) );
  INV_X1 NOT1_1574( .ZN(N6158), .A(N5095) );
  NAND2_X1 NAND2_1575( .ZN(N6159), .A1(N5095), .A2(N4763) );
  INV_X1 NOT1_1576( .ZN(N6160), .A(N5098) );
  NAND2_X1 NAND2_1577( .ZN(N6161), .A1(N5098), .A2(N4765) );
  INV_X1 NOT1_1578( .ZN(N6162), .A(N5101) );
  INV_X1 NOT1_1579( .ZN(N6163), .A(N5104) );
  NAND2_X1 NAND2_1580( .ZN(N6164), .A1(N5107), .A2(N4768) );
  INV_X1 NOT1_1581( .ZN(N6165), .A(N5107) );
  NAND2_X1 NAND2_1582( .ZN(N6166), .A1(N5451), .A2(N4776) );
  NAND2_X1 NAND2_1583( .ZN(N6170), .A1(N5452), .A2(N5453) );
  NAND2_X1 NAND2_1584( .ZN(N6174), .A1(N5454), .A2(N5455) );
  NAND2_X1 NAND2_1585( .ZN(N6177), .A1(N5456), .A2(N5457) );
  INV_X1 NOT1_1586( .ZN(N6181), .A(N5114) );
  INV_X1 NOT1_1587( .ZN(N6182), .A(N5117) );
  INV_X1 NOT1_1588( .ZN(N6183), .A(N5120) );
  INV_X1 NOT1_1589( .ZN(N6184), .A(N5123) );
  INV_X1 NOT1_1590( .ZN(N6185), .A(N5138) );
  NAND2_X1 NAND2_1591( .ZN(N6186), .A1(N5138), .A2(N4783) );
  INV_X1 NOT1_1592( .ZN(N6187), .A(N5141) );
  INV_X1 NOT1_1593( .ZN(N6188), .A(N5144) );
  INV_X1 NOT1_1594( .ZN(N6189), .A(N5147) );
  INV_X1 NOT1_1595( .ZN(N6190), .A(N5150) );
  INV_X1 NOT1_1596( .ZN(N6191), .A(N4784) );
  NAND2_X1 NAND2_1597( .ZN(N6192), .A1(N4784), .A2(N2230) );
  INV_X1 NOT1_1598( .ZN(N6193), .A(N4790) );
  NAND2_X1 NAND2_1599( .ZN(N6194), .A1(N4790), .A2(N2765) );
  INV_X1 NOT1_1600( .ZN(N6195), .A(N4796) );
  NAND2_X1 NAND2_1601( .ZN(N6196), .A1(N5476), .A2(N5477) );
  NAND2_X1 NAND2_1602( .ZN(N6199), .A1(N5474), .A2(N5475) );
  INV_X1 NOT1_1603( .ZN(N6202), .A(N4810) );
  INV_X1 NOT1_1604( .ZN(N6203), .A(N4814) );
  BUF_X4 BUFF1_1605( .Z(N6204), .A(N4769) );
  BUF_X1 BUFF1_1606( .Z(N6207), .A(N4555) );
  BUF_X1 BUFF1_1607( .Z(N6210), .A(N4769) );
  INV_X2 NOT1_1608( .ZN(N6213), .A(N4871) );
  BUF_X1 BUFF1_1609( .Z(N6214), .A(N4586) );
  NOR2_X2 NOR2_1610( .ZN(N6217), .A1(N2674), .A2(N4769) );
  BUF_X1 BUFF1_1611( .Z(N6220), .A(N4667) );
  INV_X1 NOT1_1612( .ZN(N6223), .A(N4958) );
  INV_X1 NOT1_1613( .ZN(N6224), .A(N4961) );
  INV_X1 NOT1_1614( .ZN(N6225), .A(N4964) );
  INV_X1 NOT1_1615( .ZN(N6226), .A(N4967) );
  INV_X1 NOT1_1616( .ZN(N6227), .A(N4985) );
  INV_X1 NOT1_1617( .ZN(N6228), .A(N4988) );
  INV_X1 NOT1_1618( .ZN(N6229), .A(N4991) );
  INV_X1 NOT1_1619( .ZN(N6230), .A(N4994) );
  INV_X1 NOT1_1620( .ZN(N6231), .A(N5027) );
  BUF_X1 BUFF1_1621( .Z(N6232), .A(N4711) );
  INV_X1 NOT1_1622( .ZN(N6235), .A(N5030) );
  BUF_X1 BUFF1_1623( .Z(N6236), .A(N4735) );
  INV_X1 NOT1_1624( .ZN(N6239), .A(N5052) );
  INV_X1 NOT1_1625( .ZN(N6240), .A(N5055) );
  INV_X1 NOT1_1626( .ZN(N6241), .A(N5058) );
  INV_X1 NOT1_1627( .ZN(N6242), .A(N5061) );
  NAND2_X1 NAND2_1628( .ZN(N6243), .A1(N5573), .A2(N5574) );
  NAND2_X1 NAND2_1629( .ZN(N6246), .A1(N5571), .A2(N5572) );
  NAND2_X1 NAND2_1630( .ZN(N6249), .A1(N5586), .A2(N5587) );
  NAND2_X1 NAND2_1631( .ZN(N6252), .A1(N5584), .A2(N5585) );
  INV_X1 NOT1_1632( .ZN(N6255), .A(N5126) );
  INV_X1 NOT1_1633( .ZN(N6256), .A(N5129) );
  INV_X1 NOT1_1634( .ZN(N6257), .A(N5132) );
  INV_X1 NOT1_1635( .ZN(N6258), .A(N5135) );
  INV_X1 NOT1_1636( .ZN(N6259), .A(N5153) );
  INV_X1 NOT1_1637( .ZN(N6260), .A(N5156) );
  INV_X1 NOT1_1638( .ZN(N6261), .A(N5159) );
  INV_X1 NOT1_1639( .ZN(N6262), .A(N5162) );
  NAND2_X1 NAND2_1640( .ZN(N6263), .A1(N5604), .A2(N5605) );
  NAND2_X1 NAND2_1641( .ZN(N6266), .A1(N5602), .A2(N5603) );
  NAND2_X1 NAND2_1642( .ZN(N6540), .A1(N1380), .A2(N5945) );
  NAND2_X1 NAND2_1643( .ZN(N6541), .A1(N1383), .A2(N5947) );
  NAND2_X1 NAND2_1644( .ZN(N6542), .A1(N1386), .A2(N5949) );
  NAND2_X1 NAND2_1645( .ZN(N6543), .A1(N1389), .A2(N5951) );
  NAND2_X1 NAND2_1646( .ZN(N6544), .A1(N1392), .A2(N5953) );
  NAND2_X1 NAND2_1647( .ZN(N6545), .A1(N1395), .A2(N5955) );
  NAND2_X1 NAND2_1648( .ZN(N6546), .A1(N1398), .A2(N5957) );
  NAND2_X1 NAND2_1649( .ZN(N6547), .A1(N1401), .A2(N5959) );
  NAND2_X1 NAND2_1650( .ZN(N6555), .A1(N1404), .A2(N5968) );
  NAND2_X1 NAND2_1651( .ZN(N6556), .A1(N1407), .A2(N5970) );
  NAND2_X1 NAND2_1652( .ZN(N6557), .A1(N1410), .A2(N5972) );
  NAND2_X1 NAND2_1653( .ZN(N6558), .A1(N1413), .A2(N5974) );
  NAND2_X1 NAND2_1654( .ZN(N6559), .A1(N1416), .A2(N5976) );
  NAND2_X1 NAND2_1655( .ZN(N6560), .A1(N1419), .A2(N5978) );
  NAND2_X1 NAND2_1656( .ZN(N6561), .A1(N1422), .A2(N5980) );
  NAND2_X1 NAND2_1657( .ZN(N6569), .A1(N1425), .A2(N5990) );
  NAND2_X1 NAND2_1658( .ZN(N6594), .A1(N3721), .A2(N6023) );
  NAND2_X1 NAND2_1659( .ZN(N6595), .A1(N3724), .A2(N6025) );
  NAND2_X1 NAND2_1660( .ZN(N6596), .A1(N3727), .A2(N6027) );
  NAND2_X1 NAND2_1661( .ZN(N6597), .A1(N3730), .A2(N6029) );
  NAND2_X1 NAND2_1662( .ZN(N6598), .A1(N4889), .A2(N6031) );
  NAND2_X1 NAND2_1663( .ZN(N6599), .A1(N4886), .A2(N6032) );
  NAND2_X1 NAND2_1664( .ZN(N6600), .A1(N4895), .A2(N6033) );
  NAND2_X1 NAND2_1665( .ZN(N6601), .A1(N4892), .A2(N6034) );
  NAND2_X1 NAND2_1666( .ZN(N6602), .A1(N4901), .A2(N6035) );
  NAND2_X1 NAND2_1667( .ZN(N6603), .A1(N4898), .A2(N6036) );
  NAND2_X1 NAND2_1668( .ZN(N6604), .A1(N3733), .A2(N6037) );
  NAND2_X1 NAND2_1669( .ZN(N6605), .A1(N4910), .A2(N6039) );
  NAND2_X1 NAND2_1670( .ZN(N6606), .A1(N4907), .A2(N6040) );
  NAND2_X1 NAND2_1671( .ZN(N6621), .A1(N1434), .A2(N6061) );
  NAND2_X1 NAND2_1672( .ZN(N6622), .A1(N1437), .A2(N6063) );
  NAND2_X1 NAND2_1673( .ZN(N6623), .A1(N1440), .A2(N6065) );
  NAND2_X1 NAND2_1674( .ZN(N6624), .A1(N1443), .A2(N6067) );
  NAND2_X1 NAND2_1675( .ZN(N6625), .A1(N1446), .A2(N6069) );
  NAND2_X1 NAND2_1676( .ZN(N6626), .A1(N1449), .A2(N6071) );
  NAND2_X1 NAND2_1677( .ZN(N6627), .A1(N1452), .A2(N6073) );
  NAND2_X1 NAND2_1678( .ZN(N6628), .A1(N1455), .A2(N6075) );
  NAND2_X1 NAND2_1679( .ZN(N6629), .A1(N1458), .A2(N6077) );
  NAND2_X1 NAND2_1680( .ZN(N6639), .A1(N3783), .A2(N6090) );
  NAND2_X1 NAND2_1681( .ZN(N6640), .A1(N4949), .A2(N6092) );
  NAND2_X1 NAND2_1682( .ZN(N6641), .A1(N4946), .A2(N6093) );
  NAND2_X1 NAND2_1683( .ZN(N6642), .A1(N4955), .A2(N6094) );
  NAND2_X1 NAND2_1684( .ZN(N6643), .A1(N4952), .A2(N6095) );
  NAND2_X1 NAND2_1685( .ZN(N6644), .A1(N3786), .A2(N6096) );
  NAND2_X1 NAND2_1686( .ZN(N6645), .A1(N4976), .A2(N6098) );
  NAND2_X1 NAND2_1687( .ZN(N6646), .A1(N4973), .A2(N6099) );
  NAND2_X1 NAND2_1688( .ZN(N6647), .A1(N4982), .A2(N6100) );
  NAND2_X1 NAND2_1689( .ZN(N6648), .A1(N4979), .A2(N6101) );
  NAND2_X1 NAND2_1690( .ZN(N6649), .A1(N1461), .A2(N6104) );
  NAND2_X1 NAND2_1691( .ZN(N6650), .A1(N1464), .A2(N6106) );
  NAND2_X1 NAND2_1692( .ZN(N6651), .A1(N1467), .A2(N6108) );
  NAND2_X1 NAND2_1693( .ZN(N6652), .A1(N1470), .A2(N6110) );
  NAND2_X1 NAND2_1694( .ZN(N6653), .A1(N1473), .A2(N6112) );
  NAND2_X1 NAND2_1695( .ZN(N6654), .A1(N1476), .A2(N6114) );
  NAND2_X1 NAND2_1696( .ZN(N6655), .A1(N1479), .A2(N6116) );
  NAND2_X1 NAND2_1697( .ZN(N6656), .A1(N1482), .A2(N6118) );
  NAND2_X1 NAND2_1698( .ZN(N6657), .A1(N1485), .A2(N6120) );
  NAND2_X1 NAND2_1699( .ZN(N6658), .A1(N3789), .A2(N6121) );
  NAND2_X1 NAND2_1700( .ZN(N6659), .A1(N5039), .A2(N6123) );
  NAND2_X1 NAND2_1701( .ZN(N6660), .A1(N5036), .A2(N6124) );
  NAND2_X1 NAND2_1702( .ZN(N6661), .A1(N3792), .A2(N6126) );
  NAND2_X1 NAND2_1703( .ZN(N6668), .A1(N3816), .A2(N6135) );
  NAND2_X1 NAND2_1704( .ZN(N6677), .A1(N5071), .A2(N6148) );
  NAND2_X1 NAND2_1705( .ZN(N6678), .A1(N5068), .A2(N6149) );
  NAND2_X1 NAND2_1706( .ZN(N6679), .A1(N5077), .A2(N6150) );
  NAND2_X1 NAND2_1707( .ZN(N6680), .A1(N5074), .A2(N6151) );
  NAND2_X1 NAND2_1708( .ZN(N6681), .A1(N5083), .A2(N6152) );
  NAND2_X2 NAND2_1709( .ZN(N6682), .A1(N5080), .A2(N6153) );
  NAND2_X2 NAND2_1710( .ZN(N6683), .A1(N5089), .A2(N6154) );
  NAND2_X2 NAND2_1711( .ZN(N6684), .A1(N5086), .A2(N6155) );
  NAND2_X2 NAND2_1712( .ZN(N6685), .A1(N3846), .A2(N6156) );
  NAND2_X2 NAND2_1713( .ZN(N6686), .A1(N3849), .A2(N6158) );
  NAND2_X2 NAND2_1714( .ZN(N6687), .A1(N3852), .A2(N6160) );
  NAND2_X2 NAND2_1715( .ZN(N6688), .A1(N5104), .A2(N6162) );
  NAND2_X2 NAND2_1716( .ZN(N6689), .A1(N5101), .A2(N6163) );
  NAND2_X2 NAND2_1717( .ZN(N6690), .A1(N3855), .A2(N6165) );
  NAND2_X2 NAND2_1718( .ZN(N6702), .A1(N5117), .A2(N6181) );
  NAND2_X2 NAND2_1719( .ZN(N6703), .A1(N5114), .A2(N6182) );
  NAND2_X2 NAND2_1720( .ZN(N6704), .A1(N5123), .A2(N6183) );
  NAND2_X1 NAND2_1721( .ZN(N6705), .A1(N5120), .A2(N6184) );
  NAND2_X1 NAND2_1722( .ZN(N6706), .A1(N3891), .A2(N6185) );
  NAND2_X1 NAND2_1723( .ZN(N6707), .A1(N5144), .A2(N6187) );
  NAND2_X1 NAND2_1724( .ZN(N6708), .A1(N5141), .A2(N6188) );
  NAND2_X1 NAND2_1725( .ZN(N6709), .A1(N5150), .A2(N6189) );
  NAND2_X1 NAND2_1726( .ZN(N6710), .A1(N5147), .A2(N6190) );
  NAND2_X1 NAND2_1727( .ZN(N6711), .A1(N1708), .A2(N6191) );
  NAND2_X1 NAND2_1728( .ZN(N6712), .A1(N2231), .A2(N6193) );
  NAND2_X1 NAND2_1729( .ZN(N6729), .A1(N4961), .A2(N6223) );
  NAND2_X1 NAND2_1730( .ZN(N6730), .A1(N4958), .A2(N6224) );
  NAND2_X1 NAND2_1731( .ZN(N6731), .A1(N4967), .A2(N6225) );
  NAND2_X1 NAND2_1732( .ZN(N6732), .A1(N4964), .A2(N6226) );
  NAND2_X1 NAND2_1733( .ZN(N6733), .A1(N4988), .A2(N6227) );
  NAND2_X1 NAND2_1734( .ZN(N6734), .A1(N4985), .A2(N6228) );
  NAND2_X1 NAND2_1735( .ZN(N6735), .A1(N4994), .A2(N6229) );
  NAND2_X1 NAND2_1736( .ZN(N6736), .A1(N4991), .A2(N6230) );
  NAND2_X1 NAND2_1737( .ZN(N6741), .A1(N5055), .A2(N6239) );
  NAND2_X1 NAND2_1738( .ZN(N6742), .A1(N5052), .A2(N6240) );
  NAND2_X1 NAND2_1739( .ZN(N6743), .A1(N5061), .A2(N6241) );
  NAND2_X1 NAND2_1740( .ZN(N6744), .A1(N5058), .A2(N6242) );
  NAND2_X1 NAND2_1741( .ZN(N6751), .A1(N5129), .A2(N6255) );
  NAND2_X1 NAND2_1742( .ZN(N6752), .A1(N5126), .A2(N6256) );
  NAND2_X1 NAND2_1743( .ZN(N6753), .A1(N5135), .A2(N6257) );
  NAND2_X1 NAND2_1744( .ZN(N6754), .A1(N5132), .A2(N6258) );
  NAND2_X1 NAND2_1745( .ZN(N6755), .A1(N5156), .A2(N6259) );
  NAND2_X1 NAND2_1746( .ZN(N6756), .A1(N5153), .A2(N6260) );
  NAND2_X1 NAND2_1747( .ZN(N6757), .A1(N5162), .A2(N6261) );
  NAND2_X1 NAND2_1748( .ZN(N6758), .A1(N5159), .A2(N6262) );
  INV_X2 NOT1_1749( .ZN(N6761), .A(N5892) );
  AND4_X4 AND5_1750_A( .ZN(extra0), .A1(N5683), .A2(N5670), .A3(N5654), .A4(N5640) );
  AND2_X1 AND5_1750( .ZN(N6762), .A1(extra0), .A2(N5632) );
  AND2_X1 AND2_1751( .ZN(N6766), .A1(N5632), .A2(N3097) );
  AND3_X1 AND3_1752( .ZN(N6767), .A1(N5640), .A2(N5632), .A3(N3101) );
  AND4_X1 AND4_1753( .ZN(N6768), .A1(N5654), .A2(N5632), .A3(N3107), .A4(N5640) );
  AND4_X4 AND5_1754_A( .ZN(extra1), .A1(N5670), .A2(N5654), .A3(N5632), .A4(N3114) );
  AND2_X1 AND5_1754( .ZN(N6769), .A1(extra1), .A2(N5640) );
  AND2_X1 AND2_1755( .ZN(N6770), .A1(N5640), .A2(N3101) );
  AND3_X1 AND3_1756( .ZN(N6771), .A1(N5654), .A2(N3107), .A3(N5640) );
  AND4_X1 AND4_1757( .ZN(N6772), .A1(N5670), .A2(N5654), .A3(N3114), .A4(N5640) );
  AND4_X1 AND4_1758( .ZN(N6773), .A1(N5683), .A2(N5654), .A3(N5640), .A4(N5670) );
  AND2_X1 AND2_1759( .ZN(N6774), .A1(N5640), .A2(N3101) );
  AND3_X1 AND3_1760( .ZN(N6775), .A1(N5654), .A2(N3107), .A3(N5640) );
  AND4_X1 AND4_1761( .ZN(N6776), .A1(N5670), .A2(N5654), .A3(N3114), .A4(N5640) );
  AND2_X1 AND2_1762( .ZN(N6777), .A1(N5654), .A2(N3107) );
  AND3_X1 AND3_1763( .ZN(N6778), .A1(N5670), .A2(N5654), .A3(N3114) );
  AND3_X1 AND3_1764( .ZN(N6779), .A1(N5683), .A2(N5654), .A3(N5670) );
  AND2_X1 AND2_1765( .ZN(N6780), .A1(N5654), .A2(N3107) );
  AND3_X1 AND3_1766( .ZN(N6781), .A1(N5670), .A2(N5654), .A3(N3114) );
  AND2_X1 AND2_1767( .ZN(N6782), .A1(N5670), .A2(N3114) );
  AND2_X1 AND2_1768( .ZN(N6783), .A1(N5683), .A2(N5670) );
  AND4_X4 AND5_1769_A( .ZN(extra2), .A1(N5697), .A2(N5728), .A3(N5707), .A4(N5690) );
  AND2_X1 AND5_1769( .ZN(N6784), .A1(extra2), .A2(N5718) );
  AND2_X1 AND2_1770( .ZN(N6787), .A1(N5690), .A2(N3137) );
  AND3_X1 AND3_1771( .ZN(N6788), .A1(N5697), .A2(N5690), .A3(N3140) );
  AND4_X1 AND4_1772( .ZN(N6789), .A1(N5707), .A2(N5690), .A3(N3144), .A4(N5697) );
  AND4_X4 AND5_1773_A( .ZN(extra3), .A1(N5718), .A2(N5707), .A3(N5690), .A4(N3149) );
  AND2_X1 AND5_1773( .ZN(N6790), .A1(extra3), .A2(N5697) );
  AND2_X1 AND2_1774( .ZN(N6791), .A1(N5697), .A2(N3140) );
  AND3_X1 AND3_1775( .ZN(N6792), .A1(N5707), .A2(N3144), .A3(N5697) );
  AND4_X4 AND4_1776( .ZN(N6793), .A1(N5718), .A2(N5707), .A3(N3149), .A4(N5697) );
  AND2_X1 AND2_1777( .ZN(N6794), .A1(N3144), .A2(N5707) );
  AND3_X1 AND3_1778( .ZN(N6795), .A1(N5718), .A2(N5707), .A3(N3149) );
  AND2_X1 AND2_1779( .ZN(N6796), .A1(N5718), .A2(N3149) );
  INV_X1 NOT1_1780( .ZN(N6797), .A(N5736) );
  INV_X1 NOT1_1781( .ZN(N6800), .A(N5740) );
  INV_X1 NOT1_1782( .ZN(N6803), .A(N5747) );
  INV_X1 NOT1_1783( .ZN(N6806), .A(N5751) );
  INV_X1 NOT1_1784( .ZN(N6809), .A(N5758) );
  INV_X1 NOT1_1785( .ZN(N6812), .A(N5762) );
  BUF_X4 BUFF1_1786( .Z(N6815), .A(N5744) );
  BUF_X1 BUFF1_1787( .Z(N6818), .A(N5744) );
  BUF_X1 BUFF1_1788( .Z(N6821), .A(N5755) );
  BUF_X1 BUFF1_1789( .Z(N6824), .A(N5755) );
  BUF_X1 BUFF1_1790( .Z(N6827), .A(N5766) );
  BUF_X1 BUFF1_1791( .Z(N6830), .A(N5766) );
  AND4_X1 AND4_1792( .ZN(N6833), .A1(N5850), .A2(N5789), .A3(N5778), .A4(N5771) );
  AND2_X1 AND2_1793( .ZN(N6836), .A1(N5771), .A2(N3169) );
  AND3_X1 AND3_1794( .ZN(N6837), .A1(N5778), .A2(N5771), .A3(N3173) );
  AND4_X4 AND4_1795( .ZN(N6838), .A1(N5789), .A2(N5771), .A3(N3178), .A4(N5778) );
  AND2_X1 AND2_1796( .ZN(N6839), .A1(N5778), .A2(N3173) );
  AND3_X1 AND3_1797( .ZN(N6840), .A1(N5789), .A2(N3178), .A3(N5778) );
  AND3_X1 AND3_1798( .ZN(N6841), .A1(N5850), .A2(N5789), .A3(N5778) );
  AND2_X1 AND2_1799( .ZN(N6842), .A1(N5778), .A2(N3173) );
  AND3_X1 AND3_1800( .ZN(N6843), .A1(N5789), .A2(N3178), .A3(N5778) );
  AND2_X1 AND2_1801( .ZN(N6844), .A1(N5789), .A2(N3178) );
  AND4_X1 AND5_1802_A( .ZN(extra4), .A1(N5856), .A2(N5837), .A3(N5821), .A4(N5807) );
  AND2_X1 AND5_1802( .ZN(N6845), .A1(extra4), .A2(N5799) );
  AND2_X1 AND2_1803( .ZN(N6848), .A1(N5799), .A2(N3185) );
  AND3_X1 AND3_1804( .ZN(N6849), .A1(N5807), .A2(N5799), .A3(N3189) );
  AND4_X1 AND4_1805( .ZN(N6850), .A1(N5821), .A2(N5799), .A3(N3195), .A4(N5807) );
  AND4_X4 AND5_1806_A( .ZN(extra5), .A1(N5837), .A2(N5821), .A3(N5799), .A4(N3202) );
  AND2_X1 AND5_1806( .ZN(N6851), .A1(extra5), .A2(N5807) );
  AND2_X1 AND2_1807( .ZN(N6852), .A1(N5807), .A2(N3189) );
  AND3_X1 AND3_1808( .ZN(N6853), .A1(N5821), .A2(N3195), .A3(N5807) );
  AND4_X4 AND4_1809( .ZN(N6854), .A1(N5837), .A2(N5821), .A3(N3202), .A4(N5807) );
  AND4_X1 AND4_1810( .ZN(N6855), .A1(N5856), .A2(N5821), .A3(N5807), .A4(N5837) );
  AND2_X1 AND2_1811( .ZN(N6856), .A1(N5807), .A2(N3189) );
  AND3_X1 AND3_1812( .ZN(N6857), .A1(N5821), .A2(N3195), .A3(N5807) );
  AND4_X1 AND4_1813( .ZN(N6858), .A1(N5837), .A2(N5821), .A3(N3202), .A4(N5807) );
  AND2_X1 AND2_1814( .ZN(N6859), .A1(N5821), .A2(N3195) );
  AND3_X1 AND3_1815( .ZN(N6860), .A1(N5837), .A2(N5821), .A3(N3202) );
  AND3_X1 AND3_1816( .ZN(N6861), .A1(N5856), .A2(N5821), .A3(N5837) );
  AND2_X1 AND2_1817( .ZN(N6862), .A1(N5821), .A2(N3195) );
  AND3_X1 AND3_1818( .ZN(N6863), .A1(N5837), .A2(N5821), .A3(N3202) );
  AND2_X1 AND2_1819( .ZN(N6864), .A1(N5837), .A2(N3202) );
  AND2_X1 AND2_1820( .ZN(N6865), .A1(N5850), .A2(N5789) );
  AND2_X2 AND2_1821( .ZN(N6866), .A1(N5856), .A2(N5837) );
  AND4_X1 AND4_1822( .ZN(N6867), .A1(N5870), .A2(N5892), .A3(N5881), .A4(N5863) );
  AND2_X2 AND2_1823( .ZN(N6870), .A1(N5863), .A2(N3211) );
  AND3_X1 AND3_1824( .ZN(N6871), .A1(N5870), .A2(N5863), .A3(N3215) );
  AND4_X1 AND4_1825( .ZN(N6872), .A1(N5881), .A2(N5863), .A3(N3221), .A4(N5870) );
  AND2_X2 AND2_1826( .ZN(N6873), .A1(N5870), .A2(N3215) );
  AND3_X1 AND3_1827( .ZN(N6874), .A1(N5881), .A2(N3221), .A3(N5870) );
  AND3_X1 AND3_1828( .ZN(N6875), .A1(N5892), .A2(N5881), .A3(N5870) );
  AND2_X2 AND2_1829( .ZN(N6876), .A1(N5870), .A2(N3215) );
  AND3_X1 AND3_1830( .ZN(N6877), .A1(N3221), .A2(N5881), .A3(N5870) );
  AND2_X2 AND2_1831( .ZN(N6878), .A1(N5881), .A2(N3221) );
  AND2_X1 AND2_1832( .ZN(N6879), .A1(N5892), .A2(N5881) );
  AND2_X1 AND2_1833( .ZN(N6880), .A1(N5881), .A2(N3221) );
  AND4_X1 AND5_1834_A( .ZN(extra6), .A1(N5905), .A2(N5936), .A3(N5915), .A4(N5898) );
  AND2_X1 AND5_1834( .ZN(N6881), .A1(extra6), .A2(N5926) );
  AND2_X1 AND2_1835( .ZN(N6884), .A1(N5898), .A2(N3229) );
  AND3_X1 AND3_1836( .ZN(N6885), .A1(N5905), .A2(N5898), .A3(N3232) );
  AND4_X1 AND4_1837( .ZN(N6886), .A1(N5915), .A2(N5898), .A3(N3236), .A4(N5905) );
  AND4_X1 AND5_1838_A( .ZN(extra7), .A1(N5926), .A2(N5915), .A3(N5898), .A4(N3241) );
  AND2_X1 AND5_1838( .ZN(N6887), .A1(extra7), .A2(N5905) );
  AND2_X1 AND2_1839( .ZN(N6888), .A1(N5905), .A2(N3232) );
  AND3_X1 AND3_1840( .ZN(N6889), .A1(N5915), .A2(N3236), .A3(N5905) );
  AND4_X1 AND4_1841( .ZN(N6890), .A1(N5926), .A2(N5915), .A3(N3241), .A4(N5905) );
  AND2_X1 AND2_1842( .ZN(N6891), .A1(N3236), .A2(N5915) );
  AND3_X1 AND3_1843( .ZN(N6892), .A1(N5926), .A2(N5915), .A3(N3241) );
  AND2_X1 AND2_1844( .ZN(N6893), .A1(N5926), .A2(N3241) );
  NAND2_X2 NAND2_1845( .ZN(N6894), .A1(N5944), .A2(N6540) );
  NAND2_X2 NAND2_1846( .ZN(N6901), .A1(N5946), .A2(N6541) );
  NAND2_X2 NAND2_1847( .ZN(N6912), .A1(N5948), .A2(N6542) );
  NAND2_X2 NAND2_1848( .ZN(N6923), .A1(N5950), .A2(N6543) );
  NAND2_X2 NAND2_1849( .ZN(N6929), .A1(N5952), .A2(N6544) );
  NAND2_X2 NAND2_1850( .ZN(N6936), .A1(N5954), .A2(N6545) );
  NAND2_X2 NAND2_1851( .ZN(N6946), .A1(N5956), .A2(N6546) );
  NAND2_X1 NAND2_1852( .ZN(N6957), .A1(N5958), .A2(N6547) );
  NAND2_X1 NAND2_1853( .ZN(N6967), .A1(N6204), .A2(N4575) );
  INV_X2 NOT1_1854( .ZN(N6968), .A(N6204) );
  INV_X1 NOT1_1855( .ZN(N6969), .A(N6207) );
  NAND2_X1 NAND2_1856( .ZN(N6970), .A1(N5967), .A2(N6555) );
  NAND2_X1 NAND2_1857( .ZN(N6977), .A1(N5969), .A2(N6556) );
  NAND2_X1 NAND2_1858( .ZN(N6988), .A1(N5971), .A2(N6557) );
  NAND2_X1 NAND2_1859( .ZN(N6998), .A1(N5973), .A2(N6558) );
  NAND2_X1 NAND2_1860( .ZN(N7006), .A1(N5975), .A2(N6559) );
  NAND2_X1 NAND2_1861( .ZN(N7020), .A1(N5977), .A2(N6560) );
  NAND2_X1 NAND2_1862( .ZN(N7036), .A1(N5979), .A2(N6561) );
  NAND2_X1 NAND2_1863( .ZN(N7049), .A1(N5989), .A2(N6569) );
  NAND2_X1 NAND2_1864( .ZN(N7055), .A1(N6210), .A2(N4610) );
  INV_X1 NOT1_1865( .ZN(N7056), .A(N6210) );
  AND4_X1 AND4_1866( .ZN(N7057), .A1(N6021), .A2(N6000), .A3(N5996), .A4(N5991) );
  AND2_X1 AND2_1867( .ZN(N7060), .A1(N5991), .A2(N3362) );
  AND3_X1 AND3_1868( .ZN(N7061), .A1(N5996), .A2(N5991), .A3(N3363) );
  AND4_X1 AND4_1869( .ZN(N7062), .A1(N6000), .A2(N5991), .A3(N3364), .A4(N5996) );
  AND4_X1 AND5_1870_A( .ZN(extra8), .A1(N6022), .A2(N6018), .A3(N6014), .A4(N6009) );
  AND2_X1 AND5_1870( .ZN(N7063), .A1(extra8), .A2(N6003) );
  AND2_X1 AND2_1871( .ZN(N7064), .A1(N6003), .A2(N3366) );
  AND3_X1 AND3_1872( .ZN(N7065), .A1(N6009), .A2(N6003), .A3(N3367) );
  AND4_X1 AND4_1873( .ZN(N7066), .A1(N6014), .A2(N6003), .A3(N3368), .A4(N6009) );
  AND4_X1 AND5_1874_A( .ZN(extra9), .A1(N6018), .A2(N6014), .A3(N6003), .A4(N3369) );
  AND2_X1 AND5_1874( .ZN(N7067), .A1(extra9), .A2(N6009) );
  NAND2_X1 NAND2_1875( .ZN(N7068), .A1(N6594), .A2(N6024) );
  NAND2_X1 NAND2_1876( .ZN(N7073), .A1(N6595), .A2(N6026) );
  NAND2_X1 NAND2_1877( .ZN(N7077), .A1(N6596), .A2(N6028) );
  NAND2_X1 NAND2_1878( .ZN(N7080), .A1(N6597), .A2(N6030) );
  NAND2_X1 NAND2_1879( .ZN(N7086), .A1(N6598), .A2(N6599) );
  NAND2_X1 NAND2_1880( .ZN(N7091), .A1(N6600), .A2(N6601) );
  NAND2_X1 NAND2_1881( .ZN(N7095), .A1(N6602), .A2(N6603) );
  NAND2_X1 NAND2_1882( .ZN(N7098), .A1(N6604), .A2(N6038) );
  NAND2_X1 NAND2_1883( .ZN(N7099), .A1(N6605), .A2(N6606) );
  AND4_X1 AND5_1884_A( .ZN(extra10), .A1(N6059), .A2(N6056), .A3(N6052), .A4(N6047) );
  AND2_X1 AND5_1884( .ZN(N7100), .A1(extra10), .A2(N6041) );
  AND2_X1 AND2_1885( .ZN(N7103), .A1(N6041), .A2(N3371) );
  AND3_X1 AND3_1886( .ZN(N7104), .A1(N6047), .A2(N6041), .A3(N3372) );
  AND4_X1 AND4_1887( .ZN(N7105), .A1(N6052), .A2(N6041), .A3(N3373), .A4(N6047) );
  AND4_X1 AND5_1888_A( .ZN(extra11), .A1(N6056), .A2(N6052), .A3(N6041), .A4(N3374) );
  AND2_X1 AND5_1888( .ZN(N7106), .A1(extra11), .A2(N6047) );
  NAND2_X1 NAND2_1889( .ZN(N7107), .A1(N6060), .A2(N6621) );
  NAND2_X1 NAND2_1890( .ZN(N7114), .A1(N6062), .A2(N6622) );
  NAND2_X1 NAND2_1891( .ZN(N7125), .A1(N6064), .A2(N6623) );
  NAND2_X1 NAND2_1892( .ZN(N7136), .A1(N6066), .A2(N6624) );
  NAND2_X1 NAND2_1893( .ZN(N7142), .A1(N6068), .A2(N6625) );
  NAND2_X1 NAND2_1894( .ZN(N7149), .A1(N6070), .A2(N6626) );
  NAND2_X1 NAND2_1895( .ZN(N7159), .A1(N6072), .A2(N6627) );
  NAND2_X1 NAND2_1896( .ZN(N7170), .A1(N6074), .A2(N6628) );
  NAND2_X1 NAND2_1897( .ZN(N7180), .A1(N6076), .A2(N6629) );
  INV_X1 NOT1_1898( .ZN(N7187), .A(N6220) );
  INV_X1 NOT1_1899( .ZN(N7188), .A(N6079) );
  INV_X1 NOT1_1900( .ZN(N7191), .A(N6083) );
  NAND2_X1 NAND2_1901( .ZN(N7194), .A1(N6639), .A2(N6091) );
  NAND2_X1 NAND2_1902( .ZN(N7198), .A1(N6640), .A2(N6641) );
  NAND2_X1 NAND2_1903( .ZN(N7202), .A1(N6642), .A2(N6643) );
  NAND2_X1 NAND2_1904( .ZN(N7205), .A1(N6644), .A2(N6097) );
  NAND2_X1 NAND2_1905( .ZN(N7209), .A1(N6645), .A2(N6646) );
  NAND2_X1 NAND2_1906( .ZN(N7213), .A1(N6647), .A2(N6648) );
  BUF_X4 BUFF1_1907( .Z(N7216), .A(N6087) );
  BUF_X4 BUFF1_1908( .Z(N7219), .A(N6087) );
  NAND2_X1 NAND2_1909( .ZN(N7222), .A1(N6103), .A2(N6649) );
  NAND2_X1 NAND2_1910( .ZN(N7229), .A1(N6105), .A2(N6650) );
  NAND2_X1 NAND2_1911( .ZN(N7240), .A1(N6107), .A2(N6651) );
  NAND2_X1 NAND2_1912( .ZN(N7250), .A1(N6109), .A2(N6652) );
  NAND2_X1 NAND2_1913( .ZN(N7258), .A1(N6111), .A2(N6653) );
  NAND2_X1 NAND2_1914( .ZN(N7272), .A1(N6113), .A2(N6654) );
  NAND2_X1 NAND2_1915( .ZN(N7288), .A1(N6115), .A2(N6655) );
  NAND2_X1 NAND2_1916( .ZN(N7301), .A1(N6117), .A2(N6656) );
  NAND2_X1 NAND2_1917( .ZN(N7307), .A1(N6119), .A2(N6657) );
  NAND2_X1 NAND2_1918( .ZN(N7314), .A1(N6658), .A2(N6122) );
  NAND2_X1 NAND2_1919( .ZN(N7318), .A1(N6659), .A2(N6660) );
  NAND2_X1 NAND2_1920( .ZN(N7322), .A1(N6125), .A2(N6661) );
  INV_X1 NOT1_1921( .ZN(N7325), .A(N6127) );
  INV_X1 NOT1_1922( .ZN(N7328), .A(N6131) );
  NAND2_X1 NAND2_1923( .ZN(N7331), .A1(N6668), .A2(N6136) );
  INV_X1 NOT1_1924( .ZN(N7334), .A(N6137) );
  INV_X1 NOT1_1925( .ZN(N7337), .A(N6141) );
  BUF_X1 BUFF1_1926( .Z(N7340), .A(N6145) );
  BUF_X1 BUFF1_1927( .Z(N7343), .A(N6145) );
  NAND2_X1 NAND2_1928( .ZN(N7346), .A1(N6677), .A2(N6678) );
  NAND2_X1 NAND2_1929( .ZN(N7351), .A1(N6679), .A2(N6680) );
  NAND2_X1 NAND2_1930( .ZN(N7355), .A1(N6681), .A2(N6682) );
  NAND2_X1 NAND2_1931( .ZN(N7358), .A1(N6683), .A2(N6684) );
  NAND2_X1 NAND2_1932( .ZN(N7364), .A1(N6685), .A2(N6157) );
  NAND2_X1 NAND2_1933( .ZN(N7369), .A1(N6686), .A2(N6159) );
  NAND2_X1 NAND2_1934( .ZN(N7373), .A1(N6687), .A2(N6161) );
  NAND2_X1 NAND2_1935( .ZN(N7376), .A1(N6688), .A2(N6689) );
  NAND2_X1 NAND2_1936( .ZN(N7377), .A1(N6164), .A2(N6690) );
  INV_X1 NOT1_1937( .ZN(N7378), .A(N6166) );
  INV_X1 NOT1_1938( .ZN(N7381), .A(N6170) );
  INV_X1 NOT1_1939( .ZN(N7384), .A(N6177) );
  NAND2_X1 NAND2_1940( .ZN(N7387), .A1(N6702), .A2(N6703) );
  NAND2_X1 NAND2_1941( .ZN(N7391), .A1(N6704), .A2(N6705) );
  NAND2_X1 NAND2_1942( .ZN(N7394), .A1(N6706), .A2(N6186) );
  NAND2_X1 NAND2_1943( .ZN(N7398), .A1(N6707), .A2(N6708) );
  NAND2_X1 NAND2_1944( .ZN(N7402), .A1(N6709), .A2(N6710) );
  BUF_X1 BUFF1_1945( .Z(N7405), .A(N6174) );
  BUF_X1 BUFF1_1946( .Z(N7408), .A(N6174) );
  BUF_X1 BUFF1_1947( .Z(N7411), .A(N5936) );
  BUF_X1 BUFF1_1948( .Z(N7414), .A(N5898) );
  BUF_X1 BUFF1_1949( .Z(N7417), .A(N5905) );
  BUF_X1 BUFF1_1950( .Z(N7420), .A(N5915) );
  BUF_X1 BUFF1_1951( .Z(N7423), .A(N5926) );
  BUF_X1 BUFF1_1952( .Z(N7426), .A(N5728) );
  BUF_X1 BUFF1_1953( .Z(N7429), .A(N5690) );
  BUF_X1 BUFF1_1954( .Z(N7432), .A(N5697) );
  BUF_X1 BUFF1_1955( .Z(N7435), .A(N5707) );
  BUF_X1 BUFF1_1956( .Z(N7438), .A(N5718) );
  NAND2_X1 NAND2_1957( .ZN(N7441), .A1(N6192), .A2(N6711) );
  NAND2_X1 NAND2_1958( .ZN(N7444), .A1(N6194), .A2(N6712) );
  BUF_X1 BUFF1_1959( .Z(N7447), .A(N5683) );
  BUF_X1 BUFF1_1960( .Z(N7450), .A(N5670) );
  BUF_X1 BUFF1_1961( .Z(N7453), .A(N5632) );
  BUF_X1 BUFF1_1962( .Z(N7456), .A(N5654) );
  BUF_X1 BUFF1_1963( .Z(N7459), .A(N5640) );
  BUF_X1 BUFF1_1964( .Z(N7462), .A(N5640) );
  BUF_X1 BUFF1_1965( .Z(N7465), .A(N5683) );
  BUF_X1 BUFF1_1966( .Z(N7468), .A(N5670) );
  BUF_X1 BUFF1_1967( .Z(N7471), .A(N5632) );
  BUF_X1 BUFF1_1968( .Z(N7474), .A(N5654) );
  INV_X1 NOT1_1969( .ZN(N7477), .A(N6196) );
  INV_X1 NOT1_1970( .ZN(N7478), .A(N6199) );
  BUF_X1 BUFF1_1971( .Z(N7479), .A(N5850) );
  BUF_X1 BUFF1_1972( .Z(N7482), .A(N5789) );
  BUF_X1 BUFF1_1973( .Z(N7485), .A(N5771) );
  BUF_X1 BUFF1_1974( .Z(N7488), .A(N5778) );
  BUF_X1 BUFF1_1975( .Z(N7491), .A(N5850) );
  BUF_X1 BUFF1_1976( .Z(N7494), .A(N5789) );
  BUF_X1 BUFF1_1977( .Z(N7497), .A(N5771) );
  BUF_X1 BUFF1_1978( .Z(N7500), .A(N5778) );
  BUF_X1 BUFF1_1979( .Z(N7503), .A(N5856) );
  BUF_X1 BUFF1_1980( .Z(N7506), .A(N5837) );
  BUF_X1 BUFF1_1981( .Z(N7509), .A(N5799) );
  BUF_X1 BUFF1_1982( .Z(N7512), .A(N5821) );
  BUF_X1 BUFF1_1983( .Z(N7515), .A(N5807) );
  BUF_X1 BUFF1_1984( .Z(N7518), .A(N5807) );
  BUF_X1 BUFF1_1985( .Z(N7521), .A(N5856) );
  BUF_X1 BUFF1_1986( .Z(N7524), .A(N5837) );
  BUF_X1 BUFF1_1987( .Z(N7527), .A(N5799) );
  BUF_X1 BUFF1_1988( .Z(N7530), .A(N5821) );
  BUF_X1 BUFF1_1989( .Z(N7533), .A(N5863) );
  BUF_X1 BUFF1_1990( .Z(N7536), .A(N5863) );
  BUF_X1 BUFF1_1991( .Z(N7539), .A(N5870) );
  BUF_X1 BUFF1_1992( .Z(N7542), .A(N5870) );
  BUF_X1 BUFF1_1993( .Z(N7545), .A(N5881) );
  BUF_X1 BUFF1_1994( .Z(N7548), .A(N5881) );
  INV_X2 NOT1_1995( .ZN(N7551), .A(N6214) );
  INV_X2 NOT1_1996( .ZN(N7552), .A(N6217) );
  BUF_X4 BUFF1_1997( .Z(N7553), .A(N5981) );
  INV_X1 NOT1_1998( .ZN(N7556), .A(N6249) );
  INV_X1 NOT1_1999( .ZN(N7557), .A(N6252) );
  INV_X1 NOT1_2000( .ZN(N7558), .A(N6243) );
  INV_X1 NOT1_2001( .ZN(N7559), .A(N6246) );
  NAND2_X2 NAND2_2002( .ZN(N7560), .A1(N6731), .A2(N6732) );
  NAND2_X2 NAND2_2003( .ZN(N7563), .A1(N6729), .A2(N6730) );
  NAND2_X1 NAND2_2004( .ZN(N7566), .A1(N6735), .A2(N6736) );
  NAND2_X1 NAND2_2005( .ZN(N7569), .A1(N6733), .A2(N6734) );
  INV_X1 NOT1_2006( .ZN(N7572), .A(N6232) );
  INV_X1 NOT1_2007( .ZN(N7573), .A(N6236) );
  NAND2_X1 NAND2_2008( .ZN(N7574), .A1(N6743), .A2(N6744) );
  NAND2_X1 NAND2_2009( .ZN(N7577), .A1(N6741), .A2(N6742) );
  INV_X1 NOT1_2010( .ZN(N7580), .A(N6263) );
  INV_X1 NOT1_2011( .ZN(N7581), .A(N6266) );
  NAND2_X1 NAND2_2012( .ZN(N7582), .A1(N6753), .A2(N6754) );
  NAND2_X1 NAND2_2013( .ZN(N7585), .A1(N6751), .A2(N6752) );
  NAND2_X1 NAND2_2014( .ZN(N7588), .A1(N6757), .A2(N6758) );
  NAND2_X1 NAND2_2015( .ZN(N7591), .A1(N6755), .A2(N6756) );
  OR4_X1 OR5_2016_A( .ZN(extra12), .A1(N3096), .A2(N6766), .A3(N6767), .A4(N6768) );
  OR2_X1 OR5_2016( .ZN(N7609), .A1(extra12), .A2(N6769) );
  OR2_X1 OR2_2017( .ZN(N7613), .A1(N3107), .A2(N6782) );
  OR4_X1 OR5_2018_A( .ZN(extra13), .A1(N3136), .A2(N6787), .A3(N6788), .A4(N6789) );
  OR2_X1 OR5_2018( .ZN(N7620), .A1(extra13), .A2(N6790) );
  OR4_X1 OR4_2019( .ZN(N7649), .A1(N3168), .A2(N6836), .A3(N6837), .A4(N6838) );
  OR2_X1 OR2_2020( .ZN(N7650), .A1(N3173), .A2(N6844) );
  OR4_X1 OR5_2021_A( .ZN(extra14), .A1(N3184), .A2(N6848), .A3(N6849), .A4(N6850) );
  OR2_X1 OR5_2021( .ZN(N7655), .A1(extra14), .A2(N6851) );
  OR2_X1 OR2_2022( .ZN(N7659), .A1(N3195), .A2(N6864) );
  OR4_X4 OR4_2023( .ZN(N7668), .A1(N3210), .A2(N6870), .A3(N6871), .A4(N6872) );
  OR4_X2 OR5_2024_A( .ZN(extra15), .A1(N3228), .A2(N6884), .A3(N6885), .A4(N6886) );
  OR2_X2 OR5_2024( .ZN(N7671), .A1(extra15), .A2(N6887) );
  NAND2_X1 NAND2_2025( .ZN(N7744), .A1(N3661), .A2(N6968) );
  NAND2_X1 NAND2_2026( .ZN(N7822), .A1(N3664), .A2(N7056) );
  OR4_X1 OR4_2027( .ZN(N7825), .A1(N3361), .A2(N7060), .A3(N7061), .A4(N7062) );
  OR4_X1 OR5_2028_A( .ZN(extra16), .A1(N3365), .A2(N7064), .A3(N7065), .A4(N7066) );
  OR2_X1 OR5_2028( .ZN(N7826), .A1(extra16), .A2(N7067) );
  OR4_X1 OR5_2029_A( .ZN(extra17), .A1(N3370), .A2(N7103), .A3(N7104), .A4(N7105) );
  OR2_X1 OR5_2029( .ZN(N7852), .A1(extra17), .A2(N7106) );
  OR4_X1 OR4_2030( .ZN(N8114), .A1(N3101), .A2(N6777), .A3(N6778), .A4(N6779) );
  OR4_X1 OR5_2031_A( .ZN(extra18), .A1(N3097), .A2(N6770), .A3(N6771), .A4(N6772) );
  OR2_X1 OR5_2031( .ZN(N8117), .A1(extra18), .A2(N6773) );
  NOR3_X2 NOR3_2032( .ZN(N8131), .A1(N3101), .A2(N6780), .A3(N6781) );
  NOR3_X2 NOR4_2033_A( .ZN(extra19), .A1(N3097), .A2(N6774), .A3(N6775) );
  NOR2_X1 NOR4_2033( .ZN(N8134), .A1(extra19), .A2(N6776) );
  NAND2_X1 NAND2_2034( .ZN(N8144), .A1(N6199), .A2(N7477) );
  NAND2_X1 NAND2_2035( .ZN(N8145), .A1(N6196), .A2(N7478) );
  OR4_X1 OR4_2036( .ZN(N8146), .A1(N3169), .A2(N6839), .A3(N6840), .A4(N6841) );
  NOR3_X1 NOR3_2037( .ZN(N8156), .A1(N3169), .A2(N6842), .A3(N6843) );
  OR4_X1 OR4_2038( .ZN(N8166), .A1(N3189), .A2(N6859), .A3(N6860), .A4(N6861) );
  OR4_X2 OR5_2039_A( .ZN(extra20), .A1(N3185), .A2(N6852), .A3(N6853), .A4(N6854) );
  OR2_X1 OR5_2039( .ZN(N8169), .A1(extra20), .A2(N6855) );
  NOR3_X1 NOR3_2040( .ZN(N8183), .A1(N3189), .A2(N6862), .A3(N6863) );
  NOR3_X1 NOR4_2041_A( .ZN(extra21), .A1(N3185), .A2(N6856), .A3(N6857) );
  NOR2_X1 NOR4_2041( .ZN(N8186), .A1(extra21), .A2(N6858) );
  OR4_X1 OR4_2042( .ZN(N8196), .A1(N3211), .A2(N6873), .A3(N6874), .A4(N6875) );
  NOR3_X1 NOR3_2043( .ZN(N8200), .A1(N3211), .A2(N6876), .A3(N6877) );
  OR3_X1 OR3_2044( .ZN(N8204), .A1(N3215), .A2(N6878), .A3(N6879) );
  NOR2_X1 NOR2_2045( .ZN(N8208), .A1(N3215), .A2(N6880) );
  NAND2_X1 NAND2_2046( .ZN(N8216), .A1(N6252), .A2(N7556) );
  NAND2_X1 NAND2_2047( .ZN(N8217), .A1(N6249), .A2(N7557) );
  NAND2_X1 NAND2_2048( .ZN(N8218), .A1(N6246), .A2(N7558) );
  NAND2_X1 NAND2_2049( .ZN(N8219), .A1(N6243), .A2(N7559) );
  NAND2_X1 NAND2_2050( .ZN(N8232), .A1(N6266), .A2(N7580) );
  NAND2_X1 NAND2_2051( .ZN(N8233), .A1(N6263), .A2(N7581) );
  INV_X1 NOT1_2052( .ZN(N8242), .A(N7411) );
  INV_X1 NOT1_2053( .ZN(N8243), .A(N7414) );
  INV_X1 NOT1_2054( .ZN(N8244), .A(N7417) );
  INV_X1 NOT1_2055( .ZN(N8245), .A(N7420) );
  INV_X1 NOT1_2056( .ZN(N8246), .A(N7423) );
  INV_X1 NOT1_2057( .ZN(N8247), .A(N7426) );
  INV_X1 NOT1_2058( .ZN(N8248), .A(N7429) );
  INV_X1 NOT1_2059( .ZN(N8249), .A(N7432) );
  INV_X1 NOT1_2060( .ZN(N8250), .A(N7435) );
  INV_X1 NOT1_2061( .ZN(N8251), .A(N7438) );
  INV_X1 NOT1_2062( .ZN(N8252), .A(N7136) );
  INV_X1 NOT1_2063( .ZN(N8253), .A(N6923) );
  INV_X1 NOT1_2064( .ZN(N8254), .A(N6762) );
  INV_X1 NOT1_2065( .ZN(N8260), .A(N7459) );
  INV_X1 NOT1_2066( .ZN(N8261), .A(N7462) );
  AND2_X2 AND2_2067( .ZN(N8262), .A1(N3122), .A2(N6762) );
  AND2_X1 AND2_2068( .ZN(N8269), .A1(N3155), .A2(N6784) );
  INV_X1 NOT1_2069( .ZN(N8274), .A(N6815) );
  INV_X1 NOT1_2070( .ZN(N8275), .A(N6818) );
  INV_X1 NOT1_2071( .ZN(N8276), .A(N6821) );
  INV_X1 NOT1_2072( .ZN(N8277), .A(N6824) );
  INV_X2 NOT1_2073( .ZN(N8278), .A(N6827) );
  INV_X2 NOT1_2074( .ZN(N8279), .A(N6830) );
  AND3_X1 AND3_2075( .ZN(N8280), .A1(N5740), .A2(N5736), .A3(N6815) );
  AND3_X1 AND3_2076( .ZN(N8281), .A1(N6800), .A2(N6797), .A3(N6818) );
  AND3_X1 AND3_2077( .ZN(N8282), .A1(N5751), .A2(N5747), .A3(N6821) );
  AND3_X1 AND3_2078( .ZN(N8283), .A1(N6806), .A2(N6803), .A3(N6824) );
  AND3_X1 AND3_2079( .ZN(N8284), .A1(N5762), .A2(N5758), .A3(N6827) );
  AND3_X1 AND3_2080( .ZN(N8285), .A1(N6812), .A2(N6809), .A3(N6830) );
  INV_X1 NOT1_2081( .ZN(N8288), .A(N6845) );
  INV_X1 NOT1_2082( .ZN(N8294), .A(N7488) );
  INV_X1 NOT1_2083( .ZN(N8295), .A(N7500) );
  INV_X1 NOT1_2084( .ZN(N8296), .A(N7515) );
  INV_X1 NOT1_2085( .ZN(N8297), .A(N7518) );
  AND2_X1 AND2_2086( .ZN(N8298), .A1(N6833), .A2(N6845) );
  AND2_X1 AND2_2087( .ZN(N8307), .A1(N6867), .A2(N6881) );
  INV_X1 NOT1_2088( .ZN(N8315), .A(N7533) );
  INV_X1 NOT1_2089( .ZN(N8317), .A(N7536) );
  INV_X1 NOT1_2090( .ZN(N8319), .A(N7539) );
  INV_X1 NOT1_2091( .ZN(N8321), .A(N7542) );
  NAND2_X1 NAND2_2092( .ZN(N8322), .A1(N7545), .A2(N4543) );
  INV_X1 NOT1_2093( .ZN(N8323), .A(N7545) );
  NAND2_X1 NAND2_2094( .ZN(N8324), .A1(N7548), .A2(N5943) );
  INV_X1 NOT1_2095( .ZN(N8325), .A(N7548) );
  NAND2_X1 NAND2_2096( .ZN(N8326), .A1(N6967), .A2(N7744) );
  AND4_X1 AND4_2097( .ZN(N8333), .A1(N6901), .A2(N6923), .A3(N6912), .A4(N6894) );
  AND2_X1 AND2_2098( .ZN(N8337), .A1(N6894), .A2(N4545) );
  AND3_X1 AND3_2099( .ZN(N8338), .A1(N6901), .A2(N6894), .A3(N4549) );
  AND4_X1 AND4_2100( .ZN(N8339), .A1(N6912), .A2(N6894), .A3(N4555), .A4(N6901) );
  AND2_X1 AND2_2101( .ZN(N8340), .A1(N6901), .A2(N4549) );
  AND3_X1 AND3_2102( .ZN(N8341), .A1(N6912), .A2(N4555), .A3(N6901) );
  AND3_X1 AND3_2103( .ZN(N8342), .A1(N6923), .A2(N6912), .A3(N6901) );
  AND2_X1 AND2_2104( .ZN(N8343), .A1(N6901), .A2(N4549) );
  AND3_X1 AND3_2105( .ZN(N8344), .A1(N4555), .A2(N6912), .A3(N6901) );
  AND2_X1 AND2_2106( .ZN(N8345), .A1(N6912), .A2(N4555) );
  AND2_X1 AND2_2107( .ZN(N8346), .A1(N6923), .A2(N6912) );
  AND2_X1 AND2_2108( .ZN(N8347), .A1(N6912), .A2(N4555) );
  AND2_X1 AND2_2109( .ZN(N8348), .A1(N6929), .A2(N4563) );
  AND3_X1 AND3_2110( .ZN(N8349), .A1(N6936), .A2(N6929), .A3(N4566) );
  AND4_X1 AND4_2111( .ZN(N8350), .A1(N6946), .A2(N6929), .A3(N4570), .A4(N6936) );
  AND4_X1 AND5_2112_A( .ZN(extra22), .A1(N6957), .A2(N6946), .A3(N6929), .A4(N5960) );
  AND2_X1 AND5_2112( .ZN(N8351), .A1(extra22), .A2(N6936) );
  AND2_X1 AND2_2113( .ZN(N8352), .A1(N6936), .A2(N4566) );
  AND3_X1 AND3_2114( .ZN(N8353), .A1(N6946), .A2(N4570), .A3(N6936) );
  AND4_X1 AND4_2115( .ZN(N8354), .A1(N6957), .A2(N6946), .A3(N5960), .A4(N6936) );
  AND2_X1 AND2_2116( .ZN(N8355), .A1(N4570), .A2(N6946) );
  AND3_X1 AND3_2117( .ZN(N8356), .A1(N6957), .A2(N6946), .A3(N5960) );
  AND2_X1 AND2_2118( .ZN(N8357), .A1(N6957), .A2(N5960) );
  NAND2_X1 NAND2_2119( .ZN(N8358), .A1(N7055), .A2(N7822) );
  AND4_X1 AND4_2120( .ZN(N8365), .A1(N7049), .A2(N6988), .A3(N6977), .A4(N6970) );
  AND2_X1 AND2_2121( .ZN(N8369), .A1(N6970), .A2(N4577) );
  AND3_X1 AND3_2122( .ZN(N8370), .A1(N6977), .A2(N6970), .A3(N4581) );
  AND4_X1 AND4_2123( .ZN(N8371), .A1(N6988), .A2(N6970), .A3(N4586), .A4(N6977) );
  AND2_X1 AND2_2124( .ZN(N8372), .A1(N6977), .A2(N4581) );
  AND3_X1 AND3_2125( .ZN(N8373), .A1(N6988), .A2(N4586), .A3(N6977) );
  AND3_X1 AND3_2126( .ZN(N8374), .A1(N7049), .A2(N6988), .A3(N6977) );
  AND2_X1 AND2_2127( .ZN(N8375), .A1(N6977), .A2(N4581) );
  AND3_X1 AND3_2128( .ZN(N8376), .A1(N6988), .A2(N4586), .A3(N6977) );
  AND2_X1 AND2_2129( .ZN(N8377), .A1(N6988), .A2(N4586) );
  AND2_X1 AND2_2130( .ZN(N8378), .A1(N6998), .A2(N4593) );
  AND3_X1 AND3_2131( .ZN(N8379), .A1(N7006), .A2(N6998), .A3(N4597) );
  AND4_X1 AND4_2132( .ZN(N8380), .A1(N7020), .A2(N6998), .A3(N4603), .A4(N7006) );
  AND4_X1 AND5_2133_A( .ZN(extra23), .A1(N7036), .A2(N7020), .A3(N6998), .A4(N5981) );
  AND2_X1 AND5_2133( .ZN(N8381), .A1(extra23), .A2(N7006) );
  AND2_X1 AND2_2134( .ZN(N8382), .A1(N7006), .A2(N4597) );
  AND3_X1 AND3_2135( .ZN(N8383), .A1(N7020), .A2(N4603), .A3(N7006) );
  AND4_X1 AND4_2136( .ZN(N8384), .A1(N7036), .A2(N7020), .A3(N5981), .A4(N7006) );
  AND2_X1 AND2_2137( .ZN(N8385), .A1(N7006), .A2(N4597) );
  AND3_X1 AND3_2138( .ZN(N8386), .A1(N7020), .A2(N4603), .A3(N7006) );
  AND4_X1 AND4_2139( .ZN(N8387), .A1(N7036), .A2(N7020), .A3(N5981), .A4(N7006) );
  AND2_X1 AND2_2140( .ZN(N8388), .A1(N7020), .A2(N4603) );
  AND3_X1 AND3_2141( .ZN(N8389), .A1(N7036), .A2(N7020), .A3(N5981) );
  AND2_X1 AND2_2142( .ZN(N8390), .A1(N7020), .A2(N4603) );
  AND3_X1 AND3_2143( .ZN(N8391), .A1(N7036), .A2(N7020), .A3(N5981) );
  AND2_X1 AND2_2144( .ZN(N8392), .A1(N7036), .A2(N5981) );
  AND2_X1 AND2_2145( .ZN(N8393), .A1(N7049), .A2(N6988) );
  AND2_X1 AND2_2146( .ZN(N8394), .A1(N7057), .A2(N7063) );
  AND2_X1 AND2_2147( .ZN(N8404), .A1(N7057), .A2(N7826) );
  AND4_X1 AND4_2148( .ZN(N8405), .A1(N7098), .A2(N7077), .A3(N7073), .A4(N7068) );
  AND2_X1 AND2_2149( .ZN(N8409), .A1(N7068), .A2(N4632) );
  AND3_X1 AND3_2150( .ZN(N8410), .A1(N7073), .A2(N7068), .A3(N4634) );
  AND4_X1 AND4_2151( .ZN(N8411), .A1(N7077), .A2(N7068), .A3(N4635), .A4(N7073) );
  AND4_X1 AND5_2152_A( .ZN(extra24), .A1(N7099), .A2(N7095), .A3(N7091), .A4(N7086) );
  AND2_X1 AND5_2152( .ZN(N8412), .A1(extra24), .A2(N7080) );
  AND2_X1 AND2_2153( .ZN(N8415), .A1(N7080), .A2(N4638) );
  AND3_X1 AND3_2154( .ZN(N8416), .A1(N7086), .A2(N7080), .A3(N4639) );
  AND4_X1 AND4_2155( .ZN(N8417), .A1(N7091), .A2(N7080), .A3(N4640), .A4(N7086) );
  AND4_X1 AND5_2156_A( .ZN(extra25), .A1(N7095), .A2(N7091), .A3(N7080), .A4(N4641) );
  AND2_X1 AND5_2156( .ZN(N8418), .A1(extra25), .A2(N7086) );
  AND2_X1 AND2_2157( .ZN(N8421), .A1(N3375), .A2(N7100) );
  AND4_X1 AND4_2158( .ZN(N8430), .A1(N7114), .A2(N7136), .A3(N7125), .A4(N7107) );
  AND2_X1 AND2_2159( .ZN(N8433), .A1(N7107), .A2(N4657) );
  AND3_X1 AND3_2160( .ZN(N8434), .A1(N7114), .A2(N7107), .A3(N4661) );
  AND4_X1 AND4_2161( .ZN(N8435), .A1(N7125), .A2(N7107), .A3(N4667), .A4(N7114) );
  AND2_X1 AND2_2162( .ZN(N8436), .A1(N7114), .A2(N4661) );
  AND3_X1 AND3_2163( .ZN(N8437), .A1(N7125), .A2(N4667), .A3(N7114) );
  AND3_X1 AND3_2164( .ZN(N8438), .A1(N7136), .A2(N7125), .A3(N7114) );
  AND2_X1 AND2_2165( .ZN(N8439), .A1(N7114), .A2(N4661) );
  AND3_X1 AND3_2166( .ZN(N8440), .A1(N4667), .A2(N7125), .A3(N7114) );
  AND2_X1 AND2_2167( .ZN(N8441), .A1(N7125), .A2(N4667) );
  AND2_X1 AND2_2168( .ZN(N8442), .A1(N7136), .A2(N7125) );
  AND2_X1 AND2_2169( .ZN(N8443), .A1(N7125), .A2(N4667) );
  AND4_X1 AND5_2170_A( .ZN(extra26), .A1(N7149), .A2(N7180), .A3(N7159), .A4(N7142) );
  AND2_X1 AND5_2170( .ZN(N8444), .A1(extra26), .A2(N7170) );
  AND2_X1 AND2_2171( .ZN(N8447), .A1(N7142), .A2(N4675) );
  AND3_X1 AND3_2172( .ZN(N8448), .A1(N7149), .A2(N7142), .A3(N4678) );
  AND4_X1 AND4_2173( .ZN(N8449), .A1(N7159), .A2(N7142), .A3(N4682), .A4(N7149) );
  AND4_X1 AND5_2174_A( .ZN(extra27), .A1(N7170), .A2(N7159), .A3(N7142), .A4(N4687) );
  AND2_X1 AND5_2174( .ZN(N8450), .A1(extra27), .A2(N7149) );
  AND2_X1 AND2_2175( .ZN(N8451), .A1(N7149), .A2(N4678) );
  AND3_X1 AND3_2176( .ZN(N8452), .A1(N7159), .A2(N4682), .A3(N7149) );
  AND4_X1 AND4_2177( .ZN(N8453), .A1(N7170), .A2(N7159), .A3(N4687), .A4(N7149) );
  AND2_X1 AND2_2178( .ZN(N8454), .A1(N4682), .A2(N7159) );
  AND3_X1 AND3_2179( .ZN(N8455), .A1(N7170), .A2(N7159), .A3(N4687) );
  AND2_X1 AND2_2180( .ZN(N8456), .A1(N7170), .A2(N4687) );
  INV_X2 NOT1_2181( .ZN(N8457), .A(N7194) );
  INV_X2 NOT1_2182( .ZN(N8460), .A(N7198) );
  INV_X1 NOT1_2183( .ZN(N8463), .A(N7205) );
  INV_X1 NOT1_2184( .ZN(N8466), .A(N7209) );
  INV_X1 NOT1_2185( .ZN(N8469), .A(N7216) );
  INV_X1 NOT1_2186( .ZN(N8470), .A(N7219) );
  BUF_X4 BUFF1_2187( .Z(N8471), .A(N7202) );
  BUF_X4 BUFF1_2188( .Z(N8474), .A(N7202) );
  BUF_X1 BUFF1_2189( .Z(N8477), .A(N7213) );
  BUF_X1 BUFF1_2190( .Z(N8480), .A(N7213) );
  AND3_X1 AND3_2191( .ZN(N8483), .A1(N6083), .A2(N6079), .A3(N7216) );
  AND3_X1 AND3_2192( .ZN(N8484), .A1(N7191), .A2(N7188), .A3(N7219) );
  AND4_X1 AND4_2193( .ZN(N8485), .A1(N7301), .A2(N7240), .A3(N7229), .A4(N7222) );
  AND2_X1 AND2_2194( .ZN(N8488), .A1(N7222), .A2(N4702) );
  AND3_X1 AND3_2195( .ZN(N8489), .A1(N7229), .A2(N7222), .A3(N4706) );
  AND4_X1 AND4_2196( .ZN(N8490), .A1(N7240), .A2(N7222), .A3(N4711), .A4(N7229) );
  AND2_X1 AND2_2197( .ZN(N8491), .A1(N7229), .A2(N4706) );
  AND3_X1 AND3_2198( .ZN(N8492), .A1(N7240), .A2(N4711), .A3(N7229) );
  AND3_X1 AND3_2199( .ZN(N8493), .A1(N7301), .A2(N7240), .A3(N7229) );
  AND2_X2 AND2_2200( .ZN(N8494), .A1(N7229), .A2(N4706) );
  AND3_X1 AND3_2201( .ZN(N8495), .A1(N7240), .A2(N4711), .A3(N7229) );
  AND2_X2 AND2_2202( .ZN(N8496), .A1(N7240), .A2(N4711) );
  AND4_X1 AND5_2203_A( .ZN(extra28), .A1(N7307), .A2(N7288), .A3(N7272), .A4(N7258) );
  AND2_X2 AND5_2203( .ZN(N8497), .A1(extra28), .A2(N7250) );
  AND2_X2 AND2_2204( .ZN(N8500), .A1(N7250), .A2(N4718) );
  AND3_X1 AND3_2205( .ZN(N8501), .A1(N7258), .A2(N7250), .A3(N4722) );
  AND4_X1 AND4_2206( .ZN(N8502), .A1(N7272), .A2(N7250), .A3(N4728), .A4(N7258) );
  AND4_X1 AND5_2207_A( .ZN(extra29), .A1(N7288), .A2(N7272), .A3(N7250), .A4(N4735) );
  AND2_X2 AND5_2207( .ZN(N8503), .A1(extra29), .A2(N7258) );
  AND2_X2 AND2_2208( .ZN(N8504), .A1(N7258), .A2(N4722) );
  AND3_X1 AND3_2209( .ZN(N8505), .A1(N7272), .A2(N4728), .A3(N7258) );
  AND4_X1 AND4_2210( .ZN(N8506), .A1(N7288), .A2(N7272), .A3(N4735), .A4(N7258) );
  AND4_X1 AND4_2211( .ZN(N8507), .A1(N7307), .A2(N7272), .A3(N7258), .A4(N7288) );
  AND2_X2 AND2_2212( .ZN(N8508), .A1(N7258), .A2(N4722) );
  AND3_X1 AND3_2213( .ZN(N8509), .A1(N7272), .A2(N4728), .A3(N7258) );
  AND4_X1 AND4_2214( .ZN(N8510), .A1(N7288), .A2(N7272), .A3(N4735), .A4(N7258) );
  AND2_X2 AND2_2215( .ZN(N8511), .A1(N7272), .A2(N4728) );
  AND3_X1 AND3_2216( .ZN(N8512), .A1(N7288), .A2(N7272), .A3(N4735) );
  AND3_X1 AND3_2217( .ZN(N8513), .A1(N7307), .A2(N7272), .A3(N7288) );
  AND2_X1 AND2_2218( .ZN(N8514), .A1(N7272), .A2(N4728) );
  AND3_X1 AND3_2219( .ZN(N8515), .A1(N7288), .A2(N7272), .A3(N4735) );
  AND2_X1 AND2_2220( .ZN(N8516), .A1(N7288), .A2(N4735) );
  AND2_X1 AND2_2221( .ZN(N8517), .A1(N7301), .A2(N7240) );
  AND2_X1 AND2_2222( .ZN(N8518), .A1(N7307), .A2(N7288) );
  INV_X1 NOT1_2223( .ZN(N8519), .A(N7314) );
  INV_X1 NOT1_2224( .ZN(N8522), .A(N7318) );
  BUF_X1 BUFF1_2225( .Z(N8525), .A(N7322) );
  BUF_X1 BUFF1_2226( .Z(N8528), .A(N7322) );
  BUF_X1 BUFF1_2227( .Z(N8531), .A(N7331) );
  BUF_X1 BUFF1_2228( .Z(N8534), .A(N7331) );
  INV_X1 NOT1_2229( .ZN(N8537), .A(N7340) );
  INV_X1 NOT1_2230( .ZN(N8538), .A(N7343) );
  AND3_X1 AND3_2231( .ZN(N8539), .A1(N6141), .A2(N6137), .A3(N7340) );
  AND3_X1 AND3_2232( .ZN(N8540), .A1(N7337), .A2(N7334), .A3(N7343) );
  AND4_X1 AND4_2233( .ZN(N8541), .A1(N7376), .A2(N7355), .A3(N7351), .A4(N7346) );
  AND2_X1 AND2_2234( .ZN(N8545), .A1(N7346), .A2(N4757) );
  AND3_X1 AND3_2235( .ZN(N8546), .A1(N7351), .A2(N7346), .A3(N4758) );
  AND4_X1 AND4_2236( .ZN(N8547), .A1(N7355), .A2(N7346), .A3(N4759), .A4(N7351) );
  AND4_X1 AND5_2237_A( .ZN(extra30), .A1(N7377), .A2(N7373), .A3(N7369), .A4(N7364) );
  AND2_X1 AND5_2237( .ZN(N8548), .A1(extra30), .A2(N7358) );
  AND2_X1 AND2_2238( .ZN(N8551), .A1(N7358), .A2(N4762) );
  AND3_X1 AND3_2239( .ZN(N8552), .A1(N7364), .A2(N7358), .A3(N4764) );
  AND4_X1 AND4_2240( .ZN(N8553), .A1(N7369), .A2(N7358), .A3(N4766), .A4(N7364) );
  AND4_X1 AND5_2241_A( .ZN(extra31), .A1(N7373), .A2(N7369), .A3(N7358), .A4(N4767) );
  AND2_X1 AND5_2241( .ZN(N8554), .A1(extra31), .A2(N7364) );
  INV_X1 NOT1_2242( .ZN(N8555), .A(N7387) );
  INV_X1 NOT1_2243( .ZN(N8558), .A(N7394) );
  INV_X1 NOT1_2244( .ZN(N8561), .A(N7398) );
  INV_X1 NOT1_2245( .ZN(N8564), .A(N7405) );
  INV_X1 NOT1_2246( .ZN(N8565), .A(N7408) );
  BUF_X1 BUFF1_2247( .Z(N8566), .A(N7391) );
  BUF_X1 BUFF1_2248( .Z(N8569), .A(N7391) );
  BUF_X1 BUFF1_2249( .Z(N8572), .A(N7402) );
  BUF_X1 BUFF1_2250( .Z(N8575), .A(N7402) );
  AND3_X1 AND3_2251( .ZN(N8578), .A1(N6170), .A2(N6166), .A3(N7405) );
  AND3_X1 AND3_2252( .ZN(N8579), .A1(N7381), .A2(N7378), .A3(N7408) );
  BUF_X1 BUFF1_2253( .Z(N8580), .A(N7180) );
  BUF_X1 BUFF1_2254( .Z(N8583), .A(N7142) );
  BUF_X1 BUFF1_2255( .Z(N8586), .A(N7149) );
  BUF_X1 BUFF1_2256( .Z(N8589), .A(N7159) );
  BUF_X1 BUFF1_2257( .Z(N8592), .A(N7170) );
  BUF_X1 BUFF1_2258( .Z(N8595), .A(N6929) );
  BUF_X1 BUFF1_2259( .Z(N8598), .A(N6936) );
  BUF_X1 BUFF1_2260( .Z(N8601), .A(N6946) );
  BUF_X1 BUFF1_2261( .Z(N8604), .A(N6957) );
  INV_X2 NOT1_2262( .ZN(N8607), .A(N7441) );
  NAND2_X2 NAND2_2263( .ZN(N8608), .A1(N7441), .A2(N5469) );
  INV_X2 NOT1_2264( .ZN(N8609), .A(N7444) );
  NAND2_X2 NAND2_2265( .ZN(N8610), .A1(N7444), .A2(N4793) );
  INV_X1 NOT1_2266( .ZN(N8615), .A(N7447) );
  INV_X1 NOT1_2267( .ZN(N8616), .A(N7450) );
  INV_X1 NOT1_2268( .ZN(N8617), .A(N7453) );
  INV_X1 NOT1_2269( .ZN(N8618), .A(N7456) );
  INV_X1 NOT1_2270( .ZN(N8619), .A(N7474) );
  INV_X1 NOT1_2271( .ZN(N8624), .A(N7465) );
  INV_X1 NOT1_2272( .ZN(N8625), .A(N7468) );
  INV_X1 NOT1_2273( .ZN(N8626), .A(N7471) );
  NAND2_X1 NAND2_2274( .ZN(N8627), .A1(N8144), .A2(N8145) );
  INV_X1 NOT1_2275( .ZN(N8632), .A(N7479) );
  INV_X1 NOT1_2276( .ZN(N8633), .A(N7482) );
  INV_X1 NOT1_2277( .ZN(N8634), .A(N7485) );
  INV_X1 NOT1_2278( .ZN(N8637), .A(N7491) );
  INV_X1 NOT1_2279( .ZN(N8638), .A(N7494) );
  INV_X1 NOT1_2280( .ZN(N8639), .A(N7497) );
  INV_X1 NOT1_2281( .ZN(N8644), .A(N7503) );
  INV_X1 NOT1_2282( .ZN(N8645), .A(N7506) );
  INV_X1 NOT1_2283( .ZN(N8646), .A(N7509) );
  INV_X1 NOT1_2284( .ZN(N8647), .A(N7512) );
  INV_X1 NOT1_2285( .ZN(N8648), .A(N7530) );
  INV_X1 NOT1_2286( .ZN(N8653), .A(N7521) );
  INV_X1 NOT1_2287( .ZN(N8654), .A(N7524) );
  INV_X1 NOT1_2288( .ZN(N8655), .A(N7527) );
  BUF_X4 BUFF1_2289( .Z(N8660), .A(N6894) );
  BUF_X4 BUFF1_2290( .Z(N8663), .A(N6894) );
  BUF_X4 BUFF1_2291( .Z(N8666), .A(N6901) );
  BUF_X4 BUFF1_2292( .Z(N8669), .A(N6901) );
  BUF_X4 BUFF1_2293( .Z(N8672), .A(N6912) );
  BUF_X1 BUFF1_2294( .Z(N8675), .A(N6912) );
  BUF_X1 BUFF1_2295( .Z(N8678), .A(N7049) );
  BUF_X1 BUFF1_2296( .Z(N8681), .A(N6988) );
  BUF_X1 BUFF1_2297( .Z(N8684), .A(N6970) );
  BUF_X1 BUFF1_2298( .Z(N8687), .A(N6977) );
  BUF_X1 BUFF1_2299( .Z(N8690), .A(N7049) );
  BUF_X1 BUFF1_2300( .Z(N8693), .A(N6988) );
  BUF_X1 BUFF1_2301( .Z(N8696), .A(N6970) );
  BUF_X1 BUFF1_2302( .Z(N8699), .A(N6977) );
  BUF_X1 BUFF1_2303( .Z(N8702), .A(N7036) );
  BUF_X1 BUFF1_2304( .Z(N8705), .A(N6998) );
  BUF_X1 BUFF1_2305( .Z(N8708), .A(N7020) );
  BUF_X1 BUFF1_2306( .Z(N8711), .A(N7006) );
  BUF_X1 BUFF1_2307( .Z(N8714), .A(N7006) );
  INV_X1 NOT1_2308( .ZN(N8717), .A(N7553) );
  BUF_X1 BUFF1_2309( .Z(N8718), .A(N7036) );
  BUF_X1 BUFF1_2310( .Z(N8721), .A(N6998) );
  BUF_X1 BUFF1_2311( .Z(N8724), .A(N7020) );
  NAND2_X1 NAND2_2312( .ZN(N8727), .A1(N8216), .A2(N8217) );
  NAND2_X1 NAND2_2313( .ZN(N8730), .A1(N8218), .A2(N8219) );
  INV_X1 NOT1_2314( .ZN(N8733), .A(N7574) );
  INV_X1 NOT1_2315( .ZN(N8734), .A(N7577) );
  BUF_X1 BUFF1_2316( .Z(N8735), .A(N7107) );
  BUF_X1 BUFF1_2317( .Z(N8738), .A(N7107) );
  BUF_X1 BUFF1_2318( .Z(N8741), .A(N7114) );
  BUF_X1 BUFF1_2319( .Z(N8744), .A(N7114) );
  BUF_X1 BUFF1_2320( .Z(N8747), .A(N7125) );
  BUF_X1 BUFF1_2321( .Z(N8750), .A(N7125) );
  INV_X1 NOT1_2322( .ZN(N8753), .A(N7560) );
  INV_X1 NOT1_2323( .ZN(N8754), .A(N7563) );
  INV_X1 NOT1_2324( .ZN(N8755), .A(N7566) );
  INV_X1 NOT1_2325( .ZN(N8756), .A(N7569) );
  BUF_X1 BUFF1_2326( .Z(N8757), .A(N7301) );
  BUF_X1 BUFF1_2327( .Z(N8760), .A(N7240) );
  BUF_X1 BUFF1_2328( .Z(N8763), .A(N7222) );
  BUF_X1 BUFF1_2329( .Z(N8766), .A(N7229) );
  BUF_X1 BUFF1_2330( .Z(N8769), .A(N7301) );
  BUF_X1 BUFF1_2331( .Z(N8772), .A(N7240) );
  BUF_X1 BUFF1_2332( .Z(N8775), .A(N7222) );
  BUF_X1 BUFF1_2333( .Z(N8778), .A(N7229) );
  BUF_X1 BUFF1_2334( .Z(N8781), .A(N7307) );
  BUF_X1 BUFF1_2335( .Z(N8784), .A(N7288) );
  BUF_X1 BUFF1_2336( .Z(N8787), .A(N7250) );
  BUF_X1 BUFF1_2337( .Z(N8790), .A(N7272) );
  BUF_X1 BUFF1_2338( .Z(N8793), .A(N7258) );
  BUF_X1 BUFF1_2339( .Z(N8796), .A(N7258) );
  BUF_X1 BUFF1_2340( .Z(N8799), .A(N7307) );
  BUF_X1 BUFF1_2341( .Z(N8802), .A(N7288) );
  BUF_X1 BUFF1_2342( .Z(N8805), .A(N7250) );
  BUF_X1 BUFF1_2343( .Z(N8808), .A(N7272) );
  NAND2_X1 NAND2_2344( .ZN(N8811), .A1(N8232), .A2(N8233) );
  INV_X1 NOT1_2345( .ZN(N8814), .A(N7588) );
  INV_X1 NOT1_2346( .ZN(N8815), .A(N7591) );
  INV_X1 NOT1_2347( .ZN(N8816), .A(N7582) );
  INV_X1 NOT1_2348( .ZN(N8817), .A(N7585) );
  AND2_X2 AND2_2349( .ZN(N8818), .A1(N7620), .A2(N3155) );
  AND2_X1 AND2_2350( .ZN(N8840), .A1(N3122), .A2(N7609) );
  INV_X1 NOT1_2351( .ZN(N8857), .A(N7609) );
  AND3_X1 AND3_2352( .ZN(N8861), .A1(N6797), .A2(N5740), .A3(N8274) );
  AND3_X1 AND3_2353( .ZN(N8862), .A1(N5736), .A2(N6800), .A3(N8275) );
  AND3_X1 AND3_2354( .ZN(N8863), .A1(N6803), .A2(N5751), .A3(N8276) );
  AND3_X1 AND3_2355( .ZN(N8864), .A1(N5747), .A2(N6806), .A3(N8277) );
  AND3_X1 AND3_2356( .ZN(N8865), .A1(N6809), .A2(N5762), .A3(N8278) );
  AND3_X1 AND3_2357( .ZN(N8866), .A1(N5758), .A2(N6812), .A3(N8279) );
  INV_X2 NOT1_2358( .ZN(N8871), .A(N7655) );
  AND2_X1 AND2_2359( .ZN(N8874), .A1(N6833), .A2(N7655) );
  AND2_X1 AND2_2360( .ZN(N8878), .A1(N7671), .A2(N6867) );
  INV_X2 NOT1_2361( .ZN(N8879), .A(N8196) );
  NAND2_X1 NAND2_2362( .ZN(N8880), .A1(N8196), .A2(N8315) );
  INV_X1 NOT1_2363( .ZN(N8881), .A(N8200) );
  NAND2_X1 NAND2_2364( .ZN(N8882), .A1(N8200), .A2(N8317) );
  INV_X1 NOT1_2365( .ZN(N8883), .A(N8204) );
  NAND2_X1 NAND2_2366( .ZN(N8884), .A1(N8204), .A2(N8319) );
  INV_X1 NOT1_2367( .ZN(N8885), .A(N8208) );
  NAND2_X1 NAND2_2368( .ZN(N8886), .A1(N8208), .A2(N8321) );
  NAND2_X1 NAND2_2369( .ZN(N8887), .A1(N3658), .A2(N8323) );
  NAND2_X1 NAND2_2370( .ZN(N8888), .A1(N4817), .A2(N8325) );
  OR4_X1 OR4_2371( .ZN(N8898), .A1(N4544), .A2(N8337), .A3(N8338), .A4(N8339) );
  OR4_X1 OR5_2372_A( .ZN(extra32), .A1(N4562), .A2(N8348), .A3(N8349), .A4(N8350) );
  OR2_X1 OR5_2372( .ZN(N8902), .A1(extra32), .A2(N8351) );
  OR4_X1 OR4_2373( .ZN(N8920), .A1(N4576), .A2(N8369), .A3(N8370), .A4(N8371) );
  OR2_X1 OR2_2374( .ZN(N8924), .A1(N4581), .A2(N8377) );
  OR4_X1 OR5_2375_A( .ZN(extra33), .A1(N4592), .A2(N8378), .A3(N8379), .A4(N8380) );
  OR2_X2 OR5_2375( .ZN(N8927), .A1(extra33), .A2(N8381) );
  OR2_X2 OR2_2376( .ZN(N8931), .A1(N4603), .A2(N8392) );
  OR2_X1 OR2_2377( .ZN(N8943), .A1(N7825), .A2(N8404) );
  OR4_X1 OR4_2378( .ZN(N8950), .A1(N4630), .A2(N8409), .A3(N8410), .A4(N8411) );
  OR4_X1 OR5_2379_A( .ZN(extra34), .A1(N4637), .A2(N8415), .A3(N8416), .A4(N8417) );
  OR2_X1 OR5_2379( .ZN(N8956), .A1(extra34), .A2(N8418) );
  INV_X1 NOT1_2380( .ZN(N8959), .A(N7852) );
  AND2_X1 AND2_2381( .ZN(N8960), .A1(N3375), .A2(N7852) );
  OR4_X1 OR4_2382( .ZN(N8963), .A1(N4656), .A2(N8433), .A3(N8434), .A4(N8435) );
  OR4_X1 OR5_2383_A( .ZN(extra35), .A1(N4674), .A2(N8447), .A3(N8448), .A4(N8449) );
  OR2_X1 OR5_2383( .ZN(N8966), .A1(extra35), .A2(N8450) );
  AND3_X1 AND3_2384( .ZN(N8991), .A1(N7188), .A2(N6083), .A3(N8469) );
  AND3_X1 AND3_2385( .ZN(N8992), .A1(N6079), .A2(N7191), .A3(N8470) );
  OR4_X1 OR4_2386( .ZN(N8995), .A1(N4701), .A2(N8488), .A3(N8489), .A4(N8490) );
  OR2_X1 OR2_2387( .ZN(N8996), .A1(N4706), .A2(N8496) );
  OR4_X1 OR5_2388_A( .ZN(extra36), .A1(N4717), .A2(N8500), .A3(N8501), .A4(N8502) );
  OR2_X1 OR5_2388( .ZN(N9001), .A1(extra36), .A2(N8503) );
  OR2_X1 OR2_2389( .ZN(N9005), .A1(N4728), .A2(N8516) );
  AND3_X1 AND3_2390( .ZN(N9024), .A1(N7334), .A2(N6141), .A3(N8537) );
  AND3_X1 AND3_2391( .ZN(N9025), .A1(N6137), .A2(N7337), .A3(N8538) );
  OR4_X1 OR4_2392( .ZN(N9029), .A1(N4756), .A2(N8545), .A3(N8546), .A4(N8547) );
  OR4_X1 OR5_2393_A( .ZN(extra37), .A1(N4760), .A2(N8551), .A3(N8552), .A4(N8553) );
  OR2_X1 OR5_2393( .ZN(N9035), .A1(extra37), .A2(N8554) );
  AND3_X1 AND3_2394( .ZN(N9053), .A1(N7378), .A2(N6170), .A3(N8564) );
  AND3_X1 AND3_2395( .ZN(N9054), .A1(N6166), .A2(N7381), .A3(N8565) );
  NAND2_X1 NAND2_2396( .ZN(N9064), .A1(N4303), .A2(N8607) );
  NAND2_X1 NAND2_2397( .ZN(N9065), .A1(N3507), .A2(N8609) );
  INV_X1 NOT1_2398( .ZN(N9066), .A(N8114) );
  NAND2_X1 NAND2_2399( .ZN(N9067), .A1(N8114), .A2(N4795) );
  OR2_X1 OR2_2400( .ZN(N9068), .A1(N7613), .A2(N6783) );
  INV_X1 NOT1_2401( .ZN(N9071), .A(N8117) );
  INV_X1 NOT1_2402( .ZN(N9072), .A(N8131) );
  NAND2_X1 NAND2_2403( .ZN(N9073), .A1(N8131), .A2(N6195) );
  INV_X1 NOT1_2404( .ZN(N9074), .A(N7613) );
  INV_X1 NOT1_2405( .ZN(N9077), .A(N8134) );
  OR2_X1 OR2_2406( .ZN(N9079), .A1(N7650), .A2(N6865) );
  INV_X1 NOT1_2407( .ZN(N9082), .A(N8146) );
  INV_X1 NOT1_2408( .ZN(N9083), .A(N7650) );
  INV_X1 NOT1_2409( .ZN(N9086), .A(N8156) );
  INV_X1 NOT1_2410( .ZN(N9087), .A(N8166) );
  NAND2_X1 NAND2_2411( .ZN(N9088), .A1(N8166), .A2(N4813) );
  OR2_X1 OR2_2412( .ZN(N9089), .A1(N7659), .A2(N6866) );
  INV_X1 NOT1_2413( .ZN(N9092), .A(N8169) );
  INV_X1 NOT1_2414( .ZN(N9093), .A(N8183) );
  NAND2_X1 NAND2_2415( .ZN(N9094), .A1(N8183), .A2(N6203) );
  INV_X1 NOT1_2416( .ZN(N9095), .A(N7659) );
  INV_X1 NOT1_2417( .ZN(N9098), .A(N8186) );
  OR4_X1 OR4_2418( .ZN(N9099), .A1(N4545), .A2(N8340), .A3(N8341), .A4(N8342) );
  NOR3_X2 NOR3_2419( .ZN(N9103), .A1(N4545), .A2(N8343), .A3(N8344) );
  OR3_X2 OR3_2420( .ZN(N9107), .A1(N4549), .A2(N8345), .A3(N8346) );
  NOR2_X1 NOR2_2421( .ZN(N9111), .A1(N4549), .A2(N8347) );
  OR4_X1 OR4_2422( .ZN(N9117), .A1(N4577), .A2(N8372), .A3(N8373), .A4(N8374) );
  NOR3_X1 NOR3_2423( .ZN(N9127), .A1(N4577), .A2(N8375), .A3(N8376) );
  NOR3_X1 NOR3_2424( .ZN(N9146), .A1(N4597), .A2(N8390), .A3(N8391) );
  NOR3_X1 NOR4_2425_A( .ZN(extra38), .A1(N4593), .A2(N8385), .A3(N8386) );
  NOR2_X1 NOR4_2425( .ZN(N9149), .A1(extra38), .A2(N8387) );
  NAND2_X1 NAND2_2426( .ZN(N9159), .A1(N7577), .A2(N8733) );
  NAND2_X1 NAND2_2427( .ZN(N9160), .A1(N7574), .A2(N8734) );
  OR4_X1 OR4_2428( .ZN(N9161), .A1(N4657), .A2(N8436), .A3(N8437), .A4(N8438) );
  NOR3_X1 NOR3_2429( .ZN(N9165), .A1(N4657), .A2(N8439), .A3(N8440) );
  OR3_X1 OR3_2430( .ZN(N9169), .A1(N4661), .A2(N8441), .A3(N8442) );
  NOR2_X1 NOR2_2431( .ZN(N9173), .A1(N4661), .A2(N8443) );
  NAND2_X1 NAND2_2432( .ZN(N9179), .A1(N7563), .A2(N8753) );
  NAND2_X1 NAND2_2433( .ZN(N9180), .A1(N7560), .A2(N8754) );
  NAND2_X1 NAND2_2434( .ZN(N9181), .A1(N7569), .A2(N8755) );
  NAND2_X1 NAND2_2435( .ZN(N9182), .A1(N7566), .A2(N8756) );
  OR4_X1 OR4_2436( .ZN(N9183), .A1(N4702), .A2(N8491), .A3(N8492), .A4(N8493) );
  NOR3_X1 NOR3_2437( .ZN(N9193), .A1(N4702), .A2(N8494), .A3(N8495) );
  OR4_X1 OR4_2438( .ZN(N9203), .A1(N4722), .A2(N8511), .A3(N8512), .A4(N8513) );
  OR4_X1 OR5_2439_A( .ZN(extra39), .A1(N4718), .A2(N8504), .A3(N8505), .A4(N8506) );
  OR2_X1 OR5_2439( .ZN(N9206), .A1(extra39), .A2(N8507) );
  NOR3_X1 NOR3_2440( .ZN(N9220), .A1(N4722), .A2(N8514), .A3(N8515) );
  NOR3_X1 NOR4_2441_A( .ZN(extra40), .A1(N4718), .A2(N8508), .A3(N8509) );
  NOR2_X1 NOR4_2441( .ZN(N9223), .A1(extra40), .A2(N8510) );
  NAND2_X2 NAND2_2442( .ZN(N9234), .A1(N7591), .A2(N8814) );
  NAND2_X1 NAND2_2443( .ZN(N9235), .A1(N7588), .A2(N8815) );
  NAND2_X1 NAND2_2444( .ZN(N9236), .A1(N7585), .A2(N8816) );
  NAND2_X1 NAND2_2445( .ZN(N9237), .A1(N7582), .A2(N8817) );
  OR2_X1 OR2_2446( .ZN(N9238), .A1(N3159), .A2(N8818) );
  OR2_X1 OR2_2447( .ZN(N9242), .A1(N3126), .A2(N8840) );
  NAND2_X1 NAND2_2448( .ZN(N9243), .A1(N8324), .A2(N8888) );
  INV_X2 NOT1_2449( .ZN(N9244), .A(N8580) );
  INV_X2 NOT1_2450( .ZN(N9245), .A(N8583) );
  INV_X2 NOT1_2451( .ZN(N9246), .A(N8586) );
  INV_X1 NOT1_2452( .ZN(N9247), .A(N8589) );
  INV_X1 NOT1_2453( .ZN(N9248), .A(N8592) );
  INV_X1 NOT1_2454( .ZN(N9249), .A(N8595) );
  INV_X1 NOT1_2455( .ZN(N9250), .A(N8598) );
  INV_X1 NOT1_2456( .ZN(N9251), .A(N8601) );
  INV_X1 NOT1_2457( .ZN(N9252), .A(N8604) );
  NOR2_X1 NOR2_2458( .ZN(N9256), .A1(N8861), .A2(N8280) );
  NOR2_X1 NOR2_2459( .ZN(N9257), .A1(N8862), .A2(N8281) );
  NOR2_X1 NOR2_2460( .ZN(N9258), .A1(N8863), .A2(N8282) );
  NOR2_X1 NOR2_2461( .ZN(N9259), .A1(N8864), .A2(N8283) );
  NOR2_X1 NOR2_2462( .ZN(N9260), .A1(N8865), .A2(N8284) );
  NOR2_X1 NOR2_2463( .ZN(N9261), .A1(N8866), .A2(N8285) );
  INV_X1 NOT1_2464( .ZN(N9262), .A(N8627) );
  OR2_X1 OR2_2465( .ZN(N9265), .A1(N7649), .A2(N8874) );
  OR2_X1 OR2_2466( .ZN(N9268), .A1(N7668), .A2(N8878) );
  NAND2_X1 NAND2_2467( .ZN(N9271), .A1(N7533), .A2(N8879) );
  NAND2_X1 NAND2_2468( .ZN(N9272), .A1(N7536), .A2(N8881) );
  NAND2_X1 NAND2_2469( .ZN(N9273), .A1(N7539), .A2(N8883) );
  NAND2_X1 NAND2_2470( .ZN(N9274), .A1(N7542), .A2(N8885) );
  NAND2_X1 NAND2_2471( .ZN(N9275), .A1(N8322), .A2(N8887) );
  INV_X1 NOT1_2472( .ZN(N9276), .A(N8333) );
  AND4_X1 AND5_2473_A( .ZN(extra41), .A1(N6936), .A2(N8326), .A3(N6946), .A4(N6929) );
  AND2_X2 AND5_2473( .ZN(N9280), .A1(extra41), .A2(N6957) );
  AND4_X1 AND5_2474_A( .ZN(extra42), .A1(N367), .A2(N8326), .A3(N6946), .A4(N6957) );
  AND2_X1 AND5_2474( .ZN(N9285), .A1(extra42), .A2(N6936) );
  AND4_X1 AND4_2475( .ZN(N9286), .A1(N367), .A2(N8326), .A3(N6946), .A4(N6957) );
  AND3_X1 AND3_2476( .ZN(N9287), .A1(N367), .A2(N8326), .A3(N6957) );
  AND2_X1 AND2_2477( .ZN(N9288), .A1(N367), .A2(N8326) );
  INV_X1 NOT1_2478( .ZN(N9290), .A(N8660) );
  INV_X1 NOT1_2479( .ZN(N9292), .A(N8663) );
  INV_X1 NOT1_2480( .ZN(N9294), .A(N8666) );
  INV_X1 NOT1_2481( .ZN(N9296), .A(N8669) );
  NAND2_X1 NAND2_2482( .ZN(N9297), .A1(N8672), .A2(N5966) );
  INV_X1 NOT1_2483( .ZN(N9298), .A(N8672) );
  NAND2_X1 NAND2_2484( .ZN(N9299), .A1(N8675), .A2(N6969) );
  INV_X1 NOT1_2485( .ZN(N9300), .A(N8675) );
  INV_X1 NOT1_2486( .ZN(N9301), .A(N8365) );
  AND4_X1 AND5_2487_A( .ZN(extra43), .A1(N8358), .A2(N7036), .A3(N7020), .A4(N7006) );
  AND2_X1 AND5_2487( .ZN(N9307), .A1(extra43), .A2(N6998) );
  AND4_X1 AND4_2488( .ZN(N9314), .A1(N8358), .A2(N7020), .A3(N7006), .A4(N7036) );
  AND3_X1 AND3_2489( .ZN(N9315), .A1(N8358), .A2(N7020), .A3(N7036) );
  AND2_X1 AND2_2490( .ZN(N9318), .A1(N8358), .A2(N7036) );
  INV_X1 NOT1_2491( .ZN(N9319), .A(N8687) );
  INV_X1 NOT1_2492( .ZN(N9320), .A(N8699) );
  INV_X1 NOT1_2493( .ZN(N9321), .A(N8711) );
  INV_X1 NOT1_2494( .ZN(N9322), .A(N8714) );
  INV_X1 NOT1_2495( .ZN(N9323), .A(N8727) );
  INV_X1 NOT1_2496( .ZN(N9324), .A(N8730) );
  INV_X1 NOT1_2497( .ZN(N9326), .A(N8405) );
  AND2_X1 AND2_2498( .ZN(N9332), .A1(N8405), .A2(N8412) );
  OR2_X1 OR2_2499( .ZN(N9339), .A1(N4193), .A2(N8960) );
  AND2_X1 AND2_2500( .ZN(N9344), .A1(N8430), .A2(N8444) );
  INV_X1 NOT1_2501( .ZN(N9352), .A(N8735) );
  INV_X1 NOT1_2502( .ZN(N9354), .A(N8738) );
  INV_X1 NOT1_2503( .ZN(N9356), .A(N8741) );
  INV_X1 NOT1_2504( .ZN(N9358), .A(N8744) );
  NAND2_X1 NAND2_2505( .ZN(N9359), .A1(N8747), .A2(N6078) );
  INV_X1 NOT1_2506( .ZN(N9360), .A(N8747) );
  NAND2_X1 NAND2_2507( .ZN(N9361), .A1(N8750), .A2(N7187) );
  INV_X1 NOT1_2508( .ZN(N9362), .A(N8750) );
  INV_X1 NOT1_2509( .ZN(N9363), .A(N8471) );
  INV_X1 NOT1_2510( .ZN(N9364), .A(N8474) );
  INV_X1 NOT1_2511( .ZN(N9365), .A(N8477) );
  INV_X1 NOT1_2512( .ZN(N9366), .A(N8480) );
  NOR2_X1 NOR2_2513( .ZN(N9367), .A1(N8991), .A2(N8483) );
  NOR2_X1 NOR2_2514( .ZN(N9368), .A1(N8992), .A2(N8484) );
  AND3_X1 AND3_2515( .ZN(N9369), .A1(N7198), .A2(N7194), .A3(N8471) );
  AND3_X1 AND3_2516( .ZN(N9370), .A1(N8460), .A2(N8457), .A3(N8474) );
  AND3_X1 AND3_2517( .ZN(N9371), .A1(N7209), .A2(N7205), .A3(N8477) );
  AND3_X1 AND3_2518( .ZN(N9372), .A1(N8466), .A2(N8463), .A3(N8480) );
  INV_X1 NOT1_2519( .ZN(N9375), .A(N8497) );
  INV_X1 NOT1_2520( .ZN(N9381), .A(N8766) );
  INV_X1 NOT1_2521( .ZN(N9382), .A(N8778) );
  INV_X1 NOT1_2522( .ZN(N9383), .A(N8793) );
  INV_X1 NOT1_2523( .ZN(N9384), .A(N8796) );
  AND2_X1 AND2_2524( .ZN(N9385), .A1(N8485), .A2(N8497) );
  INV_X1 NOT1_2525( .ZN(N9392), .A(N8525) );
  INV_X1 NOT1_2526( .ZN(N9393), .A(N8528) );
  INV_X1 NOT1_2527( .ZN(N9394), .A(N8531) );
  INV_X1 NOT1_2528( .ZN(N9395), .A(N8534) );
  AND3_X1 AND3_2529( .ZN(N9396), .A1(N7318), .A2(N7314), .A3(N8525) );
  AND3_X1 AND3_2530( .ZN(N9397), .A1(N8522), .A2(N8519), .A3(N8528) );
  AND3_X1 AND3_2531( .ZN(N9398), .A1(N6131), .A2(N6127), .A3(N8531) );
  AND3_X1 AND3_2532( .ZN(N9399), .A1(N7328), .A2(N7325), .A3(N8534) );
  NOR2_X1 NOR2_2533( .ZN(N9400), .A1(N9024), .A2(N8539) );
  NOR2_X1 NOR2_2534( .ZN(N9401), .A1(N9025), .A2(N8540) );
  INV_X1 NOT1_2535( .ZN(N9402), .A(N8541) );
  NAND2_X1 NAND2_2536( .ZN(N9407), .A1(N8548), .A2(N89) );
  AND2_X1 AND2_2537( .ZN(N9408), .A1(N8541), .A2(N8548) );
  INV_X1 NOT1_2538( .ZN(N9412), .A(N8811) );
  INV_X1 NOT1_2539( .ZN(N9413), .A(N8566) );
  INV_X1 NOT1_2540( .ZN(N9414), .A(N8569) );
  INV_X1 NOT1_2541( .ZN(N9415), .A(N8572) );
  INV_X1 NOT1_2542( .ZN(N9416), .A(N8575) );
  NOR2_X1 NOR2_2543( .ZN(N9417), .A1(N9053), .A2(N8578) );
  NOR2_X1 NOR2_2544( .ZN(N9418), .A1(N9054), .A2(N8579) );
  AND3_X1 AND3_2545( .ZN(N9419), .A1(N7387), .A2(N6177), .A3(N8566) );
  AND3_X1 AND3_2546( .ZN(N9420), .A1(N8555), .A2(N7384), .A3(N8569) );
  AND3_X1 AND3_2547( .ZN(N9421), .A1(N7398), .A2(N7394), .A3(N8572) );
  AND3_X1 AND3_2548( .ZN(N9422), .A1(N8561), .A2(N8558), .A3(N8575) );
  BUF_X4 BUFF1_2549( .Z(N9423), .A(N8326) );
  NAND2_X1 NAND2_2550( .ZN(N9426), .A1(N9064), .A2(N8608) );
  NAND2_X1 NAND2_2551( .ZN(N9429), .A1(N9065), .A2(N8610) );
  NAND2_X1 NAND2_2552( .ZN(N9432), .A1(N3515), .A2(N9066) );
  NAND2_X1 NAND2_2553( .ZN(N9435), .A1(N4796), .A2(N9072) );
  NAND2_X1 NAND2_2554( .ZN(N9442), .A1(N3628), .A2(N9087) );
  NAND2_X1 NAND2_2555( .ZN(N9445), .A1(N4814), .A2(N9093) );
  INV_X1 NOT1_2556( .ZN(N9454), .A(N8678) );
  INV_X1 NOT1_2557( .ZN(N9455), .A(N8681) );
  INV_X1 NOT1_2558( .ZN(N9456), .A(N8684) );
  INV_X1 NOT1_2559( .ZN(N9459), .A(N8690) );
  INV_X1 NOT1_2560( .ZN(N9460), .A(N8693) );
  INV_X1 NOT1_2561( .ZN(N9461), .A(N8696) );
  BUF_X1 BUFF1_2562( .Z(N9462), .A(N8358) );
  INV_X1 NOT1_2563( .ZN(N9465), .A(N8702) );
  INV_X1 NOT1_2564( .ZN(N9466), .A(N8705) );
  INV_X1 NOT1_2565( .ZN(N9467), .A(N8708) );
  INV_X1 NOT1_2566( .ZN(N9468), .A(N8724) );
  BUF_X1 BUFF1_2567( .Z(N9473), .A(N8358) );
  INV_X1 NOT1_2568( .ZN(N9476), .A(N8718) );
  INV_X1 NOT1_2569( .ZN(N9477), .A(N8721) );
  NAND2_X1 NAND2_2570( .ZN(N9478), .A1(N9159), .A2(N9160) );
  NAND2_X1 NAND2_2571( .ZN(N9485), .A1(N9179), .A2(N9180) );
  NAND2_X1 NAND2_2572( .ZN(N9488), .A1(N9181), .A2(N9182) );
  INV_X1 NOT1_2573( .ZN(N9493), .A(N8757) );
  INV_X1 NOT1_2574( .ZN(N9494), .A(N8760) );
  INV_X1 NOT1_2575( .ZN(N9495), .A(N8763) );
  INV_X1 NOT1_2576( .ZN(N9498), .A(N8769) );
  INV_X1 NOT1_2577( .ZN(N9499), .A(N8772) );
  INV_X1 NOT1_2578( .ZN(N9500), .A(N8775) );
  INV_X1 NOT1_2579( .ZN(N9505), .A(N8781) );
  INV_X1 NOT1_2580( .ZN(N9506), .A(N8784) );
  INV_X1 NOT1_2581( .ZN(N9507), .A(N8787) );
  INV_X1 NOT1_2582( .ZN(N9508), .A(N8790) );
  INV_X1 NOT1_2583( .ZN(N9509), .A(N8808) );
  INV_X1 NOT1_2584( .ZN(N9514), .A(N8799) );
  INV_X1 NOT1_2585( .ZN(N9515), .A(N8802) );
  INV_X1 NOT1_2586( .ZN(N9516), .A(N8805) );
  NAND2_X2 NAND2_2587( .ZN(N9517), .A1(N9234), .A2(N9235) );
  NAND2_X1 NAND2_2588( .ZN(N9520), .A1(N9236), .A2(N9237) );
  AND2_X1 AND2_2589( .ZN(N9526), .A1(N8943), .A2(N8421) );
  AND2_X1 AND2_2590( .ZN(N9531), .A1(N8943), .A2(N8421) );
  NAND2_X1 NAND2_2591( .ZN(N9539), .A1(N9271), .A2(N8880) );
  NAND2_X1 NAND2_2592( .ZN(N9540), .A1(N9273), .A2(N8884) );
  INV_X1 NOT1_2593( .ZN(N9541), .A(N9275) );
  AND2_X1 AND2_2594( .ZN(N9543), .A1(N8857), .A2(N8254) );
  AND2_X1 AND2_2595( .ZN(N9551), .A1(N8871), .A2(N8288) );
  NAND2_X1 NAND2_2596( .ZN(N9555), .A1(N9272), .A2(N8882) );
  NAND2_X1 NAND2_2597( .ZN(N9556), .A1(N9274), .A2(N8886) );
  INV_X1 NOT1_2598( .ZN(N9557), .A(N8898) );
  AND2_X1 AND2_2599( .ZN(N9560), .A1(N8902), .A2(N8333) );
  INV_X1 NOT1_2600( .ZN(N9561), .A(N9099) );
  NAND2_X1 NAND2_2601( .ZN(N9562), .A1(N9099), .A2(N9290) );
  INV_X1 NOT1_2602( .ZN(N9563), .A(N9103) );
  NAND2_X1 NAND2_2603( .ZN(N9564), .A1(N9103), .A2(N9292) );
  INV_X1 NOT1_2604( .ZN(N9565), .A(N9107) );
  NAND2_X1 NAND2_2605( .ZN(N9566), .A1(N9107), .A2(N9294) );
  INV_X1 NOT1_2606( .ZN(N9567), .A(N9111) );
  NAND2_X1 NAND2_2607( .ZN(N9568), .A1(N9111), .A2(N9296) );
  NAND2_X1 NAND2_2608( .ZN(N9569), .A1(N4844), .A2(N9298) );
  NAND2_X1 NAND2_2609( .ZN(N9570), .A1(N6207), .A2(N9300) );
  INV_X1 NOT1_2610( .ZN(N9571), .A(N8920) );
  INV_X1 NOT1_2611( .ZN(N9575), .A(N8927) );
  AND2_X1 AND2_2612( .ZN(N9579), .A1(N8365), .A2(N8927) );
  INV_X1 NOT1_2613( .ZN(N9581), .A(N8950) );
  INV_X1 NOT1_2614( .ZN(N9582), .A(N8956) );
  AND2_X2 AND2_2615( .ZN(N9585), .A1(N8405), .A2(N8956) );
  AND2_X1 AND2_2616( .ZN(N9591), .A1(N8966), .A2(N8430) );
  INV_X1 NOT1_2617( .ZN(N9592), .A(N9161) );
  NAND2_X1 NAND2_2618( .ZN(N9593), .A1(N9161), .A2(N9352) );
  INV_X1 NOT1_2619( .ZN(N9594), .A(N9165) );
  NAND2_X1 NAND2_2620( .ZN(N9595), .A1(N9165), .A2(N9354) );
  INV_X1 NOT1_2621( .ZN(N9596), .A(N9169) );
  NAND2_X1 NAND2_2622( .ZN(N9597), .A1(N9169), .A2(N9356) );
  INV_X1 NOT1_2623( .ZN(N9598), .A(N9173) );
  NAND2_X1 NAND2_2624( .ZN(N9599), .A1(N9173), .A2(N9358) );
  NAND2_X1 NAND2_2625( .ZN(N9600), .A1(N4940), .A2(N9360) );
  NAND2_X1 NAND2_2626( .ZN(N9601), .A1(N6220), .A2(N9362) );
  AND3_X1 AND3_2627( .ZN(N9602), .A1(N8457), .A2(N7198), .A3(N9363) );
  AND3_X1 AND3_2628( .ZN(N9603), .A1(N7194), .A2(N8460), .A3(N9364) );
  AND3_X1 AND3_2629( .ZN(N9604), .A1(N8463), .A2(N7209), .A3(N9365) );
  AND3_X1 AND3_2630( .ZN(N9605), .A1(N7205), .A2(N8466), .A3(N9366) );
  INV_X2 NOT1_2631( .ZN(N9608), .A(N9001) );
  AND2_X1 AND2_2632( .ZN(N9611), .A1(N8485), .A2(N9001) );
  AND3_X1 AND3_2633( .ZN(N9612), .A1(N8519), .A2(N7318), .A3(N9392) );
  AND3_X1 AND3_2634( .ZN(N9613), .A1(N7314), .A2(N8522), .A3(N9393) );
  AND3_X1 AND3_2635( .ZN(N9614), .A1(N7325), .A2(N6131), .A3(N9394) );
  AND3_X1 AND3_2636( .ZN(N9615), .A1(N6127), .A2(N7328), .A3(N9395) );
  INV_X2 NOT1_2637( .ZN(N9616), .A(N9029) );
  INV_X1 NOT1_2638( .ZN(N9617), .A(N9035) );
  AND2_X1 AND2_2639( .ZN(N9618), .A1(N8541), .A2(N9035) );
  AND3_X1 AND3_2640( .ZN(N9621), .A1(N7384), .A2(N7387), .A3(N9413) );
  AND3_X1 AND3_2641( .ZN(N9622), .A1(N6177), .A2(N8555), .A3(N9414) );
  AND3_X1 AND3_2642( .ZN(N9623), .A1(N8558), .A2(N7398), .A3(N9415) );
  AND3_X1 AND3_2643( .ZN(N9624), .A1(N7394), .A2(N8561), .A3(N9416) );
  OR4_X2 OR5_2644_A( .ZN(extra44), .A1(N4563), .A2(N8352), .A3(N8353), .A4(N8354) );
  OR2_X2 OR5_2644( .ZN(N9626), .A1(extra44), .A2(N9285) );
  OR4_X1 OR4_2645( .ZN(N9629), .A1(N4566), .A2(N8355), .A3(N8356), .A4(N9286) );
  OR3_X1 OR3_2646( .ZN(N9632), .A1(N4570), .A2(N8357), .A3(N9287) );
  OR2_X1 OR2_2647( .ZN(N9635), .A1(N5960), .A2(N9288) );
  NAND2_X1 NAND2_2648( .ZN(N9642), .A1(N9067), .A2(N9432) );
  INV_X1 NOT1_2649( .ZN(N9645), .A(N9068) );
  NAND2_X1 NAND2_2650( .ZN(N9646), .A1(N9073), .A2(N9435) );
  INV_X1 NOT1_2651( .ZN(N9649), .A(N9074) );
  NAND2_X1 NAND2_2652( .ZN(N9650), .A1(N9257), .A2(N9256) );
  NAND2_X1 NAND2_2653( .ZN(N9653), .A1(N9259), .A2(N9258) );
  NAND2_X1 NAND2_2654( .ZN(N9656), .A1(N9261), .A2(N9260) );
  INV_X1 NOT1_2655( .ZN(N9659), .A(N9079) );
  NAND2_X1 NAND2_2656( .ZN(N9660), .A1(N9079), .A2(N4809) );
  INV_X1 NOT1_2657( .ZN(N9661), .A(N9083) );
  NAND2_X1 NAND2_2658( .ZN(N9662), .A1(N9083), .A2(N6202) );
  NAND2_X1 NAND2_2659( .ZN(N9663), .A1(N9088), .A2(N9442) );
  INV_X1 NOT1_2660( .ZN(N9666), .A(N9089) );
  NAND2_X1 NAND2_2661( .ZN(N9667), .A1(N9094), .A2(N9445) );
  INV_X1 NOT1_2662( .ZN(N9670), .A(N9095) );
  OR2_X1 OR2_2663( .ZN(N9671), .A1(N8924), .A2(N8393) );
  INV_X1 NOT1_2664( .ZN(N9674), .A(N9117) );
  INV_X1 NOT1_2665( .ZN(N9675), .A(N8924) );
  INV_X1 NOT1_2666( .ZN(N9678), .A(N9127) );
  OR4_X1 OR4_2667( .ZN(N9679), .A1(N4597), .A2(N8388), .A3(N8389), .A4(N9315) );
  OR2_X1 OR2_2668( .ZN(N9682), .A1(N8931), .A2(N9318) );
  OR4_X1 OR5_2669_A( .ZN(extra45), .A1(N4593), .A2(N8382), .A3(N8383), .A4(N8384) );
  OR2_X1 OR5_2669( .ZN(N9685), .A1(extra45), .A2(N9314) );
  INV_X1 NOT1_2670( .ZN(N9690), .A(N9146) );
  NAND2_X1 NAND2_2671( .ZN(N9691), .A1(N9146), .A2(N8717) );
  INV_X1 NOT1_2672( .ZN(N9692), .A(N8931) );
  INV_X1 NOT1_2673( .ZN(N9695), .A(N9149) );
  NAND2_X1 NAND2_2674( .ZN(N9698), .A1(N9401), .A2(N9400) );
  NAND2_X1 NAND2_2675( .ZN(N9702), .A1(N9368), .A2(N9367) );
  OR2_X1 OR2_2676( .ZN(N9707), .A1(N8996), .A2(N8517) );
  INV_X1 NOT1_2677( .ZN(N9710), .A(N9183) );
  INV_X1 NOT1_2678( .ZN(N9711), .A(N8996) );
  INV_X1 NOT1_2679( .ZN(N9714), .A(N9193) );
  INV_X1 NOT1_2680( .ZN(N9715), .A(N9203) );
  NAND2_X1 NAND2_2681( .ZN(N9716), .A1(N9203), .A2(N6235) );
  OR2_X1 OR2_2682( .ZN(N9717), .A1(N9005), .A2(N8518) );
  INV_X1 NOT1_2683( .ZN(N9720), .A(N9206) );
  INV_X1 NOT1_2684( .ZN(N9721), .A(N9220) );
  NAND2_X1 NAND2_2685( .ZN(N9722), .A1(N9220), .A2(N7573) );
  INV_X1 NOT1_2686( .ZN(N9723), .A(N9005) );
  INV_X1 NOT1_2687( .ZN(N9726), .A(N9223) );
  NAND2_X1 NAND2_2688( .ZN(N9727), .A1(N9418), .A2(N9417) );
  AND2_X1 AND2_2689( .ZN(N9732), .A1(N9268), .A2(N8269) );
  NAND2_X1 NAND2_2690( .ZN(N9733), .A1(N9581), .A2(N9326) );
  AND4_X1 AND5_2691_A( .ZN(extra46), .A1(N89), .A2(N9408), .A3(N9332), .A4(N8394) );
  AND2_X1 AND5_2691( .ZN(N9734), .A1(extra46), .A2(N8421) );
  AND4_X1 AND5_2692_A( .ZN(extra47), .A1(N89), .A2(N9408), .A3(N9332), .A4(N8394) );
  AND2_X1 AND5_2692( .ZN(N9735), .A1(extra47), .A2(N8421) );
  AND2_X1 AND2_2693( .ZN(N9736), .A1(N9265), .A2(N8262) );
  INV_X1 NOT1_2694( .ZN(N9737), .A(N9555) );
  INV_X1 NOT1_2695( .ZN(N9738), .A(N9556) );
  NAND2_X1 NAND2_2696( .ZN(N9739), .A1(N9361), .A2(N9601) );
  NAND2_X1 NAND2_2697( .ZN(N9740), .A1(N9423), .A2(N1115) );
  INV_X1 NOT1_2698( .ZN(N9741), .A(N9423) );
  NAND2_X1 NAND2_2699( .ZN(N9742), .A1(N9299), .A2(N9570) );
  AND2_X1 AND2_2700( .ZN(N9754), .A1(N8333), .A2(N9280) );
  OR2_X1 OR2_2701( .ZN(N9758), .A1(N8898), .A2(N9560) );
  NAND2_X1 NAND2_2702( .ZN(N9762), .A1(N8660), .A2(N9561) );
  NAND2_X1 NAND2_2703( .ZN(N9763), .A1(N8663), .A2(N9563) );
  NAND2_X1 NAND2_2704( .ZN(N9764), .A1(N8666), .A2(N9565) );
  NAND2_X1 NAND2_2705( .ZN(N9765), .A1(N8669), .A2(N9567) );
  NAND2_X1 NAND2_2706( .ZN(N9766), .A1(N9297), .A2(N9569) );
  AND2_X1 AND2_2707( .ZN(N9767), .A1(N9280), .A2(N367) );
  NAND2_X1 NAND2_2708( .ZN(N9768), .A1(N9557), .A2(N9276) );
  INV_X1 NOT1_2709( .ZN(N9769), .A(N9307) );
  NAND2_X1 NAND2_2710( .ZN(N9773), .A1(N9307), .A2(N367) );
  NAND2_X1 NAND2_2711( .ZN(N9774), .A1(N9571), .A2(N9301) );
  AND2_X1 AND2_2712( .ZN(N9775), .A1(N8365), .A2(N9307) );
  OR2_X1 OR2_2713( .ZN(N9779), .A1(N8920), .A2(N9579) );
  INV_X1 NOT1_2714( .ZN(N9784), .A(N9478) );
  NAND2_X1 NAND2_2715( .ZN(N9785), .A1(N9616), .A2(N9402) );
  OR2_X1 OR2_2716( .ZN(N9786), .A1(N8950), .A2(N9585) );
  AND4_X1 AND4_2717( .ZN(N9790), .A1(N89), .A2(N9408), .A3(N9332), .A4(N8394) );
  OR2_X1 OR2_2718( .ZN(N9791), .A1(N8963), .A2(N9591) );
  NAND2_X1 NAND2_2719( .ZN(N9795), .A1(N8735), .A2(N9592) );
  NAND2_X1 NAND2_2720( .ZN(N9796), .A1(N8738), .A2(N9594) );
  NAND2_X2 NAND2_2721( .ZN(N9797), .A1(N8741), .A2(N9596) );
  NAND2_X2 NAND2_2722( .ZN(N9798), .A1(N8744), .A2(N9598) );
  NAND2_X1 NAND2_2723( .ZN(N9799), .A1(N9359), .A2(N9600) );
  NOR2_X1 NOR2_2724( .ZN(N9800), .A1(N9602), .A2(N9369) );
  NOR2_X1 NOR2_2725( .ZN(N9801), .A1(N9603), .A2(N9370) );
  NOR2_X2 NOR2_2726( .ZN(N9802), .A1(N9604), .A2(N9371) );
  NOR2_X2 NOR2_2727( .ZN(N9803), .A1(N9605), .A2(N9372) );
  INV_X2 NOT1_2728( .ZN(N9805), .A(N9485) );
  INV_X1 NOT1_2729( .ZN(N9806), .A(N9488) );
  OR2_X1 OR2_2730( .ZN(N9809), .A1(N8995), .A2(N9611) );
  NOR2_X1 NOR2_2731( .ZN(N9813), .A1(N9612), .A2(N9396) );
  NOR2_X1 NOR2_2732( .ZN(N9814), .A1(N9613), .A2(N9397) );
  NOR2_X1 NOR2_2733( .ZN(N9815), .A1(N9614), .A2(N9398) );
  NOR2_X1 NOR2_2734( .ZN(N9816), .A1(N9615), .A2(N9399) );
  AND2_X1 AND2_2735( .ZN(N9817), .A1(N9617), .A2(N9407) );
  OR2_X1 OR2_2736( .ZN(N9820), .A1(N9029), .A2(N9618) );
  INV_X1 NOT1_2737( .ZN(N9825), .A(N9517) );
  INV_X1 NOT1_2738( .ZN(N9826), .A(N9520) );
  NOR2_X1 NOR2_2739( .ZN(N9827), .A1(N9621), .A2(N9419) );
  NOR2_X1 NOR2_2740( .ZN(N9828), .A1(N9622), .A2(N9420) );
  NOR2_X1 NOR2_2741( .ZN(N9829), .A1(N9623), .A2(N9421) );
  NOR2_X1 NOR2_2742( .ZN(N9830), .A1(N9624), .A2(N9422) );
  INV_X1 NOT1_2743( .ZN(N9835), .A(N9426) );
  NAND2_X1 NAND2_2744( .ZN(N9836), .A1(N9426), .A2(N4789) );
  INV_X1 NOT1_2745( .ZN(N9837), .A(N9429) );
  NAND2_X1 NAND2_2746( .ZN(N9838), .A1(N9429), .A2(N4794) );
  NAND2_X1 NAND2_2747( .ZN(N9846), .A1(N3625), .A2(N9659) );
  NAND2_X1 NAND2_2748( .ZN(N9847), .A1(N4810), .A2(N9661) );
  INV_X1 NOT1_2749( .ZN(N9862), .A(N9462) );
  NAND2_X1 NAND2_2750( .ZN(N9863), .A1(N7553), .A2(N9690) );
  INV_X1 NOT1_2751( .ZN(N9866), .A(N9473) );
  NAND2_X1 NAND2_2752( .ZN(N9873), .A1(N5030), .A2(N9715) );
  NAND2_X1 NAND2_2753( .ZN(N9876), .A1(N6236), .A2(N9721) );
  NAND2_X1 NAND2_2754( .ZN(N9890), .A1(N9795), .A2(N9593) );
  NAND2_X1 NAND2_2755( .ZN(N9891), .A1(N9797), .A2(N9597) );
  INV_X1 NOT1_2756( .ZN(N9892), .A(N9799) );
  NAND2_X1 NAND2_2757( .ZN(N9893), .A1(N871), .A2(N9741) );
  NAND2_X1 NAND2_2758( .ZN(N9894), .A1(N9762), .A2(N9562) );
  NAND2_X1 NAND2_2759( .ZN(N9895), .A1(N9764), .A2(N9566) );
  INV_X1 NOT1_2760( .ZN(N9896), .A(N9766) );
  INV_X1 NOT1_2761( .ZN(N9897), .A(N9626) );
  NAND2_X1 NAND2_2762( .ZN(N9898), .A1(N9626), .A2(N9249) );
  INV_X1 NOT1_2763( .ZN(N9899), .A(N9629) );
  NAND2_X1 NAND2_2764( .ZN(N9900), .A1(N9629), .A2(N9250) );
  INV_X1 NOT1_2765( .ZN(N9901), .A(N9632) );
  NAND2_X1 NAND2_2766( .ZN(N9902), .A1(N9632), .A2(N9251) );
  INV_X1 NOT1_2767( .ZN(N9903), .A(N9635) );
  NAND2_X1 NAND2_2768( .ZN(N9904), .A1(N9635), .A2(N9252) );
  INV_X1 NOT1_2769( .ZN(N9905), .A(N9543) );
  INV_X1 NOT1_2770( .ZN(N9906), .A(N9650) );
  NAND2_X1 NAND2_2771( .ZN(N9907), .A1(N9650), .A2(N5769) );
  INV_X1 NOT1_2772( .ZN(N9908), .A(N9653) );
  NAND2_X1 NAND2_2773( .ZN(N9909), .A1(N9653), .A2(N5770) );
  INV_X1 NOT1_2774( .ZN(N9910), .A(N9656) );
  NAND2_X1 NAND2_2775( .ZN(N9911), .A1(N9656), .A2(N9262) );
  INV_X1 NOT1_2776( .ZN(N9917), .A(N9551) );
  NAND2_X1 NAND2_2777( .ZN(N9923), .A1(N9763), .A2(N9564) );
  NAND2_X1 NAND2_2778( .ZN(N9924), .A1(N9765), .A2(N9568) );
  OR2_X1 OR2_2779( .ZN(N9925), .A1(N8902), .A2(N9767) );
  AND2_X2 AND2_2780( .ZN(N9932), .A1(N9575), .A2(N9773) );
  AND2_X2 AND2_2781( .ZN(N9935), .A1(N9575), .A2(N9769) );
  INV_X1 NOT1_2782( .ZN(N9938), .A(N9698) );
  NAND2_X1 NAND2_2783( .ZN(N9939), .A1(N9698), .A2(N9323) );
  NAND2_X1 NAND2_2784( .ZN(N9945), .A1(N9796), .A2(N9595) );
  NAND2_X1 NAND2_2785( .ZN(N9946), .A1(N9798), .A2(N9599) );
  INV_X1 NOT1_2786( .ZN(N9947), .A(N9702) );
  NAND2_X1 NAND2_2787( .ZN(N9948), .A1(N9702), .A2(N6102) );
  AND2_X1 AND2_2788( .ZN(N9949), .A1(N9608), .A2(N9375) );
  INV_X1 NOT1_2789( .ZN(N9953), .A(N9727) );
  NAND2_X1 NAND2_2790( .ZN(N9954), .A1(N9727), .A2(N9412) );
  NAND2_X1 NAND2_2791( .ZN(N9955), .A1(N3502), .A2(N9835) );
  NAND2_X1 NAND2_2792( .ZN(N9956), .A1(N3510), .A2(N9837) );
  INV_X1 NOT1_2793( .ZN(N9957), .A(N9642) );
  NAND2_X1 NAND2_2794( .ZN(N9958), .A1(N9642), .A2(N9645) );
  INV_X1 NOT1_2795( .ZN(N9959), .A(N9646) );
  NAND2_X1 NAND2_2796( .ZN(N9960), .A1(N9646), .A2(N9649) );
  NAND2_X1 NAND2_2797( .ZN(N9961), .A1(N9660), .A2(N9846) );
  NAND2_X1 NAND2_2798( .ZN(N9964), .A1(N9662), .A2(N9847) );
  INV_X1 NOT1_2799( .ZN(N9967), .A(N9663) );
  NAND2_X1 NAND2_2800( .ZN(N9968), .A1(N9663), .A2(N9666) );
  INV_X1 NOT1_2801( .ZN(N9969), .A(N9667) );
  NAND2_X1 NAND2_2802( .ZN(N9970), .A1(N9667), .A2(N9670) );
  INV_X1 NOT1_2803( .ZN(N9971), .A(N9671) );
  NAND2_X1 NAND2_2804( .ZN(N9972), .A1(N9671), .A2(N6213) );
  INV_X1 NOT1_2805( .ZN(N9973), .A(N9675) );
  NAND2_X1 NAND2_2806( .ZN(N9974), .A1(N9675), .A2(N7551) );
  INV_X1 NOT1_2807( .ZN(N9975), .A(N9679) );
  NAND2_X1 NAND2_2808( .ZN(N9976), .A1(N9679), .A2(N7552) );
  INV_X1 NOT1_2809( .ZN(N9977), .A(N9682) );
  INV_X1 NOT1_2810( .ZN(N9978), .A(N9685) );
  NAND2_X1 NAND2_2811( .ZN(N9979), .A1(N9691), .A2(N9863) );
  INV_X1 NOT1_2812( .ZN(N9982), .A(N9692) );
  NAND2_X1 NAND2_2813( .ZN(N9983), .A1(N9814), .A2(N9813) );
  NAND2_X1 NAND2_2814( .ZN(N9986), .A1(N9816), .A2(N9815) );
  NAND2_X1 NAND2_2815( .ZN(N9989), .A1(N9801), .A2(N9800) );
  NAND2_X1 NAND2_2816( .ZN(N9992), .A1(N9803), .A2(N9802) );
  INV_X2 NOT1_2817( .ZN(N9995), .A(N9707) );
  NAND2_X1 NAND2_2818( .ZN(N9996), .A1(N9707), .A2(N6231) );
  INV_X1 NOT1_2819( .ZN(N9997), .A(N9711) );
  NAND2_X1 NAND2_2820( .ZN(N9998), .A1(N9711), .A2(N7572) );
  NAND2_X1 NAND2_2821( .ZN(N9999), .A1(N9716), .A2(N9873) );
  INV_X1 NOT1_2822( .ZN(N10002), .A(N9717) );
  NAND2_X1 NAND2_2823( .ZN(N10003), .A1(N9722), .A2(N9876) );
  INV_X1 NOT1_2824( .ZN(N10006), .A(N9723) );
  NAND2_X1 NAND2_2825( .ZN(N10007), .A1(N9830), .A2(N9829) );
  NAND2_X1 NAND2_2826( .ZN(N10010), .A1(N9828), .A2(N9827) );
  AND3_X1 AND3_2827( .ZN(N10013), .A1(N9791), .A2(N8307), .A3(N8269) );
  AND4_X1 AND4_2828( .ZN(N10014), .A1(N9758), .A2(N9344), .A3(N8307), .A4(N8269) );
  AND4_X1 AND5_2829_A( .ZN(extra48), .A1(N367), .A2(N9754), .A3(N9344), .A4(N8307) );
  AND2_X1 AND5_2829( .ZN(N10015), .A1(extra48), .A2(N8269) );
  AND3_X1 AND3_2830( .ZN(N10016), .A1(N9786), .A2(N8394), .A3(N8421) );
  AND4_X1 AND4_2831( .ZN(N10017), .A1(N9820), .A2(N9332), .A3(N8394), .A4(N8421) );
  AND3_X1 AND3_2832( .ZN(N10018), .A1(N9786), .A2(N8394), .A3(N8421) );
  AND4_X1 AND4_2833( .ZN(N10019), .A1(N9820), .A2(N9332), .A3(N8394), .A4(N8421) );
  AND3_X1 AND3_2834( .ZN(N10020), .A1(N9809), .A2(N8298), .A3(N8262) );
  AND4_X1 AND4_2835( .ZN(N10021), .A1(N9779), .A2(N9385), .A3(N8298), .A4(N8262) );
  AND4_X1 AND5_2836_A( .ZN(extra49), .A1(N367), .A2(N9775), .A3(N9385), .A4(N8298) );
  AND2_X1 AND5_2836( .ZN(N10022), .A1(extra49), .A2(N8262) );
  INV_X1 NOT1_2837( .ZN(N10023), .A(N9945) );
  INV_X1 NOT1_2838( .ZN(N10024), .A(N9946) );
  NAND2_X1 NAND2_2839( .ZN(N10025), .A1(N9740), .A2(N9893) );
  INV_X1 NOT1_2840( .ZN(N10026), .A(N9923) );
  INV_X1 NOT1_2841( .ZN(N10028), .A(N9924) );
  NAND2_X1 NAND2_2842( .ZN(N10032), .A1(N8595), .A2(N9897) );
  NAND2_X1 NAND2_2843( .ZN(N10033), .A1(N8598), .A2(N9899) );
  NAND2_X1 NAND2_2844( .ZN(N10034), .A1(N8601), .A2(N9901) );
  NAND2_X1 NAND2_2845( .ZN(N10035), .A1(N8604), .A2(N9903) );
  NAND2_X1 NAND2_2846( .ZN(N10036), .A1(N4803), .A2(N9906) );
  NAND2_X1 NAND2_2847( .ZN(N10037), .A1(N4806), .A2(N9908) );
  NAND2_X1 NAND2_2848( .ZN(N10038), .A1(N8627), .A2(N9910) );
  AND2_X1 AND2_2849( .ZN(N10039), .A1(N9809), .A2(N8298) );
  AND3_X1 AND3_2850( .ZN(N10040), .A1(N9779), .A2(N9385), .A3(N8298) );
  AND4_X1 AND4_2851( .ZN(N10041), .A1(N367), .A2(N9775), .A3(N9385), .A4(N8298) );
  AND2_X1 AND2_2852( .ZN(N10042), .A1(N9779), .A2(N9385) );
  AND3_X1 AND3_2853( .ZN(N10043), .A1(N367), .A2(N9775), .A3(N9385) );
  NAND2_X1 NAND2_2854( .ZN(N10050), .A1(N8727), .A2(N9938) );
  INV_X1 NOT1_2855( .ZN(N10053), .A(N9817) );
  AND2_X1 AND2_2856( .ZN(N10054), .A1(N9817), .A2(N9029) );
  AND2_X1 AND2_2857( .ZN(N10055), .A1(N9786), .A2(N8394) );
  AND3_X1 AND3_2858( .ZN(N10056), .A1(N9820), .A2(N9332), .A3(N8394) );
  AND2_X1 AND2_2859( .ZN(N10057), .A1(N9791), .A2(N8307) );
  AND3_X1 AND3_2860( .ZN(N10058), .A1(N9758), .A2(N9344), .A3(N8307) );
  AND4_X1 AND4_2861( .ZN(N10059), .A1(N367), .A2(N9754), .A3(N9344), .A4(N8307) );
  AND2_X1 AND2_2862( .ZN(N10060), .A1(N9758), .A2(N9344) );
  AND3_X1 AND3_2863( .ZN(N10061), .A1(N367), .A2(N9754), .A3(N9344) );
  NAND2_X2 NAND2_2864( .ZN(N10062), .A1(N4997), .A2(N9947) );
  NAND2_X2 NAND2_2865( .ZN(N10067), .A1(N8811), .A2(N9953) );
  NAND2_X2 NAND2_2866( .ZN(N10070), .A1(N9955), .A2(N9836) );
  NAND2_X2 NAND2_2867( .ZN(N10073), .A1(N9956), .A2(N9838) );
  NAND2_X2 NAND2_2868( .ZN(N10076), .A1(N9068), .A2(N9957) );
  NAND2_X2 NAND2_2869( .ZN(N10077), .A1(N9074), .A2(N9959) );
  NAND2_X1 NAND2_2870( .ZN(N10082), .A1(N9089), .A2(N9967) );
  NAND2_X1 NAND2_2871( .ZN(N10083), .A1(N9095), .A2(N9969) );
  NAND2_X1 NAND2_2872( .ZN(N10084), .A1(N4871), .A2(N9971) );
  NAND2_X1 NAND2_2873( .ZN(N10085), .A1(N6214), .A2(N9973) );
  NAND2_X1 NAND2_2874( .ZN(N10086), .A1(N6217), .A2(N9975) );
  NAND2_X1 NAND2_2875( .ZN(N10093), .A1(N5027), .A2(N9995) );
  NAND2_X1 NAND2_2876( .ZN(N10094), .A1(N6232), .A2(N9997) );
  OR4_X2 OR5_2877_A( .ZN(extra50), .A1(N9238), .A2(N9732), .A3(N10013), .A4(N10014) );
  OR2_X2 OR5_2877( .ZN(N10101), .A1(extra50), .A2(N10015) );
  OR4_X2 OR5_2878_A( .ZN(extra51), .A1(N9339), .A2(N9526), .A3(N10016), .A4(N10017) );
  OR2_X1 OR5_2878( .ZN(N10102), .A1(extra51), .A2(N9734) );
  OR4_X1 OR5_2879_A( .ZN(extra52), .A1(N9339), .A2(N9531), .A3(N10018), .A4(N10019) );
  OR2_X1 OR5_2879( .ZN(N10103), .A1(extra52), .A2(N9735) );
  OR4_X1 OR5_2880_A( .ZN(extra53), .A1(N9242), .A2(N9736), .A3(N10020), .A4(N10021) );
  OR2_X1 OR5_2880( .ZN(N10104), .A1(extra53), .A2(N10022) );
  AND2_X1 AND2_2881( .ZN(N10105), .A1(N9925), .A2(N9894) );
  AND2_X1 AND2_2882( .ZN(N10106), .A1(N9925), .A2(N9895) );
  AND2_X1 AND2_2883( .ZN(N10107), .A1(N9925), .A2(N9896) );
  AND2_X1 AND2_2884( .ZN(N10108), .A1(N9925), .A2(N8253) );
  NAND2_X1 NAND2_2885( .ZN(N10109), .A1(N10032), .A2(N9898) );
  NAND2_X1 NAND2_2886( .ZN(N10110), .A1(N10033), .A2(N9900) );
  NAND2_X1 NAND2_2887( .ZN(N10111), .A1(N10034), .A2(N9902) );
  NAND2_X1 NAND2_2888( .ZN(N10112), .A1(N10035), .A2(N9904) );
  NAND2_X1 NAND2_2889( .ZN(N10113), .A1(N10036), .A2(N9907) );
  NAND2_X1 NAND2_2890( .ZN(N10114), .A1(N10037), .A2(N9909) );
  NAND2_X1 NAND2_2891( .ZN(N10115), .A1(N10038), .A2(N9911) );
  OR4_X1 OR4_2892( .ZN(N10116), .A1(N9265), .A2(N10039), .A3(N10040), .A4(N10041) );
  OR3_X1 OR3_2893( .ZN(N10119), .A1(N9809), .A2(N10042), .A3(N10043) );
  INV_X1 NOT1_2894( .ZN(N10124), .A(N9925) );
  AND2_X1 AND2_2895( .ZN(N10130), .A1(N9768), .A2(N9925) );
  INV_X1 NOT1_2896( .ZN(N10131), .A(N9932) );
  INV_X1 NOT1_2897( .ZN(N10132), .A(N9935) );
  AND2_X1 AND2_2898( .ZN(N10133), .A1(N9932), .A2(N8920) );
  NAND2_X1 NAND2_2899( .ZN(N10134), .A1(N10050), .A2(N9939) );
  INV_X1 NOT1_2900( .ZN(N10135), .A(N9983) );
  NAND2_X1 NAND2_2901( .ZN(N10136), .A1(N9983), .A2(N9324) );
  INV_X1 NOT1_2902( .ZN(N10137), .A(N9986) );
  NAND2_X1 NAND2_2903( .ZN(N10138), .A1(N9986), .A2(N9784) );
  AND2_X1 AND2_2904( .ZN(N10139), .A1(N9785), .A2(N10053) );
  OR4_X1 OR4_2905( .ZN(N10140), .A1(N8943), .A2(N10055), .A3(N10056), .A4(N9790) );
  OR4_X1 OR4_2906( .ZN(N10141), .A1(N9268), .A2(N10057), .A3(N10058), .A4(N10059) );
  OR3_X1 OR3_2907( .ZN(N10148), .A1(N9791), .A2(N10060), .A3(N10061) );
  NAND2_X1 NAND2_2908( .ZN(N10155), .A1(N10062), .A2(N9948) );
  INV_X2 NOT1_2909( .ZN(N10156), .A(N9989) );
  NAND2_X1 NAND2_2910( .ZN(N10157), .A1(N9989), .A2(N9805) );
  INV_X1 NOT1_2911( .ZN(N10158), .A(N9992) );
  NAND2_X1 NAND2_2912( .ZN(N10159), .A1(N9992), .A2(N9806) );
  INV_X1 NOT1_2913( .ZN(N10160), .A(N9949) );
  NAND2_X1 NAND2_2914( .ZN(N10161), .A1(N10067), .A2(N9954) );
  INV_X1 NOT1_2915( .ZN(N10162), .A(N10007) );
  NAND2_X1 NAND2_2916( .ZN(N10163), .A1(N10007), .A2(N9825) );
  INV_X1 NOT1_2917( .ZN(N10164), .A(N10010) );
  NAND2_X1 NAND2_2918( .ZN(N10165), .A1(N10010), .A2(N9826) );
  NAND2_X1 NAND2_2919( .ZN(N10170), .A1(N10076), .A2(N9958) );
  NAND2_X1 NAND2_2920( .ZN(N10173), .A1(N10077), .A2(N9960) );
  INV_X1 NOT1_2921( .ZN(N10176), .A(N9961) );
  NAND2_X1 NAND2_2922( .ZN(N10177), .A1(N9961), .A2(N9082) );
  INV_X1 NOT1_2923( .ZN(N10178), .A(N9964) );
  NAND2_X1 NAND2_2924( .ZN(N10179), .A1(N9964), .A2(N9086) );
  NAND2_X1 NAND2_2925( .ZN(N10180), .A1(N10082), .A2(N9968) );
  NAND2_X1 NAND2_2926( .ZN(N10183), .A1(N10083), .A2(N9970) );
  NAND2_X1 NAND2_2927( .ZN(N10186), .A1(N9972), .A2(N10084) );
  NAND2_X1 NAND2_2928( .ZN(N10189), .A1(N9974), .A2(N10085) );
  NAND2_X1 NAND2_2929( .ZN(N10192), .A1(N9976), .A2(N10086) );
  INV_X1 NOT1_2930( .ZN(N10195), .A(N9979) );
  NAND2_X1 NAND2_2931( .ZN(N10196), .A1(N9979), .A2(N9982) );
  NAND2_X1 NAND2_2932( .ZN(N10197), .A1(N9996), .A2(N10093) );
  NAND2_X1 NAND2_2933( .ZN(N10200), .A1(N9998), .A2(N10094) );
  INV_X1 NOT1_2934( .ZN(N10203), .A(N9999) );
  NAND2_X1 NAND2_2935( .ZN(N10204), .A1(N9999), .A2(N10002) );
  INV_X1 NOT1_2936( .ZN(N10205), .A(N10003) );
  NAND2_X1 NAND2_2937( .ZN(N10206), .A1(N10003), .A2(N10006) );
  NAND2_X1 NAND2_2938( .ZN(N10212), .A1(N10070), .A2(N4308) );
  NAND2_X1 NAND2_2939( .ZN(N10213), .A1(N10073), .A2(N4313) );
  AND2_X2 AND2_2940( .ZN(N10230), .A1(N9774), .A2(N10131) );
  NAND2_X1 NAND2_2941( .ZN(N10231), .A1(N8730), .A2(N10135) );
  NAND2_X1 NAND2_2942( .ZN(N10232), .A1(N9478), .A2(N10137) );
  OR2_X1 OR2_2943( .ZN(N10233), .A1(N10139), .A2(N10054) );
  NAND2_X1 NAND2_2944( .ZN(N10234), .A1(N7100), .A2(N10140) );
  NAND2_X1 NAND2_2945( .ZN(N10237), .A1(N9485), .A2(N10156) );
  NAND2_X1 NAND2_2946( .ZN(N10238), .A1(N9488), .A2(N10158) );
  NAND2_X1 NAND2_2947( .ZN(N10239), .A1(N9517), .A2(N10162) );
  NAND2_X1 NAND2_2948( .ZN(N10240), .A1(N9520), .A2(N10164) );
  INV_X1 NOT1_2949( .ZN(N10241), .A(N10070) );
  INV_X1 NOT1_2950( .ZN(N10242), .A(N10073) );
  NAND2_X1 NAND2_2951( .ZN(N10247), .A1(N8146), .A2(N10176) );
  NAND2_X1 NAND2_2952( .ZN(N10248), .A1(N8156), .A2(N10178) );
  NAND2_X1 NAND2_2953( .ZN(N10259), .A1(N9692), .A2(N10195) );
  NAND2_X1 NAND2_2954( .ZN(N10264), .A1(N9717), .A2(N10203) );
  NAND2_X1 NAND2_2955( .ZN(N10265), .A1(N9723), .A2(N10205) );
  AND2_X1 AND2_2956( .ZN(N10266), .A1(N10026), .A2(N10124) );
  AND2_X1 AND2_2957( .ZN(N10267), .A1(N10028), .A2(N10124) );
  AND2_X1 AND2_2958( .ZN(N10268), .A1(N9742), .A2(N10124) );
  AND2_X1 AND2_2959( .ZN(N10269), .A1(N6923), .A2(N10124) );
  NAND2_X1 NAND2_2960( .ZN(N10270), .A1(N6762), .A2(N10116) );
  NAND2_X1 NAND2_2961( .ZN(N10271), .A1(N3061), .A2(N10241) );
  NAND2_X1 NAND2_2962( .ZN(N10272), .A1(N3064), .A2(N10242) );
  BUF_X4 BUFF1_2963( .Z(N10273), .A(N10116) );
  AND4_X1 AND5_2964_A( .ZN(extra54), .A1(N10141), .A2(N5728), .A3(N5707), .A4(N5718) );
  AND2_X1 AND5_2964( .ZN(N10278), .A1(extra54), .A2(N5697) );
  AND4_X1 AND4_2965( .ZN(N10279), .A1(N10141), .A2(N5728), .A3(N5707), .A4(N5718) );
  AND3_X1 AND3_2966( .ZN(N10280), .A1(N10141), .A2(N5728), .A3(N5718) );
  AND2_X1 AND2_2967( .ZN(N10281), .A1(N10141), .A2(N5728) );
  AND2_X1 AND2_2968( .ZN(N10282), .A1(N6784), .A2(N10141) );
  INV_X1 NOT1_2969( .ZN(N10283), .A(N10119) );
  AND4_X1 AND5_2970_A( .ZN(extra55), .A1(N10148), .A2(N5936), .A3(N5915), .A4(N5926) );
  AND2_X1 AND5_2970( .ZN(N10287), .A1(extra55), .A2(N5905) );
  AND4_X1 AND4_2971( .ZN(N10288), .A1(N10148), .A2(N5936), .A3(N5915), .A4(N5926) );
  AND3_X1 AND3_2972( .ZN(N10289), .A1(N10148), .A2(N5936), .A3(N5926) );
  AND2_X1 AND2_2973( .ZN(N10290), .A1(N10148), .A2(N5936) );
  AND2_X1 AND2_2974( .ZN(N10291), .A1(N6881), .A2(N10148) );
  AND2_X1 AND2_2975( .ZN(N10292), .A1(N8898), .A2(N10124) );
  NAND2_X1 NAND2_2976( .ZN(N10293), .A1(N10231), .A2(N10136) );
  NAND2_X1 NAND2_2977( .ZN(N10294), .A1(N10232), .A2(N10138) );
  NAND2_X1 NAND2_2978( .ZN(N10295), .A1(N8412), .A2(N10233) );
  AND2_X1 AND2_2979( .ZN(N10296), .A1(N8959), .A2(N10234) );
  NAND2_X1 NAND2_2980( .ZN(N10299), .A1(N10237), .A2(N10157) );
  NAND2_X1 NAND2_2981( .ZN(N10300), .A1(N10238), .A2(N10159) );
  OR2_X1 OR2_2982( .ZN(N10301), .A1(N10230), .A2(N10133) );
  NAND2_X1 NAND2_2983( .ZN(N10306), .A1(N10239), .A2(N10163) );
  NAND2_X1 NAND2_2984( .ZN(N10307), .A1(N10240), .A2(N10165) );
  BUF_X1 BUFF1_2985( .Z(N10308), .A(N10148) );
  BUF_X1 BUFF1_2986( .Z(N10311), .A(N10141) );
  INV_X1 NOT1_2987( .ZN(N10314), .A(N10170) );
  NAND2_X1 NAND2_2988( .ZN(N10315), .A1(N10170), .A2(N9071) );
  INV_X1 NOT1_2989( .ZN(N10316), .A(N10173) );
  NAND2_X1 NAND2_2990( .ZN(N10317), .A1(N10173), .A2(N9077) );
  NAND2_X1 NAND2_2991( .ZN(N10318), .A1(N10247), .A2(N10177) );
  NAND2_X1 NAND2_2992( .ZN(N10321), .A1(N10248), .A2(N10179) );
  INV_X1 NOT1_2993( .ZN(N10324), .A(N10180) );
  NAND2_X1 NAND2_2994( .ZN(N10325), .A1(N10180), .A2(N9092) );
  INV_X1 NOT1_2995( .ZN(N10326), .A(N10183) );
  NAND2_X1 NAND2_2996( .ZN(N10327), .A1(N10183), .A2(N9098) );
  INV_X1 NOT1_2997( .ZN(N10328), .A(N10186) );
  NAND2_X1 NAND2_2998( .ZN(N10329), .A1(N10186), .A2(N9674) );
  INV_X1 NOT1_2999( .ZN(N10330), .A(N10189) );
  NAND2_X1 NAND2_3000( .ZN(N10331), .A1(N10189), .A2(N9678) );
  INV_X2 NOT1_3001( .ZN(N10332), .A(N10192) );
  NAND2_X2 NAND2_3002( .ZN(N10333), .A1(N10192), .A2(N9977) );
  NAND2_X1 NAND2_3003( .ZN(N10334), .A1(N10259), .A2(N10196) );
  INV_X1 NOT1_3004( .ZN(N10337), .A(N10197) );
  NAND2_X1 NAND2_3005( .ZN(N10338), .A1(N10197), .A2(N9710) );
  INV_X1 NOT1_3006( .ZN(N10339), .A(N10200) );
  NAND2_X1 NAND2_3007( .ZN(N10340), .A1(N10200), .A2(N9714) );
  NAND2_X1 NAND2_3008( .ZN(N10341), .A1(N10264), .A2(N10204) );
  NAND2_X1 NAND2_3009( .ZN(N10344), .A1(N10265), .A2(N10206) );
  OR2_X1 OR2_3010( .ZN(N10350), .A1(N10266), .A2(N10105) );
  OR2_X1 OR2_3011( .ZN(N10351), .A1(N10267), .A2(N10106) );
  OR2_X1 OR2_3012( .ZN(N10352), .A1(N10268), .A2(N10107) );
  OR2_X1 OR2_3013( .ZN(N10353), .A1(N10269), .A2(N10108) );
  AND2_X1 AND2_3014( .ZN(N10354), .A1(N8857), .A2(N10270) );
  NAND2_X1 NAND2_3015( .ZN(N10357), .A1(N10271), .A2(N10212) );
  NAND2_X1 NAND2_3016( .ZN(N10360), .A1(N10272), .A2(N10213) );
  OR2_X1 OR2_3017( .ZN(N10367), .A1(N7620), .A2(N10282) );
  OR2_X1 OR2_3018( .ZN(N10375), .A1(N7671), .A2(N10291) );
  OR2_X1 OR2_3019( .ZN(N10381), .A1(N10292), .A2(N10130) );
  AND4_X1 AND4_3020( .ZN(N10388), .A1(N10114), .A2(N10134), .A3(N10293), .A4(N10294) );
  AND2_X1 AND2_3021( .ZN(N10391), .A1(N9582), .A2(N10295) );
  AND4_X1 AND4_3022( .ZN(N10399), .A1(N10113), .A2(N10115), .A3(N10299), .A4(N10300) );
  AND4_X1 AND4_3023( .ZN(N10402), .A1(N10155), .A2(N10161), .A3(N10306), .A4(N10307) );
  OR4_X2 OR5_3024_A( .ZN(extra56), .A1(N3229), .A2(N6888), .A3(N6889), .A4(N6890) );
  OR2_X2 OR5_3024( .ZN(N10406), .A1(extra56), .A2(N10287) );
  OR4_X4 OR4_3025( .ZN(N10409), .A1(N3232), .A2(N6891), .A3(N6892), .A4(N10288) );
  OR3_X1 OR3_3026( .ZN(N10412), .A1(N3236), .A2(N6893), .A3(N10289) );
  OR2_X1 OR2_3027( .ZN(N10415), .A1(N3241), .A2(N10290) );
  OR4_X1 OR5_3028_A( .ZN(extra57), .A1(N3137), .A2(N6791), .A3(N6792), .A4(N6793) );
  OR2_X1 OR5_3028( .ZN(N10419), .A1(extra57), .A2(N10278) );
  OR4_X1 OR4_3029( .ZN(N10422), .A1(N3140), .A2(N6794), .A3(N6795), .A4(N10279) );
  OR3_X1 OR3_3030( .ZN(N10425), .A1(N3144), .A2(N6796), .A3(N10280) );
  OR2_X1 OR2_3031( .ZN(N10428), .A1(N3149), .A2(N10281) );
  NAND2_X1 NAND2_3032( .ZN(N10431), .A1(N8117), .A2(N10314) );
  NAND2_X1 NAND2_3033( .ZN(N10432), .A1(N8134), .A2(N10316) );
  NAND2_X1 NAND2_3034( .ZN(N10437), .A1(N8169), .A2(N10324) );
  NAND2_X1 NAND2_3035( .ZN(N10438), .A1(N8186), .A2(N10326) );
  NAND2_X1 NAND2_3036( .ZN(N10439), .A1(N9117), .A2(N10328) );
  NAND2_X1 NAND2_3037( .ZN(N10440), .A1(N9127), .A2(N10330) );
  NAND2_X1 NAND2_3038( .ZN(N10441), .A1(N9682), .A2(N10332) );
  NAND2_X1 NAND2_3039( .ZN(N10444), .A1(N9183), .A2(N10337) );
  NAND2_X1 NAND2_3040( .ZN(N10445), .A1(N9193), .A2(N10339) );
  INV_X1 NOT1_3041( .ZN(N10450), .A(N10296) );
  AND2_X1 AND2_3042( .ZN(N10451), .A1(N10296), .A2(N4193) );
  INV_X1 NOT1_3043( .ZN(N10455), .A(N10308) );
  NAND2_X1 NAND2_3044( .ZN(N10456), .A1(N10308), .A2(N8242) );
  INV_X1 NOT1_3045( .ZN(N10465), .A(N10311) );
  NAND2_X1 NAND2_3046( .ZN(N10466), .A1(N10311), .A2(N8247) );
  INV_X1 NOT1_3047( .ZN(N10479), .A(N10273) );
  INV_X1 NOT1_3048( .ZN(N10497), .A(N10301) );
  NAND2_X1 NAND2_3049( .ZN(N10509), .A1(N10431), .A2(N10315) );
  NAND2_X1 NAND2_3050( .ZN(N10512), .A1(N10432), .A2(N10317) );
  INV_X1 NOT1_3051( .ZN(N10515), .A(N10318) );
  NAND2_X1 NAND2_3052( .ZN(N10516), .A1(N10318), .A2(N8632) );
  INV_X1 NOT1_3053( .ZN(N10517), .A(N10321) );
  NAND2_X1 NAND2_3054( .ZN(N10518), .A1(N10321), .A2(N8637) );
  NAND2_X1 NAND2_3055( .ZN(N10519), .A1(N10437), .A2(N10325) );
  NAND2_X1 NAND2_3056( .ZN(N10522), .A1(N10438), .A2(N10327) );
  NAND2_X1 NAND2_3057( .ZN(N10525), .A1(N10439), .A2(N10329) );
  NAND2_X1 NAND2_3058( .ZN(N10528), .A1(N10440), .A2(N10331) );
  NAND2_X1 NAND2_3059( .ZN(N10531), .A1(N10441), .A2(N10333) );
  INV_X1 NOT1_3060( .ZN(N10534), .A(N10334) );
  NAND2_X1 NAND2_3061( .ZN(N10535), .A1(N10334), .A2(N9695) );
  NAND2_X1 NAND2_3062( .ZN(N10536), .A1(N10444), .A2(N10338) );
  NAND2_X1 NAND2_3063( .ZN(N10539), .A1(N10445), .A2(N10340) );
  INV_X1 NOT1_3064( .ZN(N10542), .A(N10341) );
  NAND2_X1 NAND2_3065( .ZN(N10543), .A1(N10341), .A2(N9720) );
  INV_X1 NOT1_3066( .ZN(N10544), .A(N10344) );
  NAND2_X1 NAND2_3067( .ZN(N10545), .A1(N10344), .A2(N9726) );
  AND2_X1 AND2_3068( .ZN(N10546), .A1(N5631), .A2(N10450) );
  INV_X1 NOT1_3069( .ZN(N10547), .A(N10391) );
  AND2_X1 AND2_3070( .ZN(N10548), .A1(N10391), .A2(N8950) );
  AND2_X1 AND2_3071( .ZN(N10549), .A1(N5165), .A2(N10367) );
  INV_X1 NOT1_3072( .ZN(N10550), .A(N10354) );
  AND2_X2 AND2_3073( .ZN(N10551), .A1(N10354), .A2(N3126) );
  NAND2_X1 NAND2_3074( .ZN(N10552), .A1(N7411), .A2(N10455) );
  AND2_X1 AND2_3075( .ZN(N10553), .A1(N10375), .A2(N9539) );
  AND2_X1 AND2_3076( .ZN(N10554), .A1(N10375), .A2(N9540) );
  AND2_X1 AND2_3077( .ZN(N10555), .A1(N10375), .A2(N9541) );
  AND2_X1 AND2_3078( .ZN(N10556), .A1(N10375), .A2(N6761) );
  INV_X1 NOT1_3079( .ZN(N10557), .A(N10406) );
  NAND2_X1 NAND2_3080( .ZN(N10558), .A1(N10406), .A2(N8243) );
  INV_X1 NOT1_3081( .ZN(N10559), .A(N10409) );
  NAND2_X1 NAND2_3082( .ZN(N10560), .A1(N10409), .A2(N8244) );
  INV_X1 NOT1_3083( .ZN(N10561), .A(N10412) );
  NAND2_X1 NAND2_3084( .ZN(N10562), .A1(N10412), .A2(N8245) );
  INV_X1 NOT1_3085( .ZN(N10563), .A(N10415) );
  NAND2_X1 NAND2_3086( .ZN(N10564), .A1(N10415), .A2(N8246) );
  NAND2_X1 NAND2_3087( .ZN(N10565), .A1(N7426), .A2(N10465) );
  INV_X1 NOT1_3088( .ZN(N10566), .A(N10419) );
  NAND2_X1 NAND2_3089( .ZN(N10567), .A1(N10419), .A2(N8248) );
  INV_X1 NOT1_3090( .ZN(N10568), .A(N10422) );
  NAND2_X1 NAND2_3091( .ZN(N10569), .A1(N10422), .A2(N8249) );
  INV_X1 NOT1_3092( .ZN(N10570), .A(N10425) );
  NAND2_X1 NAND2_3093( .ZN(N10571), .A1(N10425), .A2(N8250) );
  INV_X2 NOT1_3094( .ZN(N10572), .A(N10428) );
  NAND2_X1 NAND2_3095( .ZN(N10573), .A1(N10428), .A2(N8251) );
  INV_X1 NOT1_3096( .ZN(N10574), .A(N10399) );
  INV_X1 NOT1_3097( .ZN(N10575), .A(N10402) );
  INV_X1 NOT1_3098( .ZN(N10576), .A(N10388) );
  AND3_X1 AND3_3099( .ZN(N10577), .A1(N10399), .A2(N10402), .A3(N10388) );
  AND3_X1 AND3_3100( .ZN(N10581), .A1(N10360), .A2(N9543), .A3(N10273) );
  AND3_X1 AND3_3101( .ZN(N10582), .A1(N10357), .A2(N9905), .A3(N10273) );
  INV_X1 NOT1_3102( .ZN(N10583), .A(N10367) );
  AND2_X1 AND2_3103( .ZN(N10587), .A1(N10367), .A2(N5735) );
  AND2_X1 AND2_3104( .ZN(N10588), .A1(N10367), .A2(N3135) );
  INV_X1 NOT1_3105( .ZN(N10589), .A(N10375) );
  AND4_X1 AND5_3106_A( .ZN(extra58), .A1(N10381), .A2(N7180), .A3(N7159), .A4(N7170) );
  AND2_X1 AND5_3106( .ZN(N10594), .A1(extra58), .A2(N7149) );
  AND4_X1 AND4_3107( .ZN(N10595), .A1(N10381), .A2(N7180), .A3(N7159), .A4(N7170) );
  AND3_X1 AND3_3108( .ZN(N10596), .A1(N10381), .A2(N7180), .A3(N7170) );
  AND2_X1 AND2_3109( .ZN(N10597), .A1(N10381), .A2(N7180) );
  AND2_X1 AND2_3110( .ZN(N10598), .A1(N8444), .A2(N10381) );
  BUF_X4 BUFF1_3111( .Z(N10602), .A(N10381) );
  NAND2_X1 NAND2_3112( .ZN(N10609), .A1(N7479), .A2(N10515) );
  NAND2_X1 NAND2_3113( .ZN(N10610), .A1(N7491), .A2(N10517) );
  NAND2_X1 NAND2_3114( .ZN(N10621), .A1(N9149), .A2(N10534) );
  NAND2_X1 NAND2_3115( .ZN(N10626), .A1(N9206), .A2(N10542) );
  NAND2_X1 NAND2_3116( .ZN(N10627), .A1(N9223), .A2(N10544) );
  OR2_X1 OR2_3117( .ZN(N10628), .A1(N10546), .A2(N10451) );
  AND2_X1 AND2_3118( .ZN(N10629), .A1(N9733), .A2(N10547) );
  AND2_X1 AND2_3119( .ZN(N10631), .A1(N5166), .A2(N10550) );
  NAND2_X1 NAND2_3120( .ZN(N10632), .A1(N10552), .A2(N10456) );
  NAND2_X1 NAND2_3121( .ZN(N10637), .A1(N7414), .A2(N10557) );
  NAND2_X1 NAND2_3122( .ZN(N10638), .A1(N7417), .A2(N10559) );
  NAND2_X1 NAND2_3123( .ZN(N10639), .A1(N7420), .A2(N10561) );
  NAND2_X1 NAND2_3124( .ZN(N10640), .A1(N7423), .A2(N10563) );
  NAND2_X1 NAND2_3125( .ZN(N10641), .A1(N10565), .A2(N10466) );
  NAND2_X1 NAND2_3126( .ZN(N10642), .A1(N7429), .A2(N10566) );
  NAND2_X1 NAND2_3127( .ZN(N10643), .A1(N7432), .A2(N10568) );
  NAND2_X1 NAND2_3128( .ZN(N10644), .A1(N7435), .A2(N10570) );
  NAND2_X1 NAND2_3129( .ZN(N10645), .A1(N7438), .A2(N10572) );
  AND3_X1 AND3_3130( .ZN(N10647), .A1(N886), .A2(N887), .A3(N10577) );
  AND3_X1 AND3_3131( .ZN(N10648), .A1(N10360), .A2(N8857), .A3(N10479) );
  AND3_X1 AND3_3132( .ZN(N10649), .A1(N10357), .A2(N7609), .A3(N10479) );
  OR2_X1 OR2_3133( .ZN(N10652), .A1(N8966), .A2(N10598) );
  OR4_X1 OR5_3134_A( .ZN(extra59), .A1(N4675), .A2(N8451), .A3(N8452), .A4(N8453) );
  OR2_X1 OR5_3134( .ZN(N10659), .A1(extra59), .A2(N10594) );
  OR4_X1 OR4_3135( .ZN(N10662), .A1(N4678), .A2(N8454), .A3(N8455), .A4(N10595) );
  OR3_X1 OR3_3136( .ZN(N10665), .A1(N4682), .A2(N8456), .A3(N10596) );
  OR2_X1 OR2_3137( .ZN(N10668), .A1(N4687), .A2(N10597) );
  INV_X1 NOT1_3138( .ZN(N10671), .A(N10509) );
  NAND2_X1 NAND2_3139( .ZN(N10672), .A1(N10509), .A2(N8615) );
  INV_X1 NOT1_3140( .ZN(N10673), .A(N10512) );
  NAND2_X1 NAND2_3141( .ZN(N10674), .A1(N10512), .A2(N8624) );
  NAND2_X1 NAND2_3142( .ZN(N10675), .A1(N10609), .A2(N10516) );
  NAND2_X1 NAND2_3143( .ZN(N10678), .A1(N10610), .A2(N10518) );
  INV_X1 NOT1_3144( .ZN(N10681), .A(N10519) );
  NAND2_X2 NAND2_3145( .ZN(N10682), .A1(N10519), .A2(N8644) );
  INV_X1 NOT1_3146( .ZN(N10683), .A(N10522) );
  NAND2_X1 NAND2_3147( .ZN(N10684), .A1(N10522), .A2(N8653) );
  INV_X1 NOT1_3148( .ZN(N10685), .A(N10525) );
  NAND2_X1 NAND2_3149( .ZN(N10686), .A1(N10525), .A2(N9454) );
  INV_X1 NOT1_3150( .ZN(N10687), .A(N10528) );
  NAND2_X1 NAND2_3151( .ZN(N10688), .A1(N10528), .A2(N9459) );
  INV_X1 NOT1_3152( .ZN(N10689), .A(N10531) );
  NAND2_X1 NAND2_3153( .ZN(N10690), .A1(N10531), .A2(N9978) );
  NAND2_X1 NAND2_3154( .ZN(N10691), .A1(N10621), .A2(N10535) );
  INV_X1 NOT1_3155( .ZN(N10694), .A(N10536) );
  NAND2_X1 NAND2_3156( .ZN(N10695), .A1(N10536), .A2(N9493) );
  INV_X1 NOT1_3157( .ZN(N10696), .A(N10539) );
  NAND2_X1 NAND2_3158( .ZN(N10697), .A1(N10539), .A2(N9498) );
  NAND2_X1 NAND2_3159( .ZN(N10698), .A1(N10626), .A2(N10543) );
  NAND2_X1 NAND2_3160( .ZN(N10701), .A1(N10627), .A2(N10545) );
  OR2_X1 OR2_3161( .ZN(N10704), .A1(N10629), .A2(N10548) );
  AND2_X1 AND2_3162( .ZN(N10705), .A1(N3159), .A2(N10583) );
  OR2_X1 OR2_3163( .ZN(N10706), .A1(N10631), .A2(N10551) );
  AND2_X1 AND2_3164( .ZN(N10707), .A1(N9737), .A2(N10589) );
  AND2_X1 AND2_3165( .ZN(N10708), .A1(N9738), .A2(N10589) );
  AND2_X1 AND2_3166( .ZN(N10709), .A1(N9243), .A2(N10589) );
  AND2_X1 AND2_3167( .ZN(N10710), .A1(N5892), .A2(N10589) );
  NAND2_X1 NAND2_3168( .ZN(N10711), .A1(N10637), .A2(N10558) );
  NAND2_X1 NAND2_3169( .ZN(N10712), .A1(N10638), .A2(N10560) );
  NAND2_X1 NAND2_3170( .ZN(N10713), .A1(N10639), .A2(N10562) );
  NAND2_X1 NAND2_3171( .ZN(N10714), .A1(N10640), .A2(N10564) );
  NAND2_X1 NAND2_3172( .ZN(N10715), .A1(N10642), .A2(N10567) );
  NAND2_X1 NAND2_3173( .ZN(N10716), .A1(N10643), .A2(N10569) );
  NAND2_X1 NAND2_3174( .ZN(N10717), .A1(N10644), .A2(N10571) );
  NAND2_X1 NAND2_3175( .ZN(N10718), .A1(N10645), .A2(N10573) );
  INV_X1 NOT1_3176( .ZN(N10719), .A(N10602) );
  NAND2_X1 NAND2_3177( .ZN(N10720), .A1(N10602), .A2(N9244) );
  INV_X1 NOT1_3178( .ZN(N10729), .A(N10647) );
  AND2_X1 AND2_3179( .ZN(N10730), .A1(N5178), .A2(N10583) );
  AND2_X1 AND2_3180( .ZN(N10731), .A1(N2533), .A2(N10583) );
  NAND2_X1 NAND2_3181( .ZN(N10737), .A1(N7447), .A2(N10671) );
  NAND2_X1 NAND2_3182( .ZN(N10738), .A1(N7465), .A2(N10673) );
  OR4_X2 OR4_3183( .ZN(N10739), .A1(N10648), .A2(N10649), .A3(N10581), .A4(N10582) );
  NAND2_X1 NAND2_3184( .ZN(N10746), .A1(N7503), .A2(N10681) );
  NAND2_X1 NAND2_3185( .ZN(N10747), .A1(N7521), .A2(N10683) );
  NAND2_X1 NAND2_3186( .ZN(N10748), .A1(N8678), .A2(N10685) );
  NAND2_X1 NAND2_3187( .ZN(N10749), .A1(N8690), .A2(N10687) );
  NAND2_X1 NAND2_3188( .ZN(N10750), .A1(N9685), .A2(N10689) );
  NAND2_X1 NAND2_3189( .ZN(N10753), .A1(N8757), .A2(N10694) );
  NAND2_X1 NAND2_3190( .ZN(N10754), .A1(N8769), .A2(N10696) );
  OR2_X1 OR2_3191( .ZN(N10759), .A1(N10705), .A2(N10549) );
  OR2_X1 OR2_3192( .ZN(N10760), .A1(N10707), .A2(N10553) );
  OR2_X1 OR2_3193( .ZN(N10761), .A1(N10708), .A2(N10554) );
  OR2_X1 OR2_3194( .ZN(N10762), .A1(N10709), .A2(N10555) );
  OR2_X1 OR2_3195( .ZN(N10763), .A1(N10710), .A2(N10556) );
  NAND2_X1 NAND2_3196( .ZN(N10764), .A1(N8580), .A2(N10719) );
  AND2_X1 AND2_3197( .ZN(N10765), .A1(N10652), .A2(N9890) );
  AND2_X1 AND2_3198( .ZN(N10766), .A1(N10652), .A2(N9891) );
  AND2_X1 AND2_3199( .ZN(N10767), .A1(N10652), .A2(N9892) );
  AND2_X1 AND2_3200( .ZN(N10768), .A1(N10652), .A2(N8252) );
  INV_X2 NOT1_3201( .ZN(N10769), .A(N10659) );
  NAND2_X1 NAND2_3202( .ZN(N10770), .A1(N10659), .A2(N9245) );
  INV_X1 NOT1_3203( .ZN(N10771), .A(N10662) );
  NAND2_X1 NAND2_3204( .ZN(N10772), .A1(N10662), .A2(N9246) );
  INV_X1 NOT1_3205( .ZN(N10773), .A(N10665) );
  NAND2_X1 NAND2_3206( .ZN(N10774), .A1(N10665), .A2(N9247) );
  INV_X1 NOT1_3207( .ZN(N10775), .A(N10668) );
  NAND2_X1 NAND2_3208( .ZN(N10776), .A1(N10668), .A2(N9248) );
  OR2_X1 OR2_3209( .ZN(N10778), .A1(N10730), .A2(N10587) );
  OR2_X1 OR2_3210( .ZN(N10781), .A1(N10731), .A2(N10588) );
  INV_X1 NOT1_3211( .ZN(N10784), .A(N10652) );
  NAND2_X1 NAND2_3212( .ZN(N10789), .A1(N10737), .A2(N10672) );
  NAND2_X1 NAND2_3213( .ZN(N10792), .A1(N10738), .A2(N10674) );
  INV_X1 NOT1_3214( .ZN(N10796), .A(N10675) );
  NAND2_X1 NAND2_3215( .ZN(N10797), .A1(N10675), .A2(N8633) );
  INV_X1 NOT1_3216( .ZN(N10798), .A(N10678) );
  NAND2_X1 NAND2_3217( .ZN(N10799), .A1(N10678), .A2(N8638) );
  NAND2_X1 NAND2_3218( .ZN(N10800), .A1(N10746), .A2(N10682) );
  NAND2_X1 NAND2_3219( .ZN(N10803), .A1(N10747), .A2(N10684) );
  NAND2_X1 NAND2_3220( .ZN(N10806), .A1(N10748), .A2(N10686) );
  NAND2_X1 NAND2_3221( .ZN(N10809), .A1(N10749), .A2(N10688) );
  NAND2_X1 NAND2_3222( .ZN(N10812), .A1(N10750), .A2(N10690) );
  INV_X1 NOT1_3223( .ZN(N10815), .A(N10691) );
  NAND2_X1 NAND2_3224( .ZN(N10816), .A1(N10691), .A2(N9866) );
  NAND2_X1 NAND2_3225( .ZN(N10817), .A1(N10753), .A2(N10695) );
  NAND2_X1 NAND2_3226( .ZN(N10820), .A1(N10754), .A2(N10697) );
  INV_X1 NOT1_3227( .ZN(N10823), .A(N10698) );
  NAND2_X1 NAND2_3228( .ZN(N10824), .A1(N10698), .A2(N9505) );
  INV_X1 NOT1_3229( .ZN(N10825), .A(N10701) );
  NAND2_X1 NAND2_3230( .ZN(N10826), .A1(N10701), .A2(N9514) );
  NAND2_X1 NAND2_3231( .ZN(N10827), .A1(N10764), .A2(N10720) );
  NAND2_X1 NAND2_3232( .ZN(N10832), .A1(N8583), .A2(N10769) );
  NAND2_X1 NAND2_3233( .ZN(N10833), .A1(N8586), .A2(N10771) );
  NAND2_X1 NAND2_3234( .ZN(N10834), .A1(N8589), .A2(N10773) );
  NAND2_X1 NAND2_3235( .ZN(N10835), .A1(N8592), .A2(N10775) );
  INV_X1 NOT1_3236( .ZN(N10836), .A(N10739) );
  BUF_X4 BUFF1_3237( .Z(N10837), .A(N10778) );
  BUF_X4 BUFF1_3238( .Z(N10838), .A(N10778) );
  BUF_X1 BUFF1_3239( .Z(N10839), .A(N10781) );
  BUF_X1 BUFF1_3240( .Z(N10840), .A(N10781) );
  NAND2_X1 NAND2_3241( .ZN(N10845), .A1(N7482), .A2(N10796) );
  NAND2_X1 NAND2_3242( .ZN(N10846), .A1(N7494), .A2(N10798) );
  NAND2_X1 NAND2_3243( .ZN(N10857), .A1(N9473), .A2(N10815) );
  NAND2_X1 NAND2_3244( .ZN(N10862), .A1(N8781), .A2(N10823) );
  NAND2_X1 NAND2_3245( .ZN(N10863), .A1(N8799), .A2(N10825) );
  AND2_X1 AND2_3246( .ZN(N10864), .A1(N10023), .A2(N10784) );
  AND2_X1 AND2_3247( .ZN(N10865), .A1(N10024), .A2(N10784) );
  AND2_X1 AND2_3248( .ZN(N10866), .A1(N9739), .A2(N10784) );
  AND2_X1 AND2_3249( .ZN(N10867), .A1(N7136), .A2(N10784) );
  NAND2_X1 NAND2_3250( .ZN(N10868), .A1(N10832), .A2(N10770) );
  NAND2_X1 NAND2_3251( .ZN(N10869), .A1(N10833), .A2(N10772) );
  NAND2_X1 NAND2_3252( .ZN(N10870), .A1(N10834), .A2(N10774) );
  NAND2_X1 NAND2_3253( .ZN(N10871), .A1(N10835), .A2(N10776) );
  INV_X1 NOT1_3254( .ZN(N10872), .A(N10789) );
  NAND2_X1 NAND2_3255( .ZN(N10873), .A1(N10789), .A2(N8616) );
  INV_X1 NOT1_3256( .ZN(N10874), .A(N10792) );
  NAND2_X1 NAND2_3257( .ZN(N10875), .A1(N10792), .A2(N8625) );
  NAND2_X1 NAND2_3258( .ZN(N10876), .A1(N10845), .A2(N10797) );
  NAND2_X1 NAND2_3259( .ZN(N10879), .A1(N10846), .A2(N10799) );
  INV_X1 NOT1_3260( .ZN(N10882), .A(N10800) );
  NAND2_X1 NAND2_3261( .ZN(N10883), .A1(N10800), .A2(N8645) );
  INV_X1 NOT1_3262( .ZN(N10884), .A(N10803) );
  NAND2_X1 NAND2_3263( .ZN(N10885), .A1(N10803), .A2(N8654) );
  INV_X1 NOT1_3264( .ZN(N10886), .A(N10806) );
  NAND2_X1 NAND2_3265( .ZN(N10887), .A1(N10806), .A2(N9455) );
  INV_X1 NOT1_3266( .ZN(N10888), .A(N10809) );
  NAND2_X1 NAND2_3267( .ZN(N10889), .A1(N10809), .A2(N9460) );
  INV_X1 NOT1_3268( .ZN(N10890), .A(N10812) );
  NAND2_X1 NAND2_3269( .ZN(N10891), .A1(N10812), .A2(N9862) );
  NAND2_X1 NAND2_3270( .ZN(N10892), .A1(N10857), .A2(N10816) );
  INV_X1 NOT1_3271( .ZN(N10895), .A(N10817) );
  NAND2_X1 NAND2_3272( .ZN(N10896), .A1(N10817), .A2(N9494) );
  INV_X1 NOT1_3273( .ZN(N10897), .A(N10820) );
  NAND2_X1 NAND2_3274( .ZN(N10898), .A1(N10820), .A2(N9499) );
  NAND2_X1 NAND2_3275( .ZN(N10899), .A1(N10862), .A2(N10824) );
  NAND2_X1 NAND2_3276( .ZN(N10902), .A1(N10863), .A2(N10826) );
  OR2_X1 OR2_3277( .ZN(N10905), .A1(N10864), .A2(N10765) );
  OR2_X1 OR2_3278( .ZN(N10906), .A1(N10865), .A2(N10766) );
  OR2_X1 OR2_3279( .ZN(N10907), .A1(N10866), .A2(N10767) );
  OR2_X1 OR2_3280( .ZN(N10908), .A1(N10867), .A2(N10768) );
  NAND2_X1 NAND2_3281( .ZN(N10909), .A1(N7450), .A2(N10872) );
  NAND2_X1 NAND2_3282( .ZN(N10910), .A1(N7468), .A2(N10874) );
  NAND2_X1 NAND2_3283( .ZN(N10915), .A1(N7506), .A2(N10882) );
  NAND2_X2 NAND2_3284( .ZN(N10916), .A1(N7524), .A2(N10884) );
  NAND2_X2 NAND2_3285( .ZN(N10917), .A1(N8681), .A2(N10886) );
  NAND2_X1 NAND2_3286( .ZN(N10918), .A1(N8693), .A2(N10888) );
  NAND2_X1 NAND2_3287( .ZN(N10919), .A1(N9462), .A2(N10890) );
  NAND2_X1 NAND2_3288( .ZN(N10922), .A1(N8760), .A2(N10895) );
  NAND2_X1 NAND2_3289( .ZN(N10923), .A1(N8772), .A2(N10897) );
  NAND2_X1 NAND2_3290( .ZN(N10928), .A1(N10909), .A2(N10873) );
  NAND2_X1 NAND2_3291( .ZN(N10931), .A1(N10910), .A2(N10875) );
  INV_X2 NOT1_3292( .ZN(N10934), .A(N10876) );
  NAND2_X1 NAND2_3293( .ZN(N10935), .A1(N10876), .A2(N8634) );
  INV_X1 NOT1_3294( .ZN(N10936), .A(N10879) );
  NAND2_X1 NAND2_3295( .ZN(N10937), .A1(N10879), .A2(N8639) );
  NAND2_X1 NAND2_3296( .ZN(N10938), .A1(N10915), .A2(N10883) );
  NAND2_X1 NAND2_3297( .ZN(N10941), .A1(N10916), .A2(N10885) );
  NAND2_X1 NAND2_3298( .ZN(N10944), .A1(N10917), .A2(N10887) );
  NAND2_X1 NAND2_3299( .ZN(N10947), .A1(N10918), .A2(N10889) );
  NAND2_X1 NAND2_3300( .ZN(N10950), .A1(N10919), .A2(N10891) );
  INV_X1 NOT1_3301( .ZN(N10953), .A(N10892) );
  NAND2_X1 NAND2_3302( .ZN(N10954), .A1(N10892), .A2(N9476) );
  NAND2_X1 NAND2_3303( .ZN(N10955), .A1(N10922), .A2(N10896) );
  NAND2_X1 NAND2_3304( .ZN(N10958), .A1(N10923), .A2(N10898) );
  INV_X1 NOT1_3305( .ZN(N10961), .A(N10899) );
  NAND2_X1 NAND2_3306( .ZN(N10962), .A1(N10899), .A2(N9506) );
  INV_X1 NOT1_3307( .ZN(N10963), .A(N10902) );
  NAND2_X1 NAND2_3308( .ZN(N10964), .A1(N10902), .A2(N9515) );
  NAND2_X1 NAND2_3309( .ZN(N10969), .A1(N7485), .A2(N10934) );
  NAND2_X1 NAND2_3310( .ZN(N10970), .A1(N7497), .A2(N10936) );
  NAND2_X1 NAND2_3311( .ZN(N10981), .A1(N8718), .A2(N10953) );
  NAND2_X1 NAND2_3312( .ZN(N10986), .A1(N8784), .A2(N10961) );
  NAND2_X1 NAND2_3313( .ZN(N10987), .A1(N8802), .A2(N10963) );
  INV_X1 NOT1_3314( .ZN(N10988), .A(N10928) );
  NAND2_X1 NAND2_3315( .ZN(N10989), .A1(N10928), .A2(N8617) );
  INV_X1 NOT1_3316( .ZN(N10990), .A(N10931) );
  NAND2_X1 NAND2_3317( .ZN(N10991), .A1(N10931), .A2(N8626) );
  NAND2_X1 NAND2_3318( .ZN(N10992), .A1(N10969), .A2(N10935) );
  NAND2_X1 NAND2_3319( .ZN(N10995), .A1(N10970), .A2(N10937) );
  INV_X1 NOT1_3320( .ZN(N10998), .A(N10938) );
  NAND2_X1 NAND2_3321( .ZN(N10999), .A1(N10938), .A2(N8646) );
  INV_X1 NOT1_3322( .ZN(N11000), .A(N10941) );
  NAND2_X1 NAND2_3323( .ZN(N11001), .A1(N10941), .A2(N8655) );
  INV_X1 NOT1_3324( .ZN(N11002), .A(N10944) );
  NAND2_X1 NAND2_3325( .ZN(N11003), .A1(N10944), .A2(N9456) );
  INV_X1 NOT1_3326( .ZN(N11004), .A(N10947) );
  NAND2_X1 NAND2_3327( .ZN(N11005), .A1(N10947), .A2(N9461) );
  INV_X1 NOT1_3328( .ZN(N11006), .A(N10950) );
  NAND2_X1 NAND2_3329( .ZN(N11007), .A1(N10950), .A2(N9465) );
  NAND2_X1 NAND2_3330( .ZN(N11008), .A1(N10981), .A2(N10954) );
  INV_X1 NOT1_3331( .ZN(N11011), .A(N10955) );
  NAND2_X1 NAND2_3332( .ZN(N11012), .A1(N10955), .A2(N9495) );
  INV_X1 NOT1_3333( .ZN(N11013), .A(N10958) );
  NAND2_X1 NAND2_3334( .ZN(N11014), .A1(N10958), .A2(N9500) );
  NAND2_X1 NAND2_3335( .ZN(N11015), .A1(N10986), .A2(N10962) );
  NAND2_X1 NAND2_3336( .ZN(N11018), .A1(N10987), .A2(N10964) );
  NAND2_X1 NAND2_3337( .ZN(N11023), .A1(N7453), .A2(N10988) );
  NAND2_X1 NAND2_3338( .ZN(N11024), .A1(N7471), .A2(N10990) );
  NAND2_X1 NAND2_3339( .ZN(N11027), .A1(N7509), .A2(N10998) );
  NAND2_X1 NAND2_3340( .ZN(N11028), .A1(N7527), .A2(N11000) );
  NAND2_X1 NAND2_3341( .ZN(N11029), .A1(N8684), .A2(N11002) );
  NAND2_X1 NAND2_3342( .ZN(N11030), .A1(N8696), .A2(N11004) );
  NAND2_X1 NAND2_3343( .ZN(N11031), .A1(N8702), .A2(N11006) );
  NAND2_X1 NAND2_3344( .ZN(N11034), .A1(N8763), .A2(N11011) );
  NAND2_X1 NAND2_3345( .ZN(N11035), .A1(N8775), .A2(N11013) );
  INV_X1 NOT1_3346( .ZN(N11040), .A(N10992) );
  NAND2_X1 NAND2_3347( .ZN(N11041), .A1(N10992), .A2(N8294) );
  INV_X1 NOT1_3348( .ZN(N11042), .A(N10995) );
  NAND2_X1 NAND2_3349( .ZN(N11043), .A1(N10995), .A2(N8295) );
  NAND2_X1 NAND2_3350( .ZN(N11044), .A1(N11023), .A2(N10989) );
  NAND2_X1 NAND2_3351( .ZN(N11047), .A1(N11024), .A2(N10991) );
  NAND2_X1 NAND2_3352( .ZN(N11050), .A1(N11027), .A2(N10999) );
  NAND2_X1 NAND2_3353( .ZN(N11053), .A1(N11028), .A2(N11001) );
  NAND2_X1 NAND2_3354( .ZN(N11056), .A1(N11029), .A2(N11003) );
  NAND2_X1 NAND2_3355( .ZN(N11059), .A1(N11030), .A2(N11005) );
  NAND2_X1 NAND2_3356( .ZN(N11062), .A1(N11031), .A2(N11007) );
  INV_X1 NOT1_3357( .ZN(N11065), .A(N11008) );
  NAND2_X1 NAND2_3358( .ZN(N11066), .A1(N11008), .A2(N9477) );
  NAND2_X1 NAND2_3359( .ZN(N11067), .A1(N11034), .A2(N11012) );
  NAND2_X1 NAND2_3360( .ZN(N11070), .A1(N11035), .A2(N11014) );
  INV_X1 NOT1_3361( .ZN(N11073), .A(N11015) );
  NAND2_X1 NAND2_3362( .ZN(N11074), .A1(N11015), .A2(N9507) );
  INV_X1 NOT1_3363( .ZN(N11075), .A(N11018) );
  NAND2_X1 NAND2_3364( .ZN(N11076), .A1(N11018), .A2(N9516) );
  NAND2_X1 NAND2_3365( .ZN(N11077), .A1(N7488), .A2(N11040) );
  NAND2_X1 NAND2_3366( .ZN(N11078), .A1(N7500), .A2(N11042) );
  NAND2_X1 NAND2_3367( .ZN(N11095), .A1(N8721), .A2(N11065) );
  NAND2_X1 NAND2_3368( .ZN(N11098), .A1(N8787), .A2(N11073) );
  NAND2_X1 NAND2_3369( .ZN(N11099), .A1(N8805), .A2(N11075) );
  NAND2_X1 NAND2_3370( .ZN(N11100), .A1(N11077), .A2(N11041) );
  NAND2_X1 NAND2_3371( .ZN(N11103), .A1(N11078), .A2(N11043) );
  INV_X1 NOT1_3372( .ZN(N11106), .A(N11056) );
  NAND2_X1 NAND2_3373( .ZN(N11107), .A1(N11056), .A2(N9319) );
  INV_X1 NOT1_3374( .ZN(N11108), .A(N11059) );
  NAND2_X1 NAND2_3375( .ZN(N11109), .A1(N11059), .A2(N9320) );
  INV_X1 NOT1_3376( .ZN(N11110), .A(N11067) );
  NAND2_X1 NAND2_3377( .ZN(N11111), .A1(N11067), .A2(N9381) );
  INV_X1 NOT1_3378( .ZN(N11112), .A(N11070) );
  NAND2_X1 NAND2_3379( .ZN(N11113), .A1(N11070), .A2(N9382) );
  INV_X2 NOT1_3380( .ZN(N11114), .A(N11044) );
  NAND2_X1 NAND2_3381( .ZN(N11115), .A1(N11044), .A2(N8618) );
  INV_X1 NOT1_3382( .ZN(N11116), .A(N11047) );
  NAND2_X1 NAND2_3383( .ZN(N11117), .A1(N11047), .A2(N8619) );
  INV_X1 NOT1_3384( .ZN(N11118), .A(N11050) );
  NAND2_X1 NAND2_3385( .ZN(N11119), .A1(N11050), .A2(N8647) );
  INV_X1 NOT1_3386( .ZN(N11120), .A(N11053) );
  NAND2_X1 NAND2_3387( .ZN(N11121), .A1(N11053), .A2(N8648) );
  INV_X1 NOT1_3388( .ZN(N11122), .A(N11062) );
  NAND2_X1 NAND2_3389( .ZN(N11123), .A1(N11062), .A2(N9466) );
  NAND2_X1 NAND2_3390( .ZN(N11124), .A1(N11095), .A2(N11066) );
  NAND2_X1 NAND2_3391( .ZN(N11127), .A1(N11098), .A2(N11074) );
  NAND2_X1 NAND2_3392( .ZN(N11130), .A1(N11099), .A2(N11076) );
  NAND2_X1 NAND2_3393( .ZN(N11137), .A1(N8687), .A2(N11106) );
  NAND2_X1 NAND2_3394( .ZN(N11138), .A1(N8699), .A2(N11108) );
  NAND2_X1 NAND2_3395( .ZN(N11139), .A1(N8766), .A2(N11110) );
  NAND2_X1 NAND2_3396( .ZN(N11140), .A1(N8778), .A2(N11112) );
  NAND2_X1 NAND2_3397( .ZN(N11141), .A1(N7456), .A2(N11114) );
  NAND2_X1 NAND2_3398( .ZN(N11142), .A1(N7474), .A2(N11116) );
  NAND2_X1 NAND2_3399( .ZN(N11143), .A1(N7512), .A2(N11118) );
  NAND2_X1 NAND2_3400( .ZN(N11144), .A1(N7530), .A2(N11120) );
  NAND2_X1 NAND2_3401( .ZN(N11145), .A1(N8705), .A2(N11122) );
  AND3_X1 AND3_3402( .ZN(N11152), .A1(N11103), .A2(N8871), .A3(N10283) );
  AND3_X1 AND3_3403( .ZN(N11153), .A1(N11100), .A2(N7655), .A3(N10283) );
  AND3_X1 AND3_3404( .ZN(N11154), .A1(N11103), .A2(N9551), .A3(N10119) );
  AND3_X1 AND3_3405( .ZN(N11155), .A1(N11100), .A2(N9917), .A3(N10119) );
  NAND2_X1 NAND2_3406( .ZN(N11156), .A1(N11137), .A2(N11107) );
  NAND2_X1 NAND2_3407( .ZN(N11159), .A1(N11138), .A2(N11109) );
  NAND2_X1 NAND2_3408( .ZN(N11162), .A1(N11139), .A2(N11111) );
  NAND2_X1 NAND2_3409( .ZN(N11165), .A1(N11140), .A2(N11113) );
  NAND2_X1 NAND2_3410( .ZN(N11168), .A1(N11141), .A2(N11115) );
  NAND2_X1 NAND2_3411( .ZN(N11171), .A1(N11142), .A2(N11117) );
  NAND2_X1 NAND2_3412( .ZN(N11174), .A1(N11143), .A2(N11119) );
  NAND2_X1 NAND2_3413( .ZN(N11177), .A1(N11144), .A2(N11121) );
  NAND2_X1 NAND2_3414( .ZN(N11180), .A1(N11145), .A2(N11123) );
  INV_X1 NOT1_3415( .ZN(N11183), .A(N11124) );
  NAND2_X1 NAND2_3416( .ZN(N11184), .A1(N11124), .A2(N9468) );
  INV_X1 NOT1_3417( .ZN(N11185), .A(N11127) );
  NAND2_X1 NAND2_3418( .ZN(N11186), .A1(N11127), .A2(N9508) );
  INV_X1 NOT1_3419( .ZN(N11187), .A(N11130) );
  NAND2_X1 NAND2_3420( .ZN(N11188), .A1(N11130), .A2(N9509) );
  OR4_X1 OR4_3421( .ZN(N11205), .A1(N11152), .A2(N11153), .A3(N11154), .A4(N11155) );
  NAND2_X1 NAND2_3422( .ZN(N11210), .A1(N8724), .A2(N11183) );
  NAND2_X1 NAND2_3423( .ZN(N11211), .A1(N8790), .A2(N11185) );
  NAND2_X1 NAND2_3424( .ZN(N11212), .A1(N8808), .A2(N11187) );
  INV_X1 NOT1_3425( .ZN(N11213), .A(N11168) );
  NAND2_X1 NAND2_3426( .ZN(N11214), .A1(N11168), .A2(N8260) );
  INV_X1 NOT1_3427( .ZN(N11215), .A(N11171) );
  NAND2_X1 NAND2_3428( .ZN(N11216), .A1(N11171), .A2(N8261) );
  INV_X1 NOT1_3429( .ZN(N11217), .A(N11174) );
  NAND2_X1 NAND2_3430( .ZN(N11218), .A1(N11174), .A2(N8296) );
  INV_X1 NOT1_3431( .ZN(N11219), .A(N11177) );
  NAND2_X1 NAND2_3432( .ZN(N11220), .A1(N11177), .A2(N8297) );
  AND3_X1 AND3_3433( .ZN(N11222), .A1(N11159), .A2(N9575), .A3(N1218) );
  AND3_X1 AND3_3434( .ZN(N11223), .A1(N11156), .A2(N8927), .A3(N1218) );
  AND3_X1 AND3_3435( .ZN(N11224), .A1(N11159), .A2(N9935), .A3(N750) );
  AND3_X1 AND3_3436( .ZN(N11225), .A1(N11156), .A2(N10132), .A3(N750) );
  AND3_X1 AND3_3437( .ZN(N11226), .A1(N11165), .A2(N9608), .A3(N10497) );
  AND3_X1 AND3_3438( .ZN(N11227), .A1(N11162), .A2(N9001), .A3(N10497) );
  AND3_X1 AND3_3439( .ZN(N11228), .A1(N11165), .A2(N9949), .A3(N10301) );
  AND3_X1 AND3_3440( .ZN(N11229), .A1(N11162), .A2(N10160), .A3(N10301) );
  INV_X1 NOT1_3441( .ZN(N11231), .A(N11180) );
  NAND2_X1 NAND2_3442( .ZN(N11232), .A1(N11180), .A2(N9467) );
  NAND2_X1 NAND2_3443( .ZN(N11233), .A1(N11210), .A2(N11184) );
  NAND2_X1 NAND2_3444( .ZN(N11236), .A1(N11211), .A2(N11186) );
  NAND2_X1 NAND2_3445( .ZN(N11239), .A1(N11212), .A2(N11188) );
  NAND2_X1 NAND2_3446( .ZN(N11242), .A1(N7459), .A2(N11213) );
  NAND2_X1 NAND2_3447( .ZN(N11243), .A1(N7462), .A2(N11215) );
  NAND2_X1 NAND2_3448( .ZN(N11244), .A1(N7515), .A2(N11217) );
  NAND2_X1 NAND2_3449( .ZN(N11245), .A1(N7518), .A2(N11219) );
  INV_X1 NOT1_3450( .ZN(N11246), .A(N11205) );
  NAND2_X1 NAND2_3451( .ZN(N11250), .A1(N8708), .A2(N11231) );
  OR4_X1 OR4_3452( .ZN(N11252), .A1(N11222), .A2(N11223), .A3(N11224), .A4(N11225) );
  OR4_X1 OR4_3453( .ZN(N11257), .A1(N11226), .A2(N11227), .A3(N11228), .A4(N11229) );
  NAND2_X1 NAND2_3454( .ZN(N11260), .A1(N11242), .A2(N11214) );
  NAND2_X1 NAND2_3455( .ZN(N11261), .A1(N11243), .A2(N11216) );
  NAND2_X1 NAND2_3456( .ZN(N11262), .A1(N11244), .A2(N11218) );
  NAND2_X1 NAND2_3457( .ZN(N11263), .A1(N11245), .A2(N11220) );
  INV_X1 NOT1_3458( .ZN(N11264), .A(N11233) );
  NAND2_X1 NAND2_3459( .ZN(N11265), .A1(N11233), .A2(N9322) );
  INV_X1 NOT1_3460( .ZN(N11267), .A(N11236) );
  NAND2_X1 NAND2_3461( .ZN(N11268), .A1(N11236), .A2(N9383) );
  INV_X1 NOT1_3462( .ZN(N11269), .A(N11239) );
  NAND2_X1 NAND2_3463( .ZN(N11270), .A1(N11239), .A2(N9384) );
  NAND2_X1 NAND2_3464( .ZN(N11272), .A1(N11250), .A2(N11232) );
  INV_X1 NOT1_3465( .ZN(N11277), .A(N11261) );
  AND2_X1 AND2_3466( .ZN(N11278), .A1(N10273), .A2(N11260) );
  INV_X1 NOT1_3467( .ZN(N11279), .A(N11263) );
  AND2_X1 AND2_3468( .ZN(N11280), .A1(N10119), .A2(N11262) );
  NAND2_X1 NAND2_3469( .ZN(N11282), .A1(N8714), .A2(N11264) );
  INV_X1 NOT1_3470( .ZN(N11283), .A(N11252) );
  NAND2_X1 NAND2_3471( .ZN(N11284), .A1(N8793), .A2(N11267) );
  NAND2_X1 NAND2_3472( .ZN(N11285), .A1(N8796), .A2(N11269) );
  INV_X1 NOT1_3473( .ZN(N11286), .A(N11257) );
  AND2_X1 AND2_3474( .ZN(N11288), .A1(N11277), .A2(N10479) );
  AND2_X1 AND2_3475( .ZN(N11289), .A1(N11279), .A2(N10283) );
  INV_X2 NOT1_3476( .ZN(N11290), .A(N11272) );
  NAND2_X1 NAND2_3477( .ZN(N11291), .A1(N11272), .A2(N9321) );
  NAND2_X1 NAND2_3478( .ZN(N11292), .A1(N11282), .A2(N11265) );
  NAND2_X1 NAND2_3479( .ZN(N11293), .A1(N11284), .A2(N11268) );
  NAND2_X1 NAND2_3480( .ZN(N11294), .A1(N11285), .A2(N11270) );
  NAND2_X1 NAND2_3481( .ZN(N11295), .A1(N8711), .A2(N11290) );
  INV_X1 NOT1_3482( .ZN(N11296), .A(N11292) );
  INV_X1 NOT1_3483( .ZN(N11297), .A(N11294) );
  AND2_X1 AND2_3484( .ZN(N11298), .A1(N10301), .A2(N11293) );
  OR2_X1 OR2_3485( .ZN(N11299), .A1(N11288), .A2(N11278) );
  OR2_X1 OR2_3486( .ZN(N11302), .A1(N11289), .A2(N11280) );
  NAND2_X1 NAND2_3487( .ZN(N11307), .A1(N11295), .A2(N11291) );
  AND2_X1 AND2_3488( .ZN(N11308), .A1(N11296), .A2(N1218) );
  AND2_X1 AND2_3489( .ZN(N11309), .A1(N11297), .A2(N10497) );
  NAND2_X1 NAND2_3490( .ZN(N11312), .A1(N11302), .A2(N11246) );
  NAND2_X1 NAND2_3491( .ZN(N11313), .A1(N11299), .A2(N10836) );
  INV_X1 NOT1_3492( .ZN(N11314), .A(N11299) );
  INV_X1 NOT1_3493( .ZN(N11315), .A(N11302) );
  AND2_X1 AND2_3494( .ZN(N11316), .A1(N750), .A2(N11307) );
  OR2_X1 OR2_3495( .ZN(N11317), .A1(N11309), .A2(N11298) );
  NAND2_X1 NAND2_3496( .ZN(N11320), .A1(N11205), .A2(N11315) );
  NAND2_X1 NAND2_3497( .ZN(N11321), .A1(N10739), .A2(N11314) );
  OR2_X1 OR2_3498( .ZN(N11323), .A1(N11308), .A2(N11316) );
  NAND2_X1 NAND2_3499( .ZN(N11327), .A1(N11312), .A2(N11320) );
  NAND2_X1 NAND2_3500( .ZN(N11328), .A1(N11313), .A2(N11321) );
  NAND2_X1 NAND2_3501( .ZN(N11329), .A1(N11317), .A2(N11286) );
  INV_X1 NOT1_3502( .ZN(N11331), .A(N11317) );
  INV_X1 NOT1_3503( .ZN(N11333), .A(N11327) );
  INV_X1 NOT1_3504( .ZN(N11334), .A(N11328) );
  NAND2_X1 NAND2_3505( .ZN(N11335), .A1(N11257), .A2(N11331) );
  NAND2_X1 NAND2_3506( .ZN(N11336), .A1(N11323), .A2(N11283) );
  INV_X1 NOT1_3507( .ZN(N11337), .A(N11323) );
  NAND2_X1 NAND2_3508( .ZN(N11338), .A1(N11329), .A2(N11335) );
  NAND2_X1 NAND2_3509( .ZN(N11339), .A1(N11252), .A2(N11337) );
  INV_X1 NOT1_3510( .ZN(N11340), .A(N11338) );
  NAND2_X1 NAND2_3511( .ZN(N11341), .A1(N11336), .A2(N11339) );
  INV_X1 NOT1_3512( .ZN(N11342), .A(N11341) );
  BUF_X1 BUFF1_3513( .Z(N241_O), .A(N241_I) );

endmodule
